magic
tech gf180mcuC
magscale 1 5
timestamp 1670238677
<< metal2 >>
rect 5516 297780 5628 298500
rect 16548 297780 16660 298500
rect 26894 297822 27538 297850
rect 27580 297836 27692 298500
rect 26894 259994 26922 297822
rect 27510 297738 27538 297822
rect 27566 297780 27692 297836
rect 38612 297780 38724 298500
rect 49644 297780 49756 298500
rect 60676 297836 60788 298500
rect 60662 297780 60788 297836
rect 71708 297780 71820 298500
rect 82740 297780 82852 298500
rect 93772 297836 93884 298500
rect 93772 297780 93898 297836
rect 104804 297780 104916 298500
rect 115836 297780 115948 298500
rect 126868 297836 126980 298500
rect 126868 297780 126994 297836
rect 137900 297780 138012 298500
rect 148932 297780 149044 298500
rect 159614 297822 159922 297850
rect 159964 297836 160076 298500
rect 27566 297738 27594 297780
rect 27510 297710 27594 297738
rect 60662 286454 60690 297780
rect 93870 295274 93898 297780
rect 126966 295330 126994 297780
rect 126966 295297 126994 295302
rect 149926 295330 149954 295335
rect 93870 295241 93898 295246
rect 60494 286426 60690 286454
rect 54166 278922 54194 278927
rect 54166 260834 54194 278894
rect 54166 260801 54194 260806
rect 60494 260050 60522 286426
rect 149926 260386 149954 295302
rect 149926 260353 149954 260358
rect 150374 295274 150402 295279
rect 60494 260017 60522 260022
rect 26894 259961 26922 259966
rect 2086 259658 2114 259663
rect 2086 258426 2114 259630
rect 2086 258393 2114 258398
rect 150374 210098 150402 295246
rect 152054 286482 152082 286487
rect 151326 260834 151354 260839
rect 151214 260386 151242 260391
rect 150430 259994 150458 259999
rect 150430 218050 150458 259966
rect 150486 259658 150514 259663
rect 150486 245882 150514 259630
rect 150486 245849 150514 245854
rect 150430 218017 150458 218022
rect 150374 210065 150402 210070
rect 151214 206122 151242 260358
rect 151270 260050 151298 260055
rect 151270 214074 151298 260022
rect 151326 241906 151354 260806
rect 151326 241873 151354 241878
rect 152054 222026 152082 286454
rect 152110 264642 152138 264647
rect 152110 226002 152138 264614
rect 159166 234402 159194 234407
rect 152110 225969 152138 225974
rect 155806 227682 155834 227687
rect 152054 221993 152082 221998
rect 151270 214041 151298 214046
rect 153286 215082 153314 215087
rect 151214 206089 151242 206094
rect 152446 181482 152474 181487
rect 151606 180194 151634 180199
rect 151606 170898 151634 180166
rect 151606 170865 151634 170870
rect 151326 169274 151354 169279
rect 151326 166922 151354 169246
rect 151326 166889 151354 166894
rect 151606 162162 151634 162167
rect 150766 142002 150794 142007
rect 150766 60130 150794 141974
rect 151606 64106 151634 162134
rect 152446 68082 152474 181454
rect 153286 91938 153314 215054
rect 153286 91905 153314 91910
rect 154126 208362 154154 208367
rect 154126 72058 154154 208334
rect 155806 76034 155834 227654
rect 159166 95914 159194 234374
rect 159614 201642 159642 297822
rect 159894 297738 159922 297822
rect 159950 297780 160076 297836
rect 170534 297822 170954 297850
rect 170996 297836 171108 298500
rect 182028 297836 182140 298500
rect 159950 297738 159978 297780
rect 159894 297710 159978 297738
rect 159614 201609 159642 201614
rect 170534 180194 170562 297822
rect 170926 297738 170954 297822
rect 170982 297780 171108 297836
rect 182014 297780 182140 297836
rect 193060 297780 193172 298500
rect 204092 297780 204204 298500
rect 215124 297836 215236 298500
rect 215110 297780 215236 297836
rect 226156 297780 226268 298500
rect 237188 297780 237300 298500
rect 248220 297780 248332 298500
rect 258734 297822 259210 297850
rect 259252 297836 259364 298500
rect 170982 297738 171010 297780
rect 170926 297710 171010 297738
rect 176806 295330 176834 295335
rect 170534 180161 170562 180166
rect 175966 295274 175994 295279
rect 175966 147042 175994 295246
rect 176806 150402 176834 295302
rect 182014 295330 182042 297780
rect 182014 295297 182042 295302
rect 204134 169274 204162 297780
rect 215110 295274 215138 297780
rect 215110 295241 215138 295246
rect 251566 280602 251594 280607
rect 204134 169241 204162 169246
rect 250726 261282 250754 261287
rect 176806 150369 176834 150374
rect 175966 147009 175994 147014
rect 250726 131082 250754 261254
rect 251566 134442 251594 280574
rect 258734 142842 258762 297822
rect 259182 297738 259210 297822
rect 259238 297780 259364 297836
rect 270284 297780 270396 298500
rect 281316 297780 281428 298500
rect 292348 297836 292460 298500
rect 292334 297780 292460 297836
rect 259238 297738 259266 297780
rect 259182 297710 259266 297738
rect 258734 142809 258762 142814
rect 292334 138642 292362 297780
rect 292334 138609 292362 138614
rect 295246 241458 295274 241463
rect 251566 134409 251594 134414
rect 250726 131049 250754 131054
rect 295246 126882 295274 241430
rect 295246 126849 295274 126854
rect 159166 95881 159194 95886
rect 166726 121842 166754 121847
rect 155806 76001 155834 76006
rect 154126 72025 154154 72030
rect 152446 68049 152474 68054
rect 151606 64073 151634 64078
rect 150766 60097 150794 60102
rect 166726 56154 166754 121814
rect 166726 56121 166754 56126
rect 295246 102690 295274 102695
rect 295246 52178 295274 102662
rect 295246 52145 295274 52150
rect 5684 -480 5796 240
rect 6636 -480 6748 240
rect 7588 -480 7700 240
rect 8540 -480 8652 240
rect 9492 -480 9604 240
rect 10444 -480 10556 240
rect 11396 -480 11508 240
rect 12348 -480 12460 240
rect 13300 -480 13412 240
rect 14252 -480 14364 240
rect 15204 -480 15316 240
rect 16156 -480 16268 240
rect 17108 -480 17220 240
rect 18060 -480 18172 240
rect 19012 -480 19124 240
rect 19964 -480 20076 240
rect 20916 -480 21028 240
rect 21868 -480 21980 240
rect 22820 -480 22932 240
rect 23772 -480 23884 240
rect 24724 -480 24836 240
rect 25676 -480 25788 240
rect 26628 -480 26740 240
rect 27580 -480 27692 240
rect 28532 -480 28644 240
rect 29484 -480 29596 240
rect 30436 -480 30548 240
rect 31388 -480 31500 240
rect 32340 -480 32452 240
rect 33292 -480 33404 240
rect 34244 -480 34356 240
rect 35196 -480 35308 240
rect 36148 -480 36260 240
rect 37100 -480 37212 240
rect 38052 -480 38164 240
rect 39004 -480 39116 240
rect 39956 -480 40068 240
rect 40908 -480 41020 240
rect 41860 -480 41972 240
rect 42812 -480 42924 240
rect 43764 -480 43876 240
rect 44716 -480 44828 240
rect 45668 -480 45780 240
rect 46620 -480 46732 240
rect 47572 -480 47684 240
rect 48524 -480 48636 240
rect 49476 -480 49588 240
rect 50428 -480 50540 240
rect 51380 -480 51492 240
rect 52332 -480 52444 240
rect 53284 -480 53396 240
rect 54236 -480 54348 240
rect 55188 -480 55300 240
rect 56140 -480 56252 240
rect 57092 -480 57204 240
rect 58044 -480 58156 240
rect 58996 -480 59108 240
rect 59948 -480 60060 240
rect 60900 -480 61012 240
rect 61852 -480 61964 240
rect 62804 -480 62916 240
rect 63756 -480 63868 240
rect 64708 -480 64820 240
rect 65660 -480 65772 240
rect 66612 -480 66724 240
rect 67564 -480 67676 240
rect 68516 -480 68628 240
rect 69468 -480 69580 240
rect 70420 -480 70532 240
rect 71372 -480 71484 240
rect 72324 -480 72436 240
rect 73276 -480 73388 240
rect 74228 -480 74340 240
rect 75180 -480 75292 240
rect 76132 -480 76244 240
rect 77084 -480 77196 240
rect 78036 -480 78148 240
rect 78988 -480 79100 240
rect 79940 -480 80052 240
rect 80892 -480 81004 240
rect 81844 -480 81956 240
rect 82796 -480 82908 240
rect 83748 -480 83860 240
rect 84700 -480 84812 240
rect 85652 -480 85764 240
rect 86604 -480 86716 240
rect 87556 -480 87668 240
rect 88508 -480 88620 240
rect 89460 -480 89572 240
rect 90412 -480 90524 240
rect 91364 -480 91476 240
rect 92316 -480 92428 240
rect 93268 -480 93380 240
rect 94220 -480 94332 240
rect 95172 -480 95284 240
rect 96124 -480 96236 240
rect 97076 -480 97188 240
rect 98028 -480 98140 240
rect 98980 -480 99092 240
rect 99932 -480 100044 240
rect 100884 -480 100996 240
rect 101836 -480 101948 240
rect 102788 -480 102900 240
rect 103740 -480 103852 240
rect 104692 -480 104804 240
rect 105644 -480 105756 240
rect 106596 -480 106708 240
rect 107548 -480 107660 240
rect 108500 -480 108612 240
rect 109452 -480 109564 240
rect 110404 -480 110516 240
rect 111356 -480 111468 240
rect 112308 -480 112420 240
rect 113260 -480 113372 240
rect 114212 -480 114324 240
rect 115164 -480 115276 240
rect 116116 -480 116228 240
rect 117068 -480 117180 240
rect 118020 -480 118132 240
rect 118972 -480 119084 240
rect 119924 -480 120036 240
rect 120876 -480 120988 240
rect 121828 -480 121940 240
rect 122780 -480 122892 240
rect 123732 -480 123844 240
rect 124684 -480 124796 240
rect 125636 -480 125748 240
rect 126588 -480 126700 240
rect 127540 -480 127652 240
rect 128492 -480 128604 240
rect 129444 -480 129556 240
rect 130396 -480 130508 240
rect 131348 -480 131460 240
rect 132300 -480 132412 240
rect 133252 -480 133364 240
rect 134204 -480 134316 240
rect 135156 -480 135268 240
rect 136108 -480 136220 240
rect 137060 -480 137172 240
rect 138012 -480 138124 240
rect 138964 -480 139076 240
rect 139916 -480 140028 240
rect 140868 -480 140980 240
rect 141820 -480 141932 240
rect 142772 -480 142884 240
rect 143724 -480 143836 240
rect 144676 -480 144788 240
rect 145628 -480 145740 240
rect 146580 -480 146692 240
rect 147532 -480 147644 240
rect 148484 -480 148596 240
rect 149436 -480 149548 240
rect 150388 -480 150500 240
rect 151340 -480 151452 240
rect 152292 -480 152404 240
rect 153244 -480 153356 240
rect 154196 -480 154308 240
rect 155148 -480 155260 240
rect 156100 -480 156212 240
rect 157052 -480 157164 240
rect 158004 -480 158116 240
rect 158956 -480 159068 240
rect 159908 -480 160020 240
rect 160860 -480 160972 240
rect 161812 -480 161924 240
rect 162764 -480 162876 240
rect 163716 -480 163828 240
rect 164668 -480 164780 240
rect 165620 -480 165732 240
rect 166572 -480 166684 240
rect 167524 -480 167636 240
rect 168476 -480 168588 240
rect 169428 -480 169540 240
rect 170380 -480 170492 240
rect 171332 -480 171444 240
rect 172284 -480 172396 240
rect 173236 -480 173348 240
rect 174188 -480 174300 240
rect 175140 -480 175252 240
rect 176092 -480 176204 240
rect 177044 -480 177156 240
rect 177996 -480 178108 240
rect 178948 -480 179060 240
rect 179900 -480 180012 240
rect 180852 -480 180964 240
rect 181804 -480 181916 240
rect 182756 -480 182868 240
rect 183708 -480 183820 240
rect 184660 -480 184772 240
rect 185612 -480 185724 240
rect 186564 -480 186676 240
rect 187516 -480 187628 240
rect 188468 -480 188580 240
rect 189420 -480 189532 240
rect 190372 -480 190484 240
rect 191324 -480 191436 240
rect 192276 -480 192388 240
rect 193228 -480 193340 240
rect 194180 -480 194292 240
rect 195132 -480 195244 240
rect 196084 -480 196196 240
rect 197036 -480 197148 240
rect 197988 -480 198100 240
rect 198940 -480 199052 240
rect 199892 -480 200004 240
rect 200844 -480 200956 240
rect 201796 -480 201908 240
rect 202748 -480 202860 240
rect 203700 -480 203812 240
rect 204652 -480 204764 240
rect 205604 -480 205716 240
rect 206556 -480 206668 240
rect 207508 -480 207620 240
rect 208460 -480 208572 240
rect 209412 -480 209524 240
rect 210364 -480 210476 240
rect 211316 -480 211428 240
rect 212268 -480 212380 240
rect 213220 -480 213332 240
rect 214172 -480 214284 240
rect 215124 -480 215236 240
rect 216076 -480 216188 240
rect 217028 -480 217140 240
rect 217980 -480 218092 240
rect 218932 -480 219044 240
rect 219884 -480 219996 240
rect 220836 -480 220948 240
rect 221788 -480 221900 240
rect 222740 -480 222852 240
rect 223692 -480 223804 240
rect 224644 -480 224756 240
rect 225596 -480 225708 240
rect 226548 -480 226660 240
rect 227500 -480 227612 240
rect 228452 -480 228564 240
rect 229404 -480 229516 240
rect 230356 -480 230468 240
rect 231308 -480 231420 240
rect 232260 -480 232372 240
rect 233212 -480 233324 240
rect 234164 -480 234276 240
rect 235116 -480 235228 240
rect 236068 -480 236180 240
rect 237020 -480 237132 240
rect 237972 -480 238084 240
rect 238924 -480 239036 240
rect 239876 -480 239988 240
rect 240828 -480 240940 240
rect 241780 -480 241892 240
rect 242732 -480 242844 240
rect 243684 -480 243796 240
rect 244636 -480 244748 240
rect 245588 -480 245700 240
rect 246540 -480 246652 240
rect 247492 -480 247604 240
rect 248444 -480 248556 240
rect 249396 -480 249508 240
rect 250348 -480 250460 240
rect 251300 -480 251412 240
rect 252252 -480 252364 240
rect 253204 -480 253316 240
rect 254156 -480 254268 240
rect 255108 -480 255220 240
rect 256060 -480 256172 240
rect 257012 -480 257124 240
rect 257964 -480 258076 240
rect 258916 -480 259028 240
rect 259868 -480 259980 240
rect 260820 -480 260932 240
rect 261772 -480 261884 240
rect 262724 -480 262836 240
rect 263676 -480 263788 240
rect 264628 -480 264740 240
rect 265580 -480 265692 240
rect 266532 -480 266644 240
rect 267484 -480 267596 240
rect 268436 -480 268548 240
rect 269388 -480 269500 240
rect 270340 -480 270452 240
rect 271292 -480 271404 240
rect 272244 -480 272356 240
rect 273196 -480 273308 240
rect 274148 -480 274260 240
rect 275100 -480 275212 240
rect 276052 -480 276164 240
rect 277004 -480 277116 240
rect 277956 -480 278068 240
rect 278908 -480 279020 240
rect 279860 -480 279972 240
rect 280812 -480 280924 240
rect 281764 -480 281876 240
rect 282716 -480 282828 240
rect 283668 -480 283780 240
rect 284620 -480 284732 240
rect 285572 -480 285684 240
rect 286524 -480 286636 240
rect 287476 -480 287588 240
rect 288428 -480 288540 240
rect 289380 -480 289492 240
rect 290332 -480 290444 240
rect 291284 -480 291396 240
rect 292236 -480 292348 240
<< via2 >>
rect 126966 295302 126994 295330
rect 149926 295302 149954 295330
rect 93870 295246 93898 295274
rect 54166 278894 54194 278922
rect 54166 260806 54194 260834
rect 149926 260358 149954 260386
rect 150374 295246 150402 295274
rect 60494 260022 60522 260050
rect 26894 259966 26922 259994
rect 2086 259630 2114 259658
rect 2086 258398 2114 258426
rect 152054 286454 152082 286482
rect 151326 260806 151354 260834
rect 151214 260358 151242 260386
rect 150430 259966 150458 259994
rect 150486 259630 150514 259658
rect 150486 245854 150514 245882
rect 150430 218022 150458 218050
rect 150374 210070 150402 210098
rect 151270 260022 151298 260050
rect 151326 241878 151354 241906
rect 152110 264614 152138 264642
rect 159166 234374 159194 234402
rect 152110 225974 152138 226002
rect 155806 227654 155834 227682
rect 152054 221998 152082 222026
rect 151270 214046 151298 214074
rect 153286 215054 153314 215082
rect 151214 206094 151242 206122
rect 152446 181454 152474 181482
rect 151606 180166 151634 180194
rect 151606 170870 151634 170898
rect 151326 169246 151354 169274
rect 151326 166894 151354 166922
rect 151606 162134 151634 162162
rect 150766 141974 150794 142002
rect 153286 91910 153314 91938
rect 154126 208334 154154 208362
rect 159614 201614 159642 201642
rect 176806 295302 176834 295330
rect 170534 180166 170562 180194
rect 175966 295246 175994 295274
rect 182014 295302 182042 295330
rect 215110 295246 215138 295274
rect 251566 280574 251594 280602
rect 204134 169246 204162 169274
rect 250726 261254 250754 261282
rect 176806 150374 176834 150402
rect 175966 147014 175994 147042
rect 258734 142814 258762 142842
rect 292334 138614 292362 138642
rect 295246 241430 295274 241458
rect 251566 134414 251594 134442
rect 250726 131054 250754 131082
rect 295246 126854 295274 126882
rect 159166 95886 159194 95914
rect 166726 121814 166754 121842
rect 155806 76006 155834 76034
rect 154126 72030 154154 72058
rect 152446 68054 152474 68082
rect 151606 64078 151634 64106
rect 150766 60102 150794 60130
rect 166726 56126 166754 56154
rect 295246 102662 295274 102690
rect 295246 52150 295274 52178
<< metal3 >>
rect 126961 295302 126966 295330
rect 126994 295302 149926 295330
rect 149954 295302 149959 295330
rect 176801 295302 176806 295330
rect 176834 295302 182014 295330
rect 182042 295302 182047 295330
rect 93865 295246 93870 295274
rect 93898 295246 150374 295274
rect 150402 295246 150407 295274
rect 175961 295246 175966 295274
rect 175994 295246 215110 295274
rect 215138 295246 215143 295274
rect 297780 294308 298500 294420
rect -480 293580 240 293692
rect 297780 287700 298500 287812
rect -480 286538 240 286636
rect -480 286524 4214 286538
rect 196 286510 4214 286524
rect 4186 286482 4214 286510
rect 4186 286454 152054 286482
rect 152082 286454 152087 286482
rect 297780 281106 298500 281204
rect 297710 281092 298500 281106
rect 297710 281078 297836 281092
rect 297710 281050 297738 281078
rect 297710 281022 297850 281050
rect 297822 280602 297850 281022
rect 251561 280574 251566 280602
rect 251594 280574 297850 280602
rect -480 279482 240 279580
rect -480 279468 266 279482
rect 196 279454 266 279468
rect 238 279426 266 279454
rect 182 279398 266 279426
rect 182 278922 210 279398
rect 182 278894 54166 278922
rect 54194 278894 54199 278922
rect 297780 274484 298500 274596
rect -480 272412 240 272524
rect 297780 267876 298500 267988
rect -480 265370 240 265468
rect -480 265356 266 265370
rect 196 265342 266 265356
rect 238 265314 266 265342
rect 182 265286 266 265314
rect 182 264642 210 265286
rect 182 264614 152110 264642
rect 152138 264614 152143 264642
rect 297780 261282 298500 261380
rect 250721 261254 250726 261282
rect 250754 261268 298500 261282
rect 250754 261254 297836 261268
rect 54161 260806 54166 260834
rect 54194 260806 151326 260834
rect 151354 260806 151359 260834
rect 149921 260358 149926 260386
rect 149954 260358 151214 260386
rect 151242 260358 151247 260386
rect 60489 260022 60494 260050
rect 60522 260022 151270 260050
rect 151298 260022 151303 260050
rect 26889 259966 26894 259994
rect 26922 259966 150430 259994
rect 150458 259966 150463 259994
rect 2081 259630 2086 259658
rect 2114 259630 150486 259658
rect 150514 259630 150519 259658
rect 196 258412 2086 258426
rect -480 258398 2086 258412
rect 2114 258398 2119 258426
rect -480 258300 240 258398
rect 297780 254660 298500 254772
rect -480 251244 240 251356
rect 297780 248052 298500 248164
rect 149940 245854 150486 245882
rect 150514 245854 150519 245882
rect -480 244188 240 244300
rect 149940 241878 151326 241906
rect 151354 241878 151359 241906
rect 297780 241458 298500 241556
rect 295241 241430 295246 241458
rect 295274 241444 298500 241458
rect 295274 241430 297836 241444
rect -480 237132 240 237244
rect 297780 234850 298500 234948
rect 297710 234836 298500 234850
rect 297710 234822 297836 234836
rect 297710 234794 297738 234822
rect 297710 234766 297850 234794
rect 297822 234402 297850 234766
rect 159161 234374 159166 234402
rect 159194 234374 297850 234402
rect -480 230076 240 230188
rect 297780 228242 298500 228340
rect 297710 228228 298500 228242
rect 297710 228214 297836 228228
rect 297710 228186 297738 228214
rect 297710 228158 297850 228186
rect 297822 227682 297850 228158
rect 155801 227654 155806 227682
rect 155834 227654 297850 227682
rect 149940 225974 152110 226002
rect 152138 225974 152143 226002
rect -480 223020 240 223132
rect 149940 221998 152054 222026
rect 152082 221998 152087 222026
rect 297780 221620 298500 221732
rect 149940 218022 150430 218050
rect 150458 218022 150463 218050
rect -480 215964 240 216076
rect 297780 215082 298500 215124
rect 153281 215054 153286 215082
rect 153314 215054 298500 215082
rect 297780 215012 298500 215054
rect 149940 214046 151270 214074
rect 151298 214046 151303 214074
rect 149940 210070 150374 210098
rect 150402 210070 150407 210098
rect -480 208908 240 209020
rect 297780 208418 298500 208516
rect 286426 208404 298500 208418
rect 286426 208390 297836 208404
rect 286426 208362 286454 208390
rect 154121 208334 154126 208362
rect 154154 208334 286454 208362
rect 149940 206094 151214 206122
rect 151242 206094 151247 206122
rect -480 201852 240 201964
rect 149926 201754 149954 202132
rect 297780 201796 298500 201908
rect 149926 201726 151214 201754
rect 151186 201642 151214 201726
rect 151186 201614 159614 201642
rect 159642 201614 159647 201642
rect 297780 195188 298500 195300
rect -480 194796 240 194908
rect 297780 188580 298500 188692
rect -480 187740 240 187852
rect 297780 181986 298500 182084
rect 297710 181972 298500 181986
rect 297710 181958 297836 181972
rect 297710 181930 297738 181958
rect 297710 181902 297850 181930
rect 297822 181482 297850 181902
rect 152441 181454 152446 181482
rect 152474 181454 297850 181482
rect -480 180684 240 180796
rect 151601 180166 151606 180194
rect 151634 180166 170534 180194
rect 170562 180166 170567 180194
rect 297780 175364 298500 175476
rect -480 173628 240 173740
rect 149940 170870 151606 170898
rect 151634 170870 151639 170898
rect 151321 169246 151326 169274
rect 151354 169246 204134 169274
rect 204162 169246 204167 169274
rect 297780 168756 298500 168868
rect 149940 166894 151326 166922
rect 151354 166894 151359 166922
rect -480 166572 240 166684
rect 297780 162162 298500 162260
rect 151601 162134 151606 162162
rect 151634 162148 298500 162162
rect 151634 162134 297836 162148
rect -480 159516 240 159628
rect 297780 155540 298500 155652
rect -480 152460 240 152572
rect 149926 150626 149954 151004
rect 149926 150598 151214 150626
rect 151186 150402 151214 150598
rect 151186 150374 176806 150402
rect 176834 150374 176839 150402
rect 297780 148932 298500 149044
rect 149940 147014 175966 147042
rect 175994 147014 175999 147042
rect -480 145404 240 145516
rect 149926 142842 149954 143052
rect 149926 142814 258734 142842
rect 258762 142814 258767 142842
rect 297780 142338 298500 142436
rect 297710 142324 298500 142338
rect 297710 142310 297836 142324
rect 297710 142282 297738 142310
rect 297710 142254 297850 142282
rect 297822 142002 297850 142254
rect 150761 141974 150766 142002
rect 150794 141974 297850 142002
rect 149926 138698 149954 139076
rect 149926 138670 151214 138698
rect 151186 138642 151214 138670
rect 151186 138614 292334 138642
rect 292362 138614 292367 138642
rect -480 138348 240 138460
rect 297780 135716 298500 135828
rect 149926 134722 149954 135100
rect 149926 134694 151214 134722
rect 151186 134442 151214 134694
rect 151186 134414 251566 134442
rect 251594 134414 251599 134442
rect -480 131292 240 131404
rect 149940 131110 151214 131138
rect 151186 131082 151214 131110
rect 151186 131054 250726 131082
rect 250754 131054 250759 131082
rect 297780 129108 298500 129220
rect 149926 126882 149954 127148
rect 149926 126854 295246 126882
rect 295274 126854 295279 126882
rect -480 124236 240 124348
rect 297780 122514 298500 122612
rect 297710 122500 298500 122514
rect 297710 122486 297836 122500
rect 297710 122458 297738 122486
rect 297710 122430 297850 122458
rect 297822 121842 297850 122430
rect 166721 121814 166726 121842
rect 166754 121814 297850 121842
rect -480 117180 240 117292
rect 297780 115892 298500 116004
rect -480 110124 240 110236
rect 297780 109284 298500 109396
rect -480 103068 240 103180
rect 297780 102690 298500 102788
rect 295241 102662 295246 102690
rect 295274 102676 298500 102690
rect 295274 102662 297836 102676
rect -480 96012 240 96124
rect 297780 96068 298500 96180
rect 119980 95886 159166 95914
rect 159194 95886 159199 95914
rect 119980 91910 153286 91938
rect 153314 91910 153319 91938
rect 297780 89460 298500 89572
rect -480 88956 240 89068
rect 297780 82852 298500 82964
rect -480 81900 240 82012
rect 297780 76244 298500 76356
rect 119980 76006 155806 76034
rect 155834 76006 155839 76034
rect -480 74844 240 74956
rect 119980 72030 154126 72058
rect 154154 72030 154159 72058
rect 297780 69636 298500 69748
rect 119980 68054 152446 68082
rect 152474 68054 152479 68082
rect -480 67788 240 67900
rect 119980 64078 151606 64106
rect 151634 64078 151639 64106
rect 297780 63028 298500 63140
rect -480 60732 240 60844
rect 119980 60102 150766 60130
rect 150794 60102 150799 60130
rect 297780 56420 298500 56532
rect 119980 56126 166726 56154
rect 166754 56126 166759 56154
rect -480 53676 240 53788
rect 119980 52150 295246 52178
rect 295274 52150 295279 52178
rect 297780 49812 298500 49924
rect -480 46620 240 46732
rect 297780 43204 298500 43316
rect -480 39564 240 39676
rect 297780 36596 298500 36708
rect -480 32508 240 32620
rect 297780 29988 298500 30100
rect -480 25452 240 25564
rect 297780 23380 298500 23492
rect -480 18396 240 18508
rect 297780 16772 298500 16884
rect -480 11340 240 11452
rect 297780 10164 298500 10276
rect -480 4284 240 4396
rect 297780 3556 298500 3668
<< metal4 >>
rect -958 299086 -648 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 -648 299086
rect -958 299024 -648 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 -648 299024
rect -958 298962 -648 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 -648 298962
rect -958 298900 -648 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 -648 298900
rect -958 293175 -648 298872
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 -648 293175
rect -958 293113 -648 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 -648 293113
rect -958 293051 -648 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 -648 293051
rect -958 292989 -648 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 -648 292989
rect -958 284175 -648 292961
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 -648 284175
rect -958 284113 -648 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 -648 284113
rect -958 284051 -648 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 -648 284051
rect -958 283989 -648 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 -648 283989
rect -958 275175 -648 283961
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 -648 275175
rect -958 275113 -648 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 -648 275113
rect -958 275051 -648 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 -648 275051
rect -958 274989 -648 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 -648 274989
rect -958 266175 -648 274961
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 -648 266175
rect -958 266113 -648 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 -648 266113
rect -958 266051 -648 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 -648 266051
rect -958 265989 -648 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 -648 265989
rect -958 257175 -648 265961
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 -648 257175
rect -958 257113 -648 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 -648 257113
rect -958 257051 -648 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 -648 257051
rect -958 256989 -648 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 -648 256989
rect -958 248175 -648 256961
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 -648 248175
rect -958 248113 -648 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 -648 248113
rect -958 248051 -648 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 -648 248051
rect -958 247989 -648 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 -648 247989
rect -958 239175 -648 247961
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 -648 239175
rect -958 239113 -648 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 -648 239113
rect -958 239051 -648 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 -648 239051
rect -958 238989 -648 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 -648 238989
rect -958 230175 -648 238961
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 -648 230175
rect -958 230113 -648 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 -648 230113
rect -958 230051 -648 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 -648 230051
rect -958 229989 -648 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 -648 229989
rect -958 221175 -648 229961
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 -648 221175
rect -958 221113 -648 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 -648 221113
rect -958 221051 -648 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 -648 221051
rect -958 220989 -648 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 -648 220989
rect -958 212175 -648 220961
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 -648 212175
rect -958 212113 -648 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 -648 212113
rect -958 212051 -648 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 -648 212051
rect -958 211989 -648 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 -648 211989
rect -958 203175 -648 211961
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 -648 203175
rect -958 203113 -648 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 -648 203113
rect -958 203051 -648 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 -648 203051
rect -958 202989 -648 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 -648 202989
rect -958 194175 -648 202961
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 -648 194175
rect -958 194113 -648 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 -648 194113
rect -958 194051 -648 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 -648 194051
rect -958 193989 -648 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 -648 193989
rect -958 185175 -648 193961
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 -648 185175
rect -958 185113 -648 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 -648 185113
rect -958 185051 -648 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 -648 185051
rect -958 184989 -648 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 -648 184989
rect -958 176175 -648 184961
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 -648 176175
rect -958 176113 -648 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 -648 176113
rect -958 176051 -648 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 -648 176051
rect -958 175989 -648 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 -648 175989
rect -958 167175 -648 175961
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 -648 167175
rect -958 167113 -648 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 -648 167113
rect -958 167051 -648 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 -648 167051
rect -958 166989 -648 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 -648 166989
rect -958 158175 -648 166961
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 -648 158175
rect -958 158113 -648 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 -648 158113
rect -958 158051 -648 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 -648 158051
rect -958 157989 -648 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 -648 157989
rect -958 149175 -648 157961
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 -648 149175
rect -958 149113 -648 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 -648 149113
rect -958 149051 -648 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 -648 149051
rect -958 148989 -648 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 -648 148989
rect -958 140175 -648 148961
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 -648 140175
rect -958 140113 -648 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 -648 140113
rect -958 140051 -648 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 -648 140051
rect -958 139989 -648 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 -648 139989
rect -958 131175 -648 139961
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 -648 131175
rect -958 131113 -648 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 -648 131113
rect -958 131051 -648 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 -648 131051
rect -958 130989 -648 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 -648 130989
rect -958 122175 -648 130961
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 -648 122175
rect -958 122113 -648 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 -648 122113
rect -958 122051 -648 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 -648 122051
rect -958 121989 -648 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 -648 121989
rect -958 113175 -648 121961
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 -648 113175
rect -958 113113 -648 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 -648 113113
rect -958 113051 -648 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 -648 113051
rect -958 112989 -648 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 -648 112989
rect -958 104175 -648 112961
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 -648 104175
rect -958 104113 -648 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 -648 104113
rect -958 104051 -648 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 -648 104051
rect -958 103989 -648 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 -648 103989
rect -958 95175 -648 103961
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 -648 95175
rect -958 95113 -648 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 -648 95113
rect -958 95051 -648 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 -648 95051
rect -958 94989 -648 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 -648 94989
rect -958 86175 -648 94961
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 -648 86175
rect -958 86113 -648 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 -648 86113
rect -958 86051 -648 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 -648 86051
rect -958 85989 -648 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 -648 85989
rect -958 77175 -648 85961
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 -648 77175
rect -958 77113 -648 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 -648 77113
rect -958 77051 -648 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 -648 77051
rect -958 76989 -648 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 -648 76989
rect -958 68175 -648 76961
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 -648 68175
rect -958 68113 -648 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 -648 68113
rect -958 68051 -648 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 -648 68051
rect -958 67989 -648 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 -648 67989
rect -958 59175 -648 67961
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 -648 59175
rect -958 59113 -648 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 -648 59113
rect -958 59051 -648 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 -648 59051
rect -958 58989 -648 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 -648 58989
rect -958 50175 -648 58961
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 -648 50175
rect -958 50113 -648 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 -648 50113
rect -958 50051 -648 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 -648 50051
rect -958 49989 -648 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 -648 49989
rect -958 41175 -648 49961
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 -648 41175
rect -958 41113 -648 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 -648 41113
rect -958 41051 -648 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 -648 41051
rect -958 40989 -648 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 -648 40989
rect -958 32175 -648 40961
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 -648 32175
rect -958 32113 -648 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 -648 32113
rect -958 32051 -648 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 -648 32051
rect -958 31989 -648 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 -648 31989
rect -958 23175 -648 31961
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 -648 23175
rect -958 23113 -648 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 -648 23113
rect -958 23051 -648 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 -648 23051
rect -958 22989 -648 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 -648 22989
rect -958 14175 -648 22961
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 -648 14175
rect -958 14113 -648 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 -648 14113
rect -958 14051 -648 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 -648 14051
rect -958 13989 -648 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 -648 13989
rect -958 5175 -648 13961
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 -648 5175
rect -958 5113 -648 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 -648 5113
rect -958 5051 -648 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 -648 5051
rect -958 4989 -648 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 -648 4989
rect -958 -560 -648 4961
rect -478 298606 -168 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 -168 298606
rect -478 298544 -168 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 -168 298544
rect -478 298482 -168 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 -168 298482
rect -478 298420 -168 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 -168 298420
rect -478 290175 -168 298392
rect -478 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 -168 290175
rect -478 290113 -168 290147
rect -478 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 -168 290113
rect -478 290051 -168 290085
rect -478 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 -168 290051
rect -478 289989 -168 290023
rect -478 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 -168 289989
rect -478 281175 -168 289961
rect -478 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 -168 281175
rect -478 281113 -168 281147
rect -478 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 -168 281113
rect -478 281051 -168 281085
rect -478 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 -168 281051
rect -478 280989 -168 281023
rect -478 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 -168 280989
rect -478 272175 -168 280961
rect -478 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 -168 272175
rect -478 272113 -168 272147
rect -478 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 -168 272113
rect -478 272051 -168 272085
rect -478 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 -168 272051
rect -478 271989 -168 272023
rect -478 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 -168 271989
rect -478 263175 -168 271961
rect -478 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 -168 263175
rect -478 263113 -168 263147
rect -478 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 -168 263113
rect -478 263051 -168 263085
rect -478 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 -168 263051
rect -478 262989 -168 263023
rect -478 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 -168 262989
rect -478 254175 -168 262961
rect -478 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 -168 254175
rect -478 254113 -168 254147
rect -478 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 -168 254113
rect -478 254051 -168 254085
rect -478 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 -168 254051
rect -478 253989 -168 254023
rect -478 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 -168 253989
rect -478 245175 -168 253961
rect -478 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 -168 245175
rect -478 245113 -168 245147
rect -478 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 -168 245113
rect -478 245051 -168 245085
rect -478 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 -168 245051
rect -478 244989 -168 245023
rect -478 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 -168 244989
rect -478 236175 -168 244961
rect -478 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 -168 236175
rect -478 236113 -168 236147
rect -478 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 -168 236113
rect -478 236051 -168 236085
rect -478 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 -168 236051
rect -478 235989 -168 236023
rect -478 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 -168 235989
rect -478 227175 -168 235961
rect -478 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 -168 227175
rect -478 227113 -168 227147
rect -478 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 -168 227113
rect -478 227051 -168 227085
rect -478 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 -168 227051
rect -478 226989 -168 227023
rect -478 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 -168 226989
rect -478 218175 -168 226961
rect -478 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 -168 218175
rect -478 218113 -168 218147
rect -478 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 -168 218113
rect -478 218051 -168 218085
rect -478 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 -168 218051
rect -478 217989 -168 218023
rect -478 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 -168 217989
rect -478 209175 -168 217961
rect -478 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 -168 209175
rect -478 209113 -168 209147
rect -478 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 -168 209113
rect -478 209051 -168 209085
rect -478 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 -168 209051
rect -478 208989 -168 209023
rect -478 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 -168 208989
rect -478 200175 -168 208961
rect -478 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 -168 200175
rect -478 200113 -168 200147
rect -478 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 -168 200113
rect -478 200051 -168 200085
rect -478 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 -168 200051
rect -478 199989 -168 200023
rect -478 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 -168 199989
rect -478 191175 -168 199961
rect -478 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 -168 191175
rect -478 191113 -168 191147
rect -478 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 -168 191113
rect -478 191051 -168 191085
rect -478 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 -168 191051
rect -478 190989 -168 191023
rect -478 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 -168 190989
rect -478 182175 -168 190961
rect -478 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 -168 182175
rect -478 182113 -168 182147
rect -478 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 -168 182113
rect -478 182051 -168 182085
rect -478 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 -168 182051
rect -478 181989 -168 182023
rect -478 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 -168 181989
rect -478 173175 -168 181961
rect -478 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 -168 173175
rect -478 173113 -168 173147
rect -478 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 -168 173113
rect -478 173051 -168 173085
rect -478 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 -168 173051
rect -478 172989 -168 173023
rect -478 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 -168 172989
rect -478 164175 -168 172961
rect -478 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 -168 164175
rect -478 164113 -168 164147
rect -478 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 -168 164113
rect -478 164051 -168 164085
rect -478 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 -168 164051
rect -478 163989 -168 164023
rect -478 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 -168 163989
rect -478 155175 -168 163961
rect -478 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 -168 155175
rect -478 155113 -168 155147
rect -478 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 -168 155113
rect -478 155051 -168 155085
rect -478 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 -168 155051
rect -478 154989 -168 155023
rect -478 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 -168 154989
rect -478 146175 -168 154961
rect -478 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 -168 146175
rect -478 146113 -168 146147
rect -478 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 -168 146113
rect -478 146051 -168 146085
rect -478 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 -168 146051
rect -478 145989 -168 146023
rect -478 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 -168 145989
rect -478 137175 -168 145961
rect -478 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 -168 137175
rect -478 137113 -168 137147
rect -478 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 -168 137113
rect -478 137051 -168 137085
rect -478 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 -168 137051
rect -478 136989 -168 137023
rect -478 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 -168 136989
rect -478 128175 -168 136961
rect -478 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 -168 128175
rect -478 128113 -168 128147
rect -478 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 -168 128113
rect -478 128051 -168 128085
rect -478 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 -168 128051
rect -478 127989 -168 128023
rect -478 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 -168 127989
rect -478 119175 -168 127961
rect -478 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 -168 119175
rect -478 119113 -168 119147
rect -478 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 -168 119113
rect -478 119051 -168 119085
rect -478 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 -168 119051
rect -478 118989 -168 119023
rect -478 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 -168 118989
rect -478 110175 -168 118961
rect -478 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 -168 110175
rect -478 110113 -168 110147
rect -478 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 -168 110113
rect -478 110051 -168 110085
rect -478 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 -168 110051
rect -478 109989 -168 110023
rect -478 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 -168 109989
rect -478 101175 -168 109961
rect -478 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 -168 101175
rect -478 101113 -168 101147
rect -478 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 -168 101113
rect -478 101051 -168 101085
rect -478 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 -168 101051
rect -478 100989 -168 101023
rect -478 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 -168 100989
rect -478 92175 -168 100961
rect -478 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 -168 92175
rect -478 92113 -168 92147
rect -478 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 -168 92113
rect -478 92051 -168 92085
rect -478 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 -168 92051
rect -478 91989 -168 92023
rect -478 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 -168 91989
rect -478 83175 -168 91961
rect -478 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 -168 83175
rect -478 83113 -168 83147
rect -478 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 -168 83113
rect -478 83051 -168 83085
rect -478 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 -168 83051
rect -478 82989 -168 83023
rect -478 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 -168 82989
rect -478 74175 -168 82961
rect -478 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 -168 74175
rect -478 74113 -168 74147
rect -478 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 -168 74113
rect -478 74051 -168 74085
rect -478 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 -168 74051
rect -478 73989 -168 74023
rect -478 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 -168 73989
rect -478 65175 -168 73961
rect -478 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 -168 65175
rect -478 65113 -168 65147
rect -478 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 -168 65113
rect -478 65051 -168 65085
rect -478 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 -168 65051
rect -478 64989 -168 65023
rect -478 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 -168 64989
rect -478 56175 -168 64961
rect -478 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 -168 56175
rect -478 56113 -168 56147
rect -478 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 -168 56113
rect -478 56051 -168 56085
rect -478 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 -168 56051
rect -478 55989 -168 56023
rect -478 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 -168 55989
rect -478 47175 -168 55961
rect -478 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 -168 47175
rect -478 47113 -168 47147
rect -478 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 -168 47113
rect -478 47051 -168 47085
rect -478 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 -168 47051
rect -478 46989 -168 47023
rect -478 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 -168 46989
rect -478 38175 -168 46961
rect -478 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 -168 38175
rect -478 38113 -168 38147
rect -478 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 -168 38113
rect -478 38051 -168 38085
rect -478 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 -168 38051
rect -478 37989 -168 38023
rect -478 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 -168 37989
rect -478 29175 -168 37961
rect -478 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 -168 29175
rect -478 29113 -168 29147
rect -478 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 -168 29113
rect -478 29051 -168 29085
rect -478 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 -168 29051
rect -478 28989 -168 29023
rect -478 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 -168 28989
rect -478 20175 -168 28961
rect -478 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 -168 20175
rect -478 20113 -168 20147
rect -478 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 -168 20113
rect -478 20051 -168 20085
rect -478 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 -168 20051
rect -478 19989 -168 20023
rect -478 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 -168 19989
rect -478 11175 -168 19961
rect -478 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 -168 11175
rect -478 11113 -168 11147
rect -478 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 -168 11113
rect -478 11051 -168 11085
rect -478 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 -168 11051
rect -478 10989 -168 11023
rect -478 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 -168 10989
rect -478 2175 -168 10961
rect -478 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 -168 2175
rect -478 2113 -168 2147
rect -478 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 -168 2113
rect -478 2051 -168 2085
rect -478 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 -168 2051
rect -478 1989 -168 2023
rect -478 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 -168 1989
rect -478 -80 -168 1961
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 -168 -80
rect -478 -142 -168 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 -168 -142
rect -478 -204 -168 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 -168 -204
rect -478 -266 -168 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 -168 -266
rect -478 -342 -168 -294
rect 1577 298606 1887 299134
rect 1577 298578 1625 298606
rect 1653 298578 1687 298606
rect 1715 298578 1749 298606
rect 1777 298578 1811 298606
rect 1839 298578 1887 298606
rect 1577 298544 1887 298578
rect 1577 298516 1625 298544
rect 1653 298516 1687 298544
rect 1715 298516 1749 298544
rect 1777 298516 1811 298544
rect 1839 298516 1887 298544
rect 1577 298482 1887 298516
rect 1577 298454 1625 298482
rect 1653 298454 1687 298482
rect 1715 298454 1749 298482
rect 1777 298454 1811 298482
rect 1839 298454 1887 298482
rect 1577 298420 1887 298454
rect 1577 298392 1625 298420
rect 1653 298392 1687 298420
rect 1715 298392 1749 298420
rect 1777 298392 1811 298420
rect 1839 298392 1887 298420
rect 1577 290175 1887 298392
rect 1577 290147 1625 290175
rect 1653 290147 1687 290175
rect 1715 290147 1749 290175
rect 1777 290147 1811 290175
rect 1839 290147 1887 290175
rect 1577 290113 1887 290147
rect 1577 290085 1625 290113
rect 1653 290085 1687 290113
rect 1715 290085 1749 290113
rect 1777 290085 1811 290113
rect 1839 290085 1887 290113
rect 1577 290051 1887 290085
rect 1577 290023 1625 290051
rect 1653 290023 1687 290051
rect 1715 290023 1749 290051
rect 1777 290023 1811 290051
rect 1839 290023 1887 290051
rect 1577 289989 1887 290023
rect 1577 289961 1625 289989
rect 1653 289961 1687 289989
rect 1715 289961 1749 289989
rect 1777 289961 1811 289989
rect 1839 289961 1887 289989
rect 1577 281175 1887 289961
rect 1577 281147 1625 281175
rect 1653 281147 1687 281175
rect 1715 281147 1749 281175
rect 1777 281147 1811 281175
rect 1839 281147 1887 281175
rect 1577 281113 1887 281147
rect 1577 281085 1625 281113
rect 1653 281085 1687 281113
rect 1715 281085 1749 281113
rect 1777 281085 1811 281113
rect 1839 281085 1887 281113
rect 1577 281051 1887 281085
rect 1577 281023 1625 281051
rect 1653 281023 1687 281051
rect 1715 281023 1749 281051
rect 1777 281023 1811 281051
rect 1839 281023 1887 281051
rect 1577 280989 1887 281023
rect 1577 280961 1625 280989
rect 1653 280961 1687 280989
rect 1715 280961 1749 280989
rect 1777 280961 1811 280989
rect 1839 280961 1887 280989
rect 1577 272175 1887 280961
rect 1577 272147 1625 272175
rect 1653 272147 1687 272175
rect 1715 272147 1749 272175
rect 1777 272147 1811 272175
rect 1839 272147 1887 272175
rect 1577 272113 1887 272147
rect 1577 272085 1625 272113
rect 1653 272085 1687 272113
rect 1715 272085 1749 272113
rect 1777 272085 1811 272113
rect 1839 272085 1887 272113
rect 1577 272051 1887 272085
rect 1577 272023 1625 272051
rect 1653 272023 1687 272051
rect 1715 272023 1749 272051
rect 1777 272023 1811 272051
rect 1839 272023 1887 272051
rect 1577 271989 1887 272023
rect 1577 271961 1625 271989
rect 1653 271961 1687 271989
rect 1715 271961 1749 271989
rect 1777 271961 1811 271989
rect 1839 271961 1887 271989
rect 1577 263175 1887 271961
rect 1577 263147 1625 263175
rect 1653 263147 1687 263175
rect 1715 263147 1749 263175
rect 1777 263147 1811 263175
rect 1839 263147 1887 263175
rect 1577 263113 1887 263147
rect 1577 263085 1625 263113
rect 1653 263085 1687 263113
rect 1715 263085 1749 263113
rect 1777 263085 1811 263113
rect 1839 263085 1887 263113
rect 1577 263051 1887 263085
rect 1577 263023 1625 263051
rect 1653 263023 1687 263051
rect 1715 263023 1749 263051
rect 1777 263023 1811 263051
rect 1839 263023 1887 263051
rect 1577 262989 1887 263023
rect 1577 262961 1625 262989
rect 1653 262961 1687 262989
rect 1715 262961 1749 262989
rect 1777 262961 1811 262989
rect 1839 262961 1887 262989
rect 1577 254175 1887 262961
rect 1577 254147 1625 254175
rect 1653 254147 1687 254175
rect 1715 254147 1749 254175
rect 1777 254147 1811 254175
rect 1839 254147 1887 254175
rect 1577 254113 1887 254147
rect 1577 254085 1625 254113
rect 1653 254085 1687 254113
rect 1715 254085 1749 254113
rect 1777 254085 1811 254113
rect 1839 254085 1887 254113
rect 1577 254051 1887 254085
rect 1577 254023 1625 254051
rect 1653 254023 1687 254051
rect 1715 254023 1749 254051
rect 1777 254023 1811 254051
rect 1839 254023 1887 254051
rect 1577 253989 1887 254023
rect 1577 253961 1625 253989
rect 1653 253961 1687 253989
rect 1715 253961 1749 253989
rect 1777 253961 1811 253989
rect 1839 253961 1887 253989
rect 1577 245175 1887 253961
rect 1577 245147 1625 245175
rect 1653 245147 1687 245175
rect 1715 245147 1749 245175
rect 1777 245147 1811 245175
rect 1839 245147 1887 245175
rect 1577 245113 1887 245147
rect 1577 245085 1625 245113
rect 1653 245085 1687 245113
rect 1715 245085 1749 245113
rect 1777 245085 1811 245113
rect 1839 245085 1887 245113
rect 1577 245051 1887 245085
rect 1577 245023 1625 245051
rect 1653 245023 1687 245051
rect 1715 245023 1749 245051
rect 1777 245023 1811 245051
rect 1839 245023 1887 245051
rect 1577 244989 1887 245023
rect 1577 244961 1625 244989
rect 1653 244961 1687 244989
rect 1715 244961 1749 244989
rect 1777 244961 1811 244989
rect 1839 244961 1887 244989
rect 1577 236175 1887 244961
rect 1577 236147 1625 236175
rect 1653 236147 1687 236175
rect 1715 236147 1749 236175
rect 1777 236147 1811 236175
rect 1839 236147 1887 236175
rect 1577 236113 1887 236147
rect 1577 236085 1625 236113
rect 1653 236085 1687 236113
rect 1715 236085 1749 236113
rect 1777 236085 1811 236113
rect 1839 236085 1887 236113
rect 1577 236051 1887 236085
rect 1577 236023 1625 236051
rect 1653 236023 1687 236051
rect 1715 236023 1749 236051
rect 1777 236023 1811 236051
rect 1839 236023 1887 236051
rect 1577 235989 1887 236023
rect 1577 235961 1625 235989
rect 1653 235961 1687 235989
rect 1715 235961 1749 235989
rect 1777 235961 1811 235989
rect 1839 235961 1887 235989
rect 1577 227175 1887 235961
rect 1577 227147 1625 227175
rect 1653 227147 1687 227175
rect 1715 227147 1749 227175
rect 1777 227147 1811 227175
rect 1839 227147 1887 227175
rect 1577 227113 1887 227147
rect 1577 227085 1625 227113
rect 1653 227085 1687 227113
rect 1715 227085 1749 227113
rect 1777 227085 1811 227113
rect 1839 227085 1887 227113
rect 1577 227051 1887 227085
rect 1577 227023 1625 227051
rect 1653 227023 1687 227051
rect 1715 227023 1749 227051
rect 1777 227023 1811 227051
rect 1839 227023 1887 227051
rect 1577 226989 1887 227023
rect 1577 226961 1625 226989
rect 1653 226961 1687 226989
rect 1715 226961 1749 226989
rect 1777 226961 1811 226989
rect 1839 226961 1887 226989
rect 1577 218175 1887 226961
rect 1577 218147 1625 218175
rect 1653 218147 1687 218175
rect 1715 218147 1749 218175
rect 1777 218147 1811 218175
rect 1839 218147 1887 218175
rect 1577 218113 1887 218147
rect 1577 218085 1625 218113
rect 1653 218085 1687 218113
rect 1715 218085 1749 218113
rect 1777 218085 1811 218113
rect 1839 218085 1887 218113
rect 1577 218051 1887 218085
rect 1577 218023 1625 218051
rect 1653 218023 1687 218051
rect 1715 218023 1749 218051
rect 1777 218023 1811 218051
rect 1839 218023 1887 218051
rect 1577 217989 1887 218023
rect 1577 217961 1625 217989
rect 1653 217961 1687 217989
rect 1715 217961 1749 217989
rect 1777 217961 1811 217989
rect 1839 217961 1887 217989
rect 1577 209175 1887 217961
rect 1577 209147 1625 209175
rect 1653 209147 1687 209175
rect 1715 209147 1749 209175
rect 1777 209147 1811 209175
rect 1839 209147 1887 209175
rect 1577 209113 1887 209147
rect 1577 209085 1625 209113
rect 1653 209085 1687 209113
rect 1715 209085 1749 209113
rect 1777 209085 1811 209113
rect 1839 209085 1887 209113
rect 1577 209051 1887 209085
rect 1577 209023 1625 209051
rect 1653 209023 1687 209051
rect 1715 209023 1749 209051
rect 1777 209023 1811 209051
rect 1839 209023 1887 209051
rect 1577 208989 1887 209023
rect 1577 208961 1625 208989
rect 1653 208961 1687 208989
rect 1715 208961 1749 208989
rect 1777 208961 1811 208989
rect 1839 208961 1887 208989
rect 1577 200175 1887 208961
rect 1577 200147 1625 200175
rect 1653 200147 1687 200175
rect 1715 200147 1749 200175
rect 1777 200147 1811 200175
rect 1839 200147 1887 200175
rect 1577 200113 1887 200147
rect 1577 200085 1625 200113
rect 1653 200085 1687 200113
rect 1715 200085 1749 200113
rect 1777 200085 1811 200113
rect 1839 200085 1887 200113
rect 1577 200051 1887 200085
rect 1577 200023 1625 200051
rect 1653 200023 1687 200051
rect 1715 200023 1749 200051
rect 1777 200023 1811 200051
rect 1839 200023 1887 200051
rect 1577 199989 1887 200023
rect 1577 199961 1625 199989
rect 1653 199961 1687 199989
rect 1715 199961 1749 199989
rect 1777 199961 1811 199989
rect 1839 199961 1887 199989
rect 1577 191175 1887 199961
rect 1577 191147 1625 191175
rect 1653 191147 1687 191175
rect 1715 191147 1749 191175
rect 1777 191147 1811 191175
rect 1839 191147 1887 191175
rect 1577 191113 1887 191147
rect 1577 191085 1625 191113
rect 1653 191085 1687 191113
rect 1715 191085 1749 191113
rect 1777 191085 1811 191113
rect 1839 191085 1887 191113
rect 1577 191051 1887 191085
rect 1577 191023 1625 191051
rect 1653 191023 1687 191051
rect 1715 191023 1749 191051
rect 1777 191023 1811 191051
rect 1839 191023 1887 191051
rect 1577 190989 1887 191023
rect 1577 190961 1625 190989
rect 1653 190961 1687 190989
rect 1715 190961 1749 190989
rect 1777 190961 1811 190989
rect 1839 190961 1887 190989
rect 1577 182175 1887 190961
rect 1577 182147 1625 182175
rect 1653 182147 1687 182175
rect 1715 182147 1749 182175
rect 1777 182147 1811 182175
rect 1839 182147 1887 182175
rect 1577 182113 1887 182147
rect 1577 182085 1625 182113
rect 1653 182085 1687 182113
rect 1715 182085 1749 182113
rect 1777 182085 1811 182113
rect 1839 182085 1887 182113
rect 1577 182051 1887 182085
rect 1577 182023 1625 182051
rect 1653 182023 1687 182051
rect 1715 182023 1749 182051
rect 1777 182023 1811 182051
rect 1839 182023 1887 182051
rect 1577 181989 1887 182023
rect 1577 181961 1625 181989
rect 1653 181961 1687 181989
rect 1715 181961 1749 181989
rect 1777 181961 1811 181989
rect 1839 181961 1887 181989
rect 1577 173175 1887 181961
rect 1577 173147 1625 173175
rect 1653 173147 1687 173175
rect 1715 173147 1749 173175
rect 1777 173147 1811 173175
rect 1839 173147 1887 173175
rect 1577 173113 1887 173147
rect 1577 173085 1625 173113
rect 1653 173085 1687 173113
rect 1715 173085 1749 173113
rect 1777 173085 1811 173113
rect 1839 173085 1887 173113
rect 1577 173051 1887 173085
rect 1577 173023 1625 173051
rect 1653 173023 1687 173051
rect 1715 173023 1749 173051
rect 1777 173023 1811 173051
rect 1839 173023 1887 173051
rect 1577 172989 1887 173023
rect 1577 172961 1625 172989
rect 1653 172961 1687 172989
rect 1715 172961 1749 172989
rect 1777 172961 1811 172989
rect 1839 172961 1887 172989
rect 1577 164175 1887 172961
rect 1577 164147 1625 164175
rect 1653 164147 1687 164175
rect 1715 164147 1749 164175
rect 1777 164147 1811 164175
rect 1839 164147 1887 164175
rect 1577 164113 1887 164147
rect 1577 164085 1625 164113
rect 1653 164085 1687 164113
rect 1715 164085 1749 164113
rect 1777 164085 1811 164113
rect 1839 164085 1887 164113
rect 1577 164051 1887 164085
rect 1577 164023 1625 164051
rect 1653 164023 1687 164051
rect 1715 164023 1749 164051
rect 1777 164023 1811 164051
rect 1839 164023 1887 164051
rect 1577 163989 1887 164023
rect 1577 163961 1625 163989
rect 1653 163961 1687 163989
rect 1715 163961 1749 163989
rect 1777 163961 1811 163989
rect 1839 163961 1887 163989
rect 1577 155175 1887 163961
rect 1577 155147 1625 155175
rect 1653 155147 1687 155175
rect 1715 155147 1749 155175
rect 1777 155147 1811 155175
rect 1839 155147 1887 155175
rect 1577 155113 1887 155147
rect 1577 155085 1625 155113
rect 1653 155085 1687 155113
rect 1715 155085 1749 155113
rect 1777 155085 1811 155113
rect 1839 155085 1887 155113
rect 1577 155051 1887 155085
rect 1577 155023 1625 155051
rect 1653 155023 1687 155051
rect 1715 155023 1749 155051
rect 1777 155023 1811 155051
rect 1839 155023 1887 155051
rect 1577 154989 1887 155023
rect 1577 154961 1625 154989
rect 1653 154961 1687 154989
rect 1715 154961 1749 154989
rect 1777 154961 1811 154989
rect 1839 154961 1887 154989
rect 1577 146175 1887 154961
rect 1577 146147 1625 146175
rect 1653 146147 1687 146175
rect 1715 146147 1749 146175
rect 1777 146147 1811 146175
rect 1839 146147 1887 146175
rect 1577 146113 1887 146147
rect 1577 146085 1625 146113
rect 1653 146085 1687 146113
rect 1715 146085 1749 146113
rect 1777 146085 1811 146113
rect 1839 146085 1887 146113
rect 1577 146051 1887 146085
rect 1577 146023 1625 146051
rect 1653 146023 1687 146051
rect 1715 146023 1749 146051
rect 1777 146023 1811 146051
rect 1839 146023 1887 146051
rect 1577 145989 1887 146023
rect 1577 145961 1625 145989
rect 1653 145961 1687 145989
rect 1715 145961 1749 145989
rect 1777 145961 1811 145989
rect 1839 145961 1887 145989
rect 1577 137175 1887 145961
rect 1577 137147 1625 137175
rect 1653 137147 1687 137175
rect 1715 137147 1749 137175
rect 1777 137147 1811 137175
rect 1839 137147 1887 137175
rect 1577 137113 1887 137147
rect 1577 137085 1625 137113
rect 1653 137085 1687 137113
rect 1715 137085 1749 137113
rect 1777 137085 1811 137113
rect 1839 137085 1887 137113
rect 1577 137051 1887 137085
rect 1577 137023 1625 137051
rect 1653 137023 1687 137051
rect 1715 137023 1749 137051
rect 1777 137023 1811 137051
rect 1839 137023 1887 137051
rect 1577 136989 1887 137023
rect 1577 136961 1625 136989
rect 1653 136961 1687 136989
rect 1715 136961 1749 136989
rect 1777 136961 1811 136989
rect 1839 136961 1887 136989
rect 1577 128175 1887 136961
rect 1577 128147 1625 128175
rect 1653 128147 1687 128175
rect 1715 128147 1749 128175
rect 1777 128147 1811 128175
rect 1839 128147 1887 128175
rect 1577 128113 1887 128147
rect 1577 128085 1625 128113
rect 1653 128085 1687 128113
rect 1715 128085 1749 128113
rect 1777 128085 1811 128113
rect 1839 128085 1887 128113
rect 1577 128051 1887 128085
rect 1577 128023 1625 128051
rect 1653 128023 1687 128051
rect 1715 128023 1749 128051
rect 1777 128023 1811 128051
rect 1839 128023 1887 128051
rect 1577 127989 1887 128023
rect 1577 127961 1625 127989
rect 1653 127961 1687 127989
rect 1715 127961 1749 127989
rect 1777 127961 1811 127989
rect 1839 127961 1887 127989
rect 1577 119175 1887 127961
rect 1577 119147 1625 119175
rect 1653 119147 1687 119175
rect 1715 119147 1749 119175
rect 1777 119147 1811 119175
rect 1839 119147 1887 119175
rect 1577 119113 1887 119147
rect 1577 119085 1625 119113
rect 1653 119085 1687 119113
rect 1715 119085 1749 119113
rect 1777 119085 1811 119113
rect 1839 119085 1887 119113
rect 1577 119051 1887 119085
rect 1577 119023 1625 119051
rect 1653 119023 1687 119051
rect 1715 119023 1749 119051
rect 1777 119023 1811 119051
rect 1839 119023 1887 119051
rect 1577 118989 1887 119023
rect 1577 118961 1625 118989
rect 1653 118961 1687 118989
rect 1715 118961 1749 118989
rect 1777 118961 1811 118989
rect 1839 118961 1887 118989
rect 1577 110175 1887 118961
rect 1577 110147 1625 110175
rect 1653 110147 1687 110175
rect 1715 110147 1749 110175
rect 1777 110147 1811 110175
rect 1839 110147 1887 110175
rect 1577 110113 1887 110147
rect 1577 110085 1625 110113
rect 1653 110085 1687 110113
rect 1715 110085 1749 110113
rect 1777 110085 1811 110113
rect 1839 110085 1887 110113
rect 1577 110051 1887 110085
rect 1577 110023 1625 110051
rect 1653 110023 1687 110051
rect 1715 110023 1749 110051
rect 1777 110023 1811 110051
rect 1839 110023 1887 110051
rect 1577 109989 1887 110023
rect 1577 109961 1625 109989
rect 1653 109961 1687 109989
rect 1715 109961 1749 109989
rect 1777 109961 1811 109989
rect 1839 109961 1887 109989
rect 1577 101175 1887 109961
rect 1577 101147 1625 101175
rect 1653 101147 1687 101175
rect 1715 101147 1749 101175
rect 1777 101147 1811 101175
rect 1839 101147 1887 101175
rect 1577 101113 1887 101147
rect 1577 101085 1625 101113
rect 1653 101085 1687 101113
rect 1715 101085 1749 101113
rect 1777 101085 1811 101113
rect 1839 101085 1887 101113
rect 1577 101051 1887 101085
rect 1577 101023 1625 101051
rect 1653 101023 1687 101051
rect 1715 101023 1749 101051
rect 1777 101023 1811 101051
rect 1839 101023 1887 101051
rect 1577 100989 1887 101023
rect 1577 100961 1625 100989
rect 1653 100961 1687 100989
rect 1715 100961 1749 100989
rect 1777 100961 1811 100989
rect 1839 100961 1887 100989
rect 1577 92175 1887 100961
rect 1577 92147 1625 92175
rect 1653 92147 1687 92175
rect 1715 92147 1749 92175
rect 1777 92147 1811 92175
rect 1839 92147 1887 92175
rect 1577 92113 1887 92147
rect 1577 92085 1625 92113
rect 1653 92085 1687 92113
rect 1715 92085 1749 92113
rect 1777 92085 1811 92113
rect 1839 92085 1887 92113
rect 1577 92051 1887 92085
rect 1577 92023 1625 92051
rect 1653 92023 1687 92051
rect 1715 92023 1749 92051
rect 1777 92023 1811 92051
rect 1839 92023 1887 92051
rect 1577 91989 1887 92023
rect 1577 91961 1625 91989
rect 1653 91961 1687 91989
rect 1715 91961 1749 91989
rect 1777 91961 1811 91989
rect 1839 91961 1887 91989
rect 1577 83175 1887 91961
rect 1577 83147 1625 83175
rect 1653 83147 1687 83175
rect 1715 83147 1749 83175
rect 1777 83147 1811 83175
rect 1839 83147 1887 83175
rect 1577 83113 1887 83147
rect 1577 83085 1625 83113
rect 1653 83085 1687 83113
rect 1715 83085 1749 83113
rect 1777 83085 1811 83113
rect 1839 83085 1887 83113
rect 1577 83051 1887 83085
rect 1577 83023 1625 83051
rect 1653 83023 1687 83051
rect 1715 83023 1749 83051
rect 1777 83023 1811 83051
rect 1839 83023 1887 83051
rect 1577 82989 1887 83023
rect 1577 82961 1625 82989
rect 1653 82961 1687 82989
rect 1715 82961 1749 82989
rect 1777 82961 1811 82989
rect 1839 82961 1887 82989
rect 1577 74175 1887 82961
rect 1577 74147 1625 74175
rect 1653 74147 1687 74175
rect 1715 74147 1749 74175
rect 1777 74147 1811 74175
rect 1839 74147 1887 74175
rect 1577 74113 1887 74147
rect 1577 74085 1625 74113
rect 1653 74085 1687 74113
rect 1715 74085 1749 74113
rect 1777 74085 1811 74113
rect 1839 74085 1887 74113
rect 1577 74051 1887 74085
rect 1577 74023 1625 74051
rect 1653 74023 1687 74051
rect 1715 74023 1749 74051
rect 1777 74023 1811 74051
rect 1839 74023 1887 74051
rect 1577 73989 1887 74023
rect 1577 73961 1625 73989
rect 1653 73961 1687 73989
rect 1715 73961 1749 73989
rect 1777 73961 1811 73989
rect 1839 73961 1887 73989
rect 1577 65175 1887 73961
rect 1577 65147 1625 65175
rect 1653 65147 1687 65175
rect 1715 65147 1749 65175
rect 1777 65147 1811 65175
rect 1839 65147 1887 65175
rect 1577 65113 1887 65147
rect 1577 65085 1625 65113
rect 1653 65085 1687 65113
rect 1715 65085 1749 65113
rect 1777 65085 1811 65113
rect 1839 65085 1887 65113
rect 1577 65051 1887 65085
rect 1577 65023 1625 65051
rect 1653 65023 1687 65051
rect 1715 65023 1749 65051
rect 1777 65023 1811 65051
rect 1839 65023 1887 65051
rect 1577 64989 1887 65023
rect 1577 64961 1625 64989
rect 1653 64961 1687 64989
rect 1715 64961 1749 64989
rect 1777 64961 1811 64989
rect 1839 64961 1887 64989
rect 1577 56175 1887 64961
rect 1577 56147 1625 56175
rect 1653 56147 1687 56175
rect 1715 56147 1749 56175
rect 1777 56147 1811 56175
rect 1839 56147 1887 56175
rect 1577 56113 1887 56147
rect 1577 56085 1625 56113
rect 1653 56085 1687 56113
rect 1715 56085 1749 56113
rect 1777 56085 1811 56113
rect 1839 56085 1887 56113
rect 1577 56051 1887 56085
rect 1577 56023 1625 56051
rect 1653 56023 1687 56051
rect 1715 56023 1749 56051
rect 1777 56023 1811 56051
rect 1839 56023 1887 56051
rect 1577 55989 1887 56023
rect 1577 55961 1625 55989
rect 1653 55961 1687 55989
rect 1715 55961 1749 55989
rect 1777 55961 1811 55989
rect 1839 55961 1887 55989
rect 1577 47175 1887 55961
rect 1577 47147 1625 47175
rect 1653 47147 1687 47175
rect 1715 47147 1749 47175
rect 1777 47147 1811 47175
rect 1839 47147 1887 47175
rect 1577 47113 1887 47147
rect 1577 47085 1625 47113
rect 1653 47085 1687 47113
rect 1715 47085 1749 47113
rect 1777 47085 1811 47113
rect 1839 47085 1887 47113
rect 1577 47051 1887 47085
rect 1577 47023 1625 47051
rect 1653 47023 1687 47051
rect 1715 47023 1749 47051
rect 1777 47023 1811 47051
rect 1839 47023 1887 47051
rect 1577 46989 1887 47023
rect 1577 46961 1625 46989
rect 1653 46961 1687 46989
rect 1715 46961 1749 46989
rect 1777 46961 1811 46989
rect 1839 46961 1887 46989
rect 1577 38175 1887 46961
rect 1577 38147 1625 38175
rect 1653 38147 1687 38175
rect 1715 38147 1749 38175
rect 1777 38147 1811 38175
rect 1839 38147 1887 38175
rect 1577 38113 1887 38147
rect 1577 38085 1625 38113
rect 1653 38085 1687 38113
rect 1715 38085 1749 38113
rect 1777 38085 1811 38113
rect 1839 38085 1887 38113
rect 1577 38051 1887 38085
rect 1577 38023 1625 38051
rect 1653 38023 1687 38051
rect 1715 38023 1749 38051
rect 1777 38023 1811 38051
rect 1839 38023 1887 38051
rect 1577 37989 1887 38023
rect 1577 37961 1625 37989
rect 1653 37961 1687 37989
rect 1715 37961 1749 37989
rect 1777 37961 1811 37989
rect 1839 37961 1887 37989
rect 1577 29175 1887 37961
rect 1577 29147 1625 29175
rect 1653 29147 1687 29175
rect 1715 29147 1749 29175
rect 1777 29147 1811 29175
rect 1839 29147 1887 29175
rect 1577 29113 1887 29147
rect 1577 29085 1625 29113
rect 1653 29085 1687 29113
rect 1715 29085 1749 29113
rect 1777 29085 1811 29113
rect 1839 29085 1887 29113
rect 1577 29051 1887 29085
rect 1577 29023 1625 29051
rect 1653 29023 1687 29051
rect 1715 29023 1749 29051
rect 1777 29023 1811 29051
rect 1839 29023 1887 29051
rect 1577 28989 1887 29023
rect 1577 28961 1625 28989
rect 1653 28961 1687 28989
rect 1715 28961 1749 28989
rect 1777 28961 1811 28989
rect 1839 28961 1887 28989
rect 1577 20175 1887 28961
rect 1577 20147 1625 20175
rect 1653 20147 1687 20175
rect 1715 20147 1749 20175
rect 1777 20147 1811 20175
rect 1839 20147 1887 20175
rect 1577 20113 1887 20147
rect 1577 20085 1625 20113
rect 1653 20085 1687 20113
rect 1715 20085 1749 20113
rect 1777 20085 1811 20113
rect 1839 20085 1887 20113
rect 1577 20051 1887 20085
rect 1577 20023 1625 20051
rect 1653 20023 1687 20051
rect 1715 20023 1749 20051
rect 1777 20023 1811 20051
rect 1839 20023 1887 20051
rect 1577 19989 1887 20023
rect 1577 19961 1625 19989
rect 1653 19961 1687 19989
rect 1715 19961 1749 19989
rect 1777 19961 1811 19989
rect 1839 19961 1887 19989
rect 1577 11175 1887 19961
rect 1577 11147 1625 11175
rect 1653 11147 1687 11175
rect 1715 11147 1749 11175
rect 1777 11147 1811 11175
rect 1839 11147 1887 11175
rect 1577 11113 1887 11147
rect 1577 11085 1625 11113
rect 1653 11085 1687 11113
rect 1715 11085 1749 11113
rect 1777 11085 1811 11113
rect 1839 11085 1887 11113
rect 1577 11051 1887 11085
rect 1577 11023 1625 11051
rect 1653 11023 1687 11051
rect 1715 11023 1749 11051
rect 1777 11023 1811 11051
rect 1839 11023 1887 11051
rect 1577 10989 1887 11023
rect 1577 10961 1625 10989
rect 1653 10961 1687 10989
rect 1715 10961 1749 10989
rect 1777 10961 1811 10989
rect 1839 10961 1887 10989
rect 1577 2175 1887 10961
rect 1577 2147 1625 2175
rect 1653 2147 1687 2175
rect 1715 2147 1749 2175
rect 1777 2147 1811 2175
rect 1839 2147 1887 2175
rect 1577 2113 1887 2147
rect 1577 2085 1625 2113
rect 1653 2085 1687 2113
rect 1715 2085 1749 2113
rect 1777 2085 1811 2113
rect 1839 2085 1887 2113
rect 1577 2051 1887 2085
rect 1577 2023 1625 2051
rect 1653 2023 1687 2051
rect 1715 2023 1749 2051
rect 1777 2023 1811 2051
rect 1839 2023 1887 2051
rect 1577 1989 1887 2023
rect 1577 1961 1625 1989
rect 1653 1961 1687 1989
rect 1715 1961 1749 1989
rect 1777 1961 1811 1989
rect 1839 1961 1887 1989
rect 1577 -80 1887 1961
rect 1577 -108 1625 -80
rect 1653 -108 1687 -80
rect 1715 -108 1749 -80
rect 1777 -108 1811 -80
rect 1839 -108 1887 -80
rect 1577 -142 1887 -108
rect 1577 -170 1625 -142
rect 1653 -170 1687 -142
rect 1715 -170 1749 -142
rect 1777 -170 1811 -142
rect 1839 -170 1887 -142
rect 1577 -204 1887 -170
rect 1577 -232 1625 -204
rect 1653 -232 1687 -204
rect 1715 -232 1749 -204
rect 1777 -232 1811 -204
rect 1839 -232 1887 -204
rect 1577 -266 1887 -232
rect 1577 -294 1625 -266
rect 1653 -294 1687 -266
rect 1715 -294 1749 -266
rect 1777 -294 1811 -266
rect 1839 -294 1887 -266
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 -648 -560
rect -958 -622 -648 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 -648 -622
rect -958 -684 -648 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 -648 -684
rect -958 -746 -648 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 -648 -746
rect -958 -822 -648 -774
rect 1577 -822 1887 -294
rect 3437 299086 3747 299134
rect 3437 299058 3485 299086
rect 3513 299058 3547 299086
rect 3575 299058 3609 299086
rect 3637 299058 3671 299086
rect 3699 299058 3747 299086
rect 3437 299024 3747 299058
rect 3437 298996 3485 299024
rect 3513 298996 3547 299024
rect 3575 298996 3609 299024
rect 3637 298996 3671 299024
rect 3699 298996 3747 299024
rect 3437 298962 3747 298996
rect 3437 298934 3485 298962
rect 3513 298934 3547 298962
rect 3575 298934 3609 298962
rect 3637 298934 3671 298962
rect 3699 298934 3747 298962
rect 3437 298900 3747 298934
rect 3437 298872 3485 298900
rect 3513 298872 3547 298900
rect 3575 298872 3609 298900
rect 3637 298872 3671 298900
rect 3699 298872 3747 298900
rect 3437 293175 3747 298872
rect 3437 293147 3485 293175
rect 3513 293147 3547 293175
rect 3575 293147 3609 293175
rect 3637 293147 3671 293175
rect 3699 293147 3747 293175
rect 3437 293113 3747 293147
rect 3437 293085 3485 293113
rect 3513 293085 3547 293113
rect 3575 293085 3609 293113
rect 3637 293085 3671 293113
rect 3699 293085 3747 293113
rect 3437 293051 3747 293085
rect 3437 293023 3485 293051
rect 3513 293023 3547 293051
rect 3575 293023 3609 293051
rect 3637 293023 3671 293051
rect 3699 293023 3747 293051
rect 3437 292989 3747 293023
rect 3437 292961 3485 292989
rect 3513 292961 3547 292989
rect 3575 292961 3609 292989
rect 3637 292961 3671 292989
rect 3699 292961 3747 292989
rect 3437 284175 3747 292961
rect 3437 284147 3485 284175
rect 3513 284147 3547 284175
rect 3575 284147 3609 284175
rect 3637 284147 3671 284175
rect 3699 284147 3747 284175
rect 3437 284113 3747 284147
rect 3437 284085 3485 284113
rect 3513 284085 3547 284113
rect 3575 284085 3609 284113
rect 3637 284085 3671 284113
rect 3699 284085 3747 284113
rect 3437 284051 3747 284085
rect 3437 284023 3485 284051
rect 3513 284023 3547 284051
rect 3575 284023 3609 284051
rect 3637 284023 3671 284051
rect 3699 284023 3747 284051
rect 3437 283989 3747 284023
rect 3437 283961 3485 283989
rect 3513 283961 3547 283989
rect 3575 283961 3609 283989
rect 3637 283961 3671 283989
rect 3699 283961 3747 283989
rect 3437 275175 3747 283961
rect 3437 275147 3485 275175
rect 3513 275147 3547 275175
rect 3575 275147 3609 275175
rect 3637 275147 3671 275175
rect 3699 275147 3747 275175
rect 3437 275113 3747 275147
rect 3437 275085 3485 275113
rect 3513 275085 3547 275113
rect 3575 275085 3609 275113
rect 3637 275085 3671 275113
rect 3699 275085 3747 275113
rect 3437 275051 3747 275085
rect 3437 275023 3485 275051
rect 3513 275023 3547 275051
rect 3575 275023 3609 275051
rect 3637 275023 3671 275051
rect 3699 275023 3747 275051
rect 3437 274989 3747 275023
rect 3437 274961 3485 274989
rect 3513 274961 3547 274989
rect 3575 274961 3609 274989
rect 3637 274961 3671 274989
rect 3699 274961 3747 274989
rect 3437 266175 3747 274961
rect 3437 266147 3485 266175
rect 3513 266147 3547 266175
rect 3575 266147 3609 266175
rect 3637 266147 3671 266175
rect 3699 266147 3747 266175
rect 3437 266113 3747 266147
rect 3437 266085 3485 266113
rect 3513 266085 3547 266113
rect 3575 266085 3609 266113
rect 3637 266085 3671 266113
rect 3699 266085 3747 266113
rect 3437 266051 3747 266085
rect 3437 266023 3485 266051
rect 3513 266023 3547 266051
rect 3575 266023 3609 266051
rect 3637 266023 3671 266051
rect 3699 266023 3747 266051
rect 3437 265989 3747 266023
rect 3437 265961 3485 265989
rect 3513 265961 3547 265989
rect 3575 265961 3609 265989
rect 3637 265961 3671 265989
rect 3699 265961 3747 265989
rect 3437 257175 3747 265961
rect 3437 257147 3485 257175
rect 3513 257147 3547 257175
rect 3575 257147 3609 257175
rect 3637 257147 3671 257175
rect 3699 257147 3747 257175
rect 3437 257113 3747 257147
rect 3437 257085 3485 257113
rect 3513 257085 3547 257113
rect 3575 257085 3609 257113
rect 3637 257085 3671 257113
rect 3699 257085 3747 257113
rect 3437 257051 3747 257085
rect 3437 257023 3485 257051
rect 3513 257023 3547 257051
rect 3575 257023 3609 257051
rect 3637 257023 3671 257051
rect 3699 257023 3747 257051
rect 3437 256989 3747 257023
rect 3437 256961 3485 256989
rect 3513 256961 3547 256989
rect 3575 256961 3609 256989
rect 3637 256961 3671 256989
rect 3699 256961 3747 256989
rect 3437 248175 3747 256961
rect 3437 248147 3485 248175
rect 3513 248147 3547 248175
rect 3575 248147 3609 248175
rect 3637 248147 3671 248175
rect 3699 248147 3747 248175
rect 3437 248113 3747 248147
rect 3437 248085 3485 248113
rect 3513 248085 3547 248113
rect 3575 248085 3609 248113
rect 3637 248085 3671 248113
rect 3699 248085 3747 248113
rect 3437 248051 3747 248085
rect 3437 248023 3485 248051
rect 3513 248023 3547 248051
rect 3575 248023 3609 248051
rect 3637 248023 3671 248051
rect 3699 248023 3747 248051
rect 3437 247989 3747 248023
rect 3437 247961 3485 247989
rect 3513 247961 3547 247989
rect 3575 247961 3609 247989
rect 3637 247961 3671 247989
rect 3699 247961 3747 247989
rect 3437 239175 3747 247961
rect 3437 239147 3485 239175
rect 3513 239147 3547 239175
rect 3575 239147 3609 239175
rect 3637 239147 3671 239175
rect 3699 239147 3747 239175
rect 3437 239113 3747 239147
rect 3437 239085 3485 239113
rect 3513 239085 3547 239113
rect 3575 239085 3609 239113
rect 3637 239085 3671 239113
rect 3699 239085 3747 239113
rect 3437 239051 3747 239085
rect 3437 239023 3485 239051
rect 3513 239023 3547 239051
rect 3575 239023 3609 239051
rect 3637 239023 3671 239051
rect 3699 239023 3747 239051
rect 3437 238989 3747 239023
rect 3437 238961 3485 238989
rect 3513 238961 3547 238989
rect 3575 238961 3609 238989
rect 3637 238961 3671 238989
rect 3699 238961 3747 238989
rect 3437 230175 3747 238961
rect 3437 230147 3485 230175
rect 3513 230147 3547 230175
rect 3575 230147 3609 230175
rect 3637 230147 3671 230175
rect 3699 230147 3747 230175
rect 3437 230113 3747 230147
rect 3437 230085 3485 230113
rect 3513 230085 3547 230113
rect 3575 230085 3609 230113
rect 3637 230085 3671 230113
rect 3699 230085 3747 230113
rect 3437 230051 3747 230085
rect 3437 230023 3485 230051
rect 3513 230023 3547 230051
rect 3575 230023 3609 230051
rect 3637 230023 3671 230051
rect 3699 230023 3747 230051
rect 3437 229989 3747 230023
rect 3437 229961 3485 229989
rect 3513 229961 3547 229989
rect 3575 229961 3609 229989
rect 3637 229961 3671 229989
rect 3699 229961 3747 229989
rect 3437 221175 3747 229961
rect 3437 221147 3485 221175
rect 3513 221147 3547 221175
rect 3575 221147 3609 221175
rect 3637 221147 3671 221175
rect 3699 221147 3747 221175
rect 3437 221113 3747 221147
rect 3437 221085 3485 221113
rect 3513 221085 3547 221113
rect 3575 221085 3609 221113
rect 3637 221085 3671 221113
rect 3699 221085 3747 221113
rect 3437 221051 3747 221085
rect 3437 221023 3485 221051
rect 3513 221023 3547 221051
rect 3575 221023 3609 221051
rect 3637 221023 3671 221051
rect 3699 221023 3747 221051
rect 3437 220989 3747 221023
rect 3437 220961 3485 220989
rect 3513 220961 3547 220989
rect 3575 220961 3609 220989
rect 3637 220961 3671 220989
rect 3699 220961 3747 220989
rect 3437 212175 3747 220961
rect 3437 212147 3485 212175
rect 3513 212147 3547 212175
rect 3575 212147 3609 212175
rect 3637 212147 3671 212175
rect 3699 212147 3747 212175
rect 3437 212113 3747 212147
rect 3437 212085 3485 212113
rect 3513 212085 3547 212113
rect 3575 212085 3609 212113
rect 3637 212085 3671 212113
rect 3699 212085 3747 212113
rect 3437 212051 3747 212085
rect 3437 212023 3485 212051
rect 3513 212023 3547 212051
rect 3575 212023 3609 212051
rect 3637 212023 3671 212051
rect 3699 212023 3747 212051
rect 3437 211989 3747 212023
rect 3437 211961 3485 211989
rect 3513 211961 3547 211989
rect 3575 211961 3609 211989
rect 3637 211961 3671 211989
rect 3699 211961 3747 211989
rect 3437 203175 3747 211961
rect 3437 203147 3485 203175
rect 3513 203147 3547 203175
rect 3575 203147 3609 203175
rect 3637 203147 3671 203175
rect 3699 203147 3747 203175
rect 3437 203113 3747 203147
rect 3437 203085 3485 203113
rect 3513 203085 3547 203113
rect 3575 203085 3609 203113
rect 3637 203085 3671 203113
rect 3699 203085 3747 203113
rect 3437 203051 3747 203085
rect 3437 203023 3485 203051
rect 3513 203023 3547 203051
rect 3575 203023 3609 203051
rect 3637 203023 3671 203051
rect 3699 203023 3747 203051
rect 3437 202989 3747 203023
rect 3437 202961 3485 202989
rect 3513 202961 3547 202989
rect 3575 202961 3609 202989
rect 3637 202961 3671 202989
rect 3699 202961 3747 202989
rect 3437 194175 3747 202961
rect 3437 194147 3485 194175
rect 3513 194147 3547 194175
rect 3575 194147 3609 194175
rect 3637 194147 3671 194175
rect 3699 194147 3747 194175
rect 3437 194113 3747 194147
rect 3437 194085 3485 194113
rect 3513 194085 3547 194113
rect 3575 194085 3609 194113
rect 3637 194085 3671 194113
rect 3699 194085 3747 194113
rect 3437 194051 3747 194085
rect 3437 194023 3485 194051
rect 3513 194023 3547 194051
rect 3575 194023 3609 194051
rect 3637 194023 3671 194051
rect 3699 194023 3747 194051
rect 3437 193989 3747 194023
rect 3437 193961 3485 193989
rect 3513 193961 3547 193989
rect 3575 193961 3609 193989
rect 3637 193961 3671 193989
rect 3699 193961 3747 193989
rect 3437 185175 3747 193961
rect 3437 185147 3485 185175
rect 3513 185147 3547 185175
rect 3575 185147 3609 185175
rect 3637 185147 3671 185175
rect 3699 185147 3747 185175
rect 3437 185113 3747 185147
rect 3437 185085 3485 185113
rect 3513 185085 3547 185113
rect 3575 185085 3609 185113
rect 3637 185085 3671 185113
rect 3699 185085 3747 185113
rect 3437 185051 3747 185085
rect 3437 185023 3485 185051
rect 3513 185023 3547 185051
rect 3575 185023 3609 185051
rect 3637 185023 3671 185051
rect 3699 185023 3747 185051
rect 3437 184989 3747 185023
rect 3437 184961 3485 184989
rect 3513 184961 3547 184989
rect 3575 184961 3609 184989
rect 3637 184961 3671 184989
rect 3699 184961 3747 184989
rect 3437 176175 3747 184961
rect 3437 176147 3485 176175
rect 3513 176147 3547 176175
rect 3575 176147 3609 176175
rect 3637 176147 3671 176175
rect 3699 176147 3747 176175
rect 3437 176113 3747 176147
rect 3437 176085 3485 176113
rect 3513 176085 3547 176113
rect 3575 176085 3609 176113
rect 3637 176085 3671 176113
rect 3699 176085 3747 176113
rect 3437 176051 3747 176085
rect 3437 176023 3485 176051
rect 3513 176023 3547 176051
rect 3575 176023 3609 176051
rect 3637 176023 3671 176051
rect 3699 176023 3747 176051
rect 3437 175989 3747 176023
rect 3437 175961 3485 175989
rect 3513 175961 3547 175989
rect 3575 175961 3609 175989
rect 3637 175961 3671 175989
rect 3699 175961 3747 175989
rect 3437 167175 3747 175961
rect 3437 167147 3485 167175
rect 3513 167147 3547 167175
rect 3575 167147 3609 167175
rect 3637 167147 3671 167175
rect 3699 167147 3747 167175
rect 3437 167113 3747 167147
rect 3437 167085 3485 167113
rect 3513 167085 3547 167113
rect 3575 167085 3609 167113
rect 3637 167085 3671 167113
rect 3699 167085 3747 167113
rect 3437 167051 3747 167085
rect 3437 167023 3485 167051
rect 3513 167023 3547 167051
rect 3575 167023 3609 167051
rect 3637 167023 3671 167051
rect 3699 167023 3747 167051
rect 3437 166989 3747 167023
rect 3437 166961 3485 166989
rect 3513 166961 3547 166989
rect 3575 166961 3609 166989
rect 3637 166961 3671 166989
rect 3699 166961 3747 166989
rect 3437 158175 3747 166961
rect 3437 158147 3485 158175
rect 3513 158147 3547 158175
rect 3575 158147 3609 158175
rect 3637 158147 3671 158175
rect 3699 158147 3747 158175
rect 3437 158113 3747 158147
rect 3437 158085 3485 158113
rect 3513 158085 3547 158113
rect 3575 158085 3609 158113
rect 3637 158085 3671 158113
rect 3699 158085 3747 158113
rect 3437 158051 3747 158085
rect 3437 158023 3485 158051
rect 3513 158023 3547 158051
rect 3575 158023 3609 158051
rect 3637 158023 3671 158051
rect 3699 158023 3747 158051
rect 3437 157989 3747 158023
rect 3437 157961 3485 157989
rect 3513 157961 3547 157989
rect 3575 157961 3609 157989
rect 3637 157961 3671 157989
rect 3699 157961 3747 157989
rect 3437 149175 3747 157961
rect 3437 149147 3485 149175
rect 3513 149147 3547 149175
rect 3575 149147 3609 149175
rect 3637 149147 3671 149175
rect 3699 149147 3747 149175
rect 3437 149113 3747 149147
rect 3437 149085 3485 149113
rect 3513 149085 3547 149113
rect 3575 149085 3609 149113
rect 3637 149085 3671 149113
rect 3699 149085 3747 149113
rect 3437 149051 3747 149085
rect 3437 149023 3485 149051
rect 3513 149023 3547 149051
rect 3575 149023 3609 149051
rect 3637 149023 3671 149051
rect 3699 149023 3747 149051
rect 3437 148989 3747 149023
rect 3437 148961 3485 148989
rect 3513 148961 3547 148989
rect 3575 148961 3609 148989
rect 3637 148961 3671 148989
rect 3699 148961 3747 148989
rect 3437 140175 3747 148961
rect 3437 140147 3485 140175
rect 3513 140147 3547 140175
rect 3575 140147 3609 140175
rect 3637 140147 3671 140175
rect 3699 140147 3747 140175
rect 3437 140113 3747 140147
rect 3437 140085 3485 140113
rect 3513 140085 3547 140113
rect 3575 140085 3609 140113
rect 3637 140085 3671 140113
rect 3699 140085 3747 140113
rect 3437 140051 3747 140085
rect 3437 140023 3485 140051
rect 3513 140023 3547 140051
rect 3575 140023 3609 140051
rect 3637 140023 3671 140051
rect 3699 140023 3747 140051
rect 3437 139989 3747 140023
rect 3437 139961 3485 139989
rect 3513 139961 3547 139989
rect 3575 139961 3609 139989
rect 3637 139961 3671 139989
rect 3699 139961 3747 139989
rect 3437 131175 3747 139961
rect 3437 131147 3485 131175
rect 3513 131147 3547 131175
rect 3575 131147 3609 131175
rect 3637 131147 3671 131175
rect 3699 131147 3747 131175
rect 3437 131113 3747 131147
rect 3437 131085 3485 131113
rect 3513 131085 3547 131113
rect 3575 131085 3609 131113
rect 3637 131085 3671 131113
rect 3699 131085 3747 131113
rect 3437 131051 3747 131085
rect 3437 131023 3485 131051
rect 3513 131023 3547 131051
rect 3575 131023 3609 131051
rect 3637 131023 3671 131051
rect 3699 131023 3747 131051
rect 3437 130989 3747 131023
rect 3437 130961 3485 130989
rect 3513 130961 3547 130989
rect 3575 130961 3609 130989
rect 3637 130961 3671 130989
rect 3699 130961 3747 130989
rect 3437 122175 3747 130961
rect 3437 122147 3485 122175
rect 3513 122147 3547 122175
rect 3575 122147 3609 122175
rect 3637 122147 3671 122175
rect 3699 122147 3747 122175
rect 3437 122113 3747 122147
rect 3437 122085 3485 122113
rect 3513 122085 3547 122113
rect 3575 122085 3609 122113
rect 3637 122085 3671 122113
rect 3699 122085 3747 122113
rect 3437 122051 3747 122085
rect 3437 122023 3485 122051
rect 3513 122023 3547 122051
rect 3575 122023 3609 122051
rect 3637 122023 3671 122051
rect 3699 122023 3747 122051
rect 3437 121989 3747 122023
rect 3437 121961 3485 121989
rect 3513 121961 3547 121989
rect 3575 121961 3609 121989
rect 3637 121961 3671 121989
rect 3699 121961 3747 121989
rect 3437 113175 3747 121961
rect 3437 113147 3485 113175
rect 3513 113147 3547 113175
rect 3575 113147 3609 113175
rect 3637 113147 3671 113175
rect 3699 113147 3747 113175
rect 3437 113113 3747 113147
rect 3437 113085 3485 113113
rect 3513 113085 3547 113113
rect 3575 113085 3609 113113
rect 3637 113085 3671 113113
rect 3699 113085 3747 113113
rect 3437 113051 3747 113085
rect 3437 113023 3485 113051
rect 3513 113023 3547 113051
rect 3575 113023 3609 113051
rect 3637 113023 3671 113051
rect 3699 113023 3747 113051
rect 3437 112989 3747 113023
rect 3437 112961 3485 112989
rect 3513 112961 3547 112989
rect 3575 112961 3609 112989
rect 3637 112961 3671 112989
rect 3699 112961 3747 112989
rect 3437 104175 3747 112961
rect 3437 104147 3485 104175
rect 3513 104147 3547 104175
rect 3575 104147 3609 104175
rect 3637 104147 3671 104175
rect 3699 104147 3747 104175
rect 3437 104113 3747 104147
rect 3437 104085 3485 104113
rect 3513 104085 3547 104113
rect 3575 104085 3609 104113
rect 3637 104085 3671 104113
rect 3699 104085 3747 104113
rect 3437 104051 3747 104085
rect 3437 104023 3485 104051
rect 3513 104023 3547 104051
rect 3575 104023 3609 104051
rect 3637 104023 3671 104051
rect 3699 104023 3747 104051
rect 3437 103989 3747 104023
rect 3437 103961 3485 103989
rect 3513 103961 3547 103989
rect 3575 103961 3609 103989
rect 3637 103961 3671 103989
rect 3699 103961 3747 103989
rect 3437 95175 3747 103961
rect 3437 95147 3485 95175
rect 3513 95147 3547 95175
rect 3575 95147 3609 95175
rect 3637 95147 3671 95175
rect 3699 95147 3747 95175
rect 3437 95113 3747 95147
rect 3437 95085 3485 95113
rect 3513 95085 3547 95113
rect 3575 95085 3609 95113
rect 3637 95085 3671 95113
rect 3699 95085 3747 95113
rect 3437 95051 3747 95085
rect 3437 95023 3485 95051
rect 3513 95023 3547 95051
rect 3575 95023 3609 95051
rect 3637 95023 3671 95051
rect 3699 95023 3747 95051
rect 3437 94989 3747 95023
rect 3437 94961 3485 94989
rect 3513 94961 3547 94989
rect 3575 94961 3609 94989
rect 3637 94961 3671 94989
rect 3699 94961 3747 94989
rect 3437 86175 3747 94961
rect 3437 86147 3485 86175
rect 3513 86147 3547 86175
rect 3575 86147 3609 86175
rect 3637 86147 3671 86175
rect 3699 86147 3747 86175
rect 3437 86113 3747 86147
rect 3437 86085 3485 86113
rect 3513 86085 3547 86113
rect 3575 86085 3609 86113
rect 3637 86085 3671 86113
rect 3699 86085 3747 86113
rect 3437 86051 3747 86085
rect 3437 86023 3485 86051
rect 3513 86023 3547 86051
rect 3575 86023 3609 86051
rect 3637 86023 3671 86051
rect 3699 86023 3747 86051
rect 3437 85989 3747 86023
rect 3437 85961 3485 85989
rect 3513 85961 3547 85989
rect 3575 85961 3609 85989
rect 3637 85961 3671 85989
rect 3699 85961 3747 85989
rect 3437 77175 3747 85961
rect 3437 77147 3485 77175
rect 3513 77147 3547 77175
rect 3575 77147 3609 77175
rect 3637 77147 3671 77175
rect 3699 77147 3747 77175
rect 3437 77113 3747 77147
rect 3437 77085 3485 77113
rect 3513 77085 3547 77113
rect 3575 77085 3609 77113
rect 3637 77085 3671 77113
rect 3699 77085 3747 77113
rect 3437 77051 3747 77085
rect 3437 77023 3485 77051
rect 3513 77023 3547 77051
rect 3575 77023 3609 77051
rect 3637 77023 3671 77051
rect 3699 77023 3747 77051
rect 3437 76989 3747 77023
rect 3437 76961 3485 76989
rect 3513 76961 3547 76989
rect 3575 76961 3609 76989
rect 3637 76961 3671 76989
rect 3699 76961 3747 76989
rect 3437 68175 3747 76961
rect 3437 68147 3485 68175
rect 3513 68147 3547 68175
rect 3575 68147 3609 68175
rect 3637 68147 3671 68175
rect 3699 68147 3747 68175
rect 3437 68113 3747 68147
rect 3437 68085 3485 68113
rect 3513 68085 3547 68113
rect 3575 68085 3609 68113
rect 3637 68085 3671 68113
rect 3699 68085 3747 68113
rect 3437 68051 3747 68085
rect 3437 68023 3485 68051
rect 3513 68023 3547 68051
rect 3575 68023 3609 68051
rect 3637 68023 3671 68051
rect 3699 68023 3747 68051
rect 3437 67989 3747 68023
rect 3437 67961 3485 67989
rect 3513 67961 3547 67989
rect 3575 67961 3609 67989
rect 3637 67961 3671 67989
rect 3699 67961 3747 67989
rect 3437 59175 3747 67961
rect 3437 59147 3485 59175
rect 3513 59147 3547 59175
rect 3575 59147 3609 59175
rect 3637 59147 3671 59175
rect 3699 59147 3747 59175
rect 3437 59113 3747 59147
rect 3437 59085 3485 59113
rect 3513 59085 3547 59113
rect 3575 59085 3609 59113
rect 3637 59085 3671 59113
rect 3699 59085 3747 59113
rect 3437 59051 3747 59085
rect 3437 59023 3485 59051
rect 3513 59023 3547 59051
rect 3575 59023 3609 59051
rect 3637 59023 3671 59051
rect 3699 59023 3747 59051
rect 3437 58989 3747 59023
rect 3437 58961 3485 58989
rect 3513 58961 3547 58989
rect 3575 58961 3609 58989
rect 3637 58961 3671 58989
rect 3699 58961 3747 58989
rect 3437 50175 3747 58961
rect 3437 50147 3485 50175
rect 3513 50147 3547 50175
rect 3575 50147 3609 50175
rect 3637 50147 3671 50175
rect 3699 50147 3747 50175
rect 3437 50113 3747 50147
rect 3437 50085 3485 50113
rect 3513 50085 3547 50113
rect 3575 50085 3609 50113
rect 3637 50085 3671 50113
rect 3699 50085 3747 50113
rect 3437 50051 3747 50085
rect 3437 50023 3485 50051
rect 3513 50023 3547 50051
rect 3575 50023 3609 50051
rect 3637 50023 3671 50051
rect 3699 50023 3747 50051
rect 3437 49989 3747 50023
rect 3437 49961 3485 49989
rect 3513 49961 3547 49989
rect 3575 49961 3609 49989
rect 3637 49961 3671 49989
rect 3699 49961 3747 49989
rect 3437 41175 3747 49961
rect 3437 41147 3485 41175
rect 3513 41147 3547 41175
rect 3575 41147 3609 41175
rect 3637 41147 3671 41175
rect 3699 41147 3747 41175
rect 3437 41113 3747 41147
rect 3437 41085 3485 41113
rect 3513 41085 3547 41113
rect 3575 41085 3609 41113
rect 3637 41085 3671 41113
rect 3699 41085 3747 41113
rect 3437 41051 3747 41085
rect 3437 41023 3485 41051
rect 3513 41023 3547 41051
rect 3575 41023 3609 41051
rect 3637 41023 3671 41051
rect 3699 41023 3747 41051
rect 3437 40989 3747 41023
rect 3437 40961 3485 40989
rect 3513 40961 3547 40989
rect 3575 40961 3609 40989
rect 3637 40961 3671 40989
rect 3699 40961 3747 40989
rect 3437 32175 3747 40961
rect 3437 32147 3485 32175
rect 3513 32147 3547 32175
rect 3575 32147 3609 32175
rect 3637 32147 3671 32175
rect 3699 32147 3747 32175
rect 3437 32113 3747 32147
rect 3437 32085 3485 32113
rect 3513 32085 3547 32113
rect 3575 32085 3609 32113
rect 3637 32085 3671 32113
rect 3699 32085 3747 32113
rect 3437 32051 3747 32085
rect 3437 32023 3485 32051
rect 3513 32023 3547 32051
rect 3575 32023 3609 32051
rect 3637 32023 3671 32051
rect 3699 32023 3747 32051
rect 3437 31989 3747 32023
rect 3437 31961 3485 31989
rect 3513 31961 3547 31989
rect 3575 31961 3609 31989
rect 3637 31961 3671 31989
rect 3699 31961 3747 31989
rect 3437 23175 3747 31961
rect 3437 23147 3485 23175
rect 3513 23147 3547 23175
rect 3575 23147 3609 23175
rect 3637 23147 3671 23175
rect 3699 23147 3747 23175
rect 3437 23113 3747 23147
rect 3437 23085 3485 23113
rect 3513 23085 3547 23113
rect 3575 23085 3609 23113
rect 3637 23085 3671 23113
rect 3699 23085 3747 23113
rect 3437 23051 3747 23085
rect 3437 23023 3485 23051
rect 3513 23023 3547 23051
rect 3575 23023 3609 23051
rect 3637 23023 3671 23051
rect 3699 23023 3747 23051
rect 3437 22989 3747 23023
rect 3437 22961 3485 22989
rect 3513 22961 3547 22989
rect 3575 22961 3609 22989
rect 3637 22961 3671 22989
rect 3699 22961 3747 22989
rect 3437 14175 3747 22961
rect 3437 14147 3485 14175
rect 3513 14147 3547 14175
rect 3575 14147 3609 14175
rect 3637 14147 3671 14175
rect 3699 14147 3747 14175
rect 3437 14113 3747 14147
rect 3437 14085 3485 14113
rect 3513 14085 3547 14113
rect 3575 14085 3609 14113
rect 3637 14085 3671 14113
rect 3699 14085 3747 14113
rect 3437 14051 3747 14085
rect 3437 14023 3485 14051
rect 3513 14023 3547 14051
rect 3575 14023 3609 14051
rect 3637 14023 3671 14051
rect 3699 14023 3747 14051
rect 3437 13989 3747 14023
rect 3437 13961 3485 13989
rect 3513 13961 3547 13989
rect 3575 13961 3609 13989
rect 3637 13961 3671 13989
rect 3699 13961 3747 13989
rect 3437 5175 3747 13961
rect 3437 5147 3485 5175
rect 3513 5147 3547 5175
rect 3575 5147 3609 5175
rect 3637 5147 3671 5175
rect 3699 5147 3747 5175
rect 3437 5113 3747 5147
rect 3437 5085 3485 5113
rect 3513 5085 3547 5113
rect 3575 5085 3609 5113
rect 3637 5085 3671 5113
rect 3699 5085 3747 5113
rect 3437 5051 3747 5085
rect 3437 5023 3485 5051
rect 3513 5023 3547 5051
rect 3575 5023 3609 5051
rect 3637 5023 3671 5051
rect 3699 5023 3747 5051
rect 3437 4989 3747 5023
rect 3437 4961 3485 4989
rect 3513 4961 3547 4989
rect 3575 4961 3609 4989
rect 3637 4961 3671 4989
rect 3699 4961 3747 4989
rect 3437 -560 3747 4961
rect 3437 -588 3485 -560
rect 3513 -588 3547 -560
rect 3575 -588 3609 -560
rect 3637 -588 3671 -560
rect 3699 -588 3747 -560
rect 3437 -622 3747 -588
rect 3437 -650 3485 -622
rect 3513 -650 3547 -622
rect 3575 -650 3609 -622
rect 3637 -650 3671 -622
rect 3699 -650 3747 -622
rect 3437 -684 3747 -650
rect 3437 -712 3485 -684
rect 3513 -712 3547 -684
rect 3575 -712 3609 -684
rect 3637 -712 3671 -684
rect 3699 -712 3747 -684
rect 3437 -746 3747 -712
rect 3437 -774 3485 -746
rect 3513 -774 3547 -746
rect 3575 -774 3609 -746
rect 3637 -774 3671 -746
rect 3699 -774 3747 -746
rect 3437 -822 3747 -774
rect 10577 298606 10887 299134
rect 10577 298578 10625 298606
rect 10653 298578 10687 298606
rect 10715 298578 10749 298606
rect 10777 298578 10811 298606
rect 10839 298578 10887 298606
rect 10577 298544 10887 298578
rect 10577 298516 10625 298544
rect 10653 298516 10687 298544
rect 10715 298516 10749 298544
rect 10777 298516 10811 298544
rect 10839 298516 10887 298544
rect 10577 298482 10887 298516
rect 10577 298454 10625 298482
rect 10653 298454 10687 298482
rect 10715 298454 10749 298482
rect 10777 298454 10811 298482
rect 10839 298454 10887 298482
rect 10577 298420 10887 298454
rect 10577 298392 10625 298420
rect 10653 298392 10687 298420
rect 10715 298392 10749 298420
rect 10777 298392 10811 298420
rect 10839 298392 10887 298420
rect 10577 290175 10887 298392
rect 10577 290147 10625 290175
rect 10653 290147 10687 290175
rect 10715 290147 10749 290175
rect 10777 290147 10811 290175
rect 10839 290147 10887 290175
rect 10577 290113 10887 290147
rect 10577 290085 10625 290113
rect 10653 290085 10687 290113
rect 10715 290085 10749 290113
rect 10777 290085 10811 290113
rect 10839 290085 10887 290113
rect 10577 290051 10887 290085
rect 10577 290023 10625 290051
rect 10653 290023 10687 290051
rect 10715 290023 10749 290051
rect 10777 290023 10811 290051
rect 10839 290023 10887 290051
rect 10577 289989 10887 290023
rect 10577 289961 10625 289989
rect 10653 289961 10687 289989
rect 10715 289961 10749 289989
rect 10777 289961 10811 289989
rect 10839 289961 10887 289989
rect 10577 281175 10887 289961
rect 10577 281147 10625 281175
rect 10653 281147 10687 281175
rect 10715 281147 10749 281175
rect 10777 281147 10811 281175
rect 10839 281147 10887 281175
rect 10577 281113 10887 281147
rect 10577 281085 10625 281113
rect 10653 281085 10687 281113
rect 10715 281085 10749 281113
rect 10777 281085 10811 281113
rect 10839 281085 10887 281113
rect 10577 281051 10887 281085
rect 10577 281023 10625 281051
rect 10653 281023 10687 281051
rect 10715 281023 10749 281051
rect 10777 281023 10811 281051
rect 10839 281023 10887 281051
rect 10577 280989 10887 281023
rect 10577 280961 10625 280989
rect 10653 280961 10687 280989
rect 10715 280961 10749 280989
rect 10777 280961 10811 280989
rect 10839 280961 10887 280989
rect 10577 272175 10887 280961
rect 10577 272147 10625 272175
rect 10653 272147 10687 272175
rect 10715 272147 10749 272175
rect 10777 272147 10811 272175
rect 10839 272147 10887 272175
rect 10577 272113 10887 272147
rect 10577 272085 10625 272113
rect 10653 272085 10687 272113
rect 10715 272085 10749 272113
rect 10777 272085 10811 272113
rect 10839 272085 10887 272113
rect 10577 272051 10887 272085
rect 10577 272023 10625 272051
rect 10653 272023 10687 272051
rect 10715 272023 10749 272051
rect 10777 272023 10811 272051
rect 10839 272023 10887 272051
rect 10577 271989 10887 272023
rect 10577 271961 10625 271989
rect 10653 271961 10687 271989
rect 10715 271961 10749 271989
rect 10777 271961 10811 271989
rect 10839 271961 10887 271989
rect 10577 263175 10887 271961
rect 10577 263147 10625 263175
rect 10653 263147 10687 263175
rect 10715 263147 10749 263175
rect 10777 263147 10811 263175
rect 10839 263147 10887 263175
rect 10577 263113 10887 263147
rect 10577 263085 10625 263113
rect 10653 263085 10687 263113
rect 10715 263085 10749 263113
rect 10777 263085 10811 263113
rect 10839 263085 10887 263113
rect 10577 263051 10887 263085
rect 10577 263023 10625 263051
rect 10653 263023 10687 263051
rect 10715 263023 10749 263051
rect 10777 263023 10811 263051
rect 10839 263023 10887 263051
rect 10577 262989 10887 263023
rect 10577 262961 10625 262989
rect 10653 262961 10687 262989
rect 10715 262961 10749 262989
rect 10777 262961 10811 262989
rect 10839 262961 10887 262989
rect 10577 254175 10887 262961
rect 10577 254147 10625 254175
rect 10653 254147 10687 254175
rect 10715 254147 10749 254175
rect 10777 254147 10811 254175
rect 10839 254147 10887 254175
rect 10577 254113 10887 254147
rect 10577 254085 10625 254113
rect 10653 254085 10687 254113
rect 10715 254085 10749 254113
rect 10777 254085 10811 254113
rect 10839 254085 10887 254113
rect 10577 254051 10887 254085
rect 10577 254023 10625 254051
rect 10653 254023 10687 254051
rect 10715 254023 10749 254051
rect 10777 254023 10811 254051
rect 10839 254023 10887 254051
rect 10577 253989 10887 254023
rect 10577 253961 10625 253989
rect 10653 253961 10687 253989
rect 10715 253961 10749 253989
rect 10777 253961 10811 253989
rect 10839 253961 10887 253989
rect 10577 245175 10887 253961
rect 10577 245147 10625 245175
rect 10653 245147 10687 245175
rect 10715 245147 10749 245175
rect 10777 245147 10811 245175
rect 10839 245147 10887 245175
rect 10577 245113 10887 245147
rect 10577 245085 10625 245113
rect 10653 245085 10687 245113
rect 10715 245085 10749 245113
rect 10777 245085 10811 245113
rect 10839 245085 10887 245113
rect 10577 245051 10887 245085
rect 10577 245023 10625 245051
rect 10653 245023 10687 245051
rect 10715 245023 10749 245051
rect 10777 245023 10811 245051
rect 10839 245023 10887 245051
rect 10577 244989 10887 245023
rect 10577 244961 10625 244989
rect 10653 244961 10687 244989
rect 10715 244961 10749 244989
rect 10777 244961 10811 244989
rect 10839 244961 10887 244989
rect 10577 236175 10887 244961
rect 10577 236147 10625 236175
rect 10653 236147 10687 236175
rect 10715 236147 10749 236175
rect 10777 236147 10811 236175
rect 10839 236147 10887 236175
rect 10577 236113 10887 236147
rect 10577 236085 10625 236113
rect 10653 236085 10687 236113
rect 10715 236085 10749 236113
rect 10777 236085 10811 236113
rect 10839 236085 10887 236113
rect 10577 236051 10887 236085
rect 10577 236023 10625 236051
rect 10653 236023 10687 236051
rect 10715 236023 10749 236051
rect 10777 236023 10811 236051
rect 10839 236023 10887 236051
rect 10577 235989 10887 236023
rect 10577 235961 10625 235989
rect 10653 235961 10687 235989
rect 10715 235961 10749 235989
rect 10777 235961 10811 235989
rect 10839 235961 10887 235989
rect 10577 227175 10887 235961
rect 10577 227147 10625 227175
rect 10653 227147 10687 227175
rect 10715 227147 10749 227175
rect 10777 227147 10811 227175
rect 10839 227147 10887 227175
rect 10577 227113 10887 227147
rect 10577 227085 10625 227113
rect 10653 227085 10687 227113
rect 10715 227085 10749 227113
rect 10777 227085 10811 227113
rect 10839 227085 10887 227113
rect 10577 227051 10887 227085
rect 10577 227023 10625 227051
rect 10653 227023 10687 227051
rect 10715 227023 10749 227051
rect 10777 227023 10811 227051
rect 10839 227023 10887 227051
rect 10577 226989 10887 227023
rect 10577 226961 10625 226989
rect 10653 226961 10687 226989
rect 10715 226961 10749 226989
rect 10777 226961 10811 226989
rect 10839 226961 10887 226989
rect 10577 218175 10887 226961
rect 10577 218147 10625 218175
rect 10653 218147 10687 218175
rect 10715 218147 10749 218175
rect 10777 218147 10811 218175
rect 10839 218147 10887 218175
rect 10577 218113 10887 218147
rect 10577 218085 10625 218113
rect 10653 218085 10687 218113
rect 10715 218085 10749 218113
rect 10777 218085 10811 218113
rect 10839 218085 10887 218113
rect 10577 218051 10887 218085
rect 10577 218023 10625 218051
rect 10653 218023 10687 218051
rect 10715 218023 10749 218051
rect 10777 218023 10811 218051
rect 10839 218023 10887 218051
rect 10577 217989 10887 218023
rect 10577 217961 10625 217989
rect 10653 217961 10687 217989
rect 10715 217961 10749 217989
rect 10777 217961 10811 217989
rect 10839 217961 10887 217989
rect 10577 209175 10887 217961
rect 10577 209147 10625 209175
rect 10653 209147 10687 209175
rect 10715 209147 10749 209175
rect 10777 209147 10811 209175
rect 10839 209147 10887 209175
rect 10577 209113 10887 209147
rect 10577 209085 10625 209113
rect 10653 209085 10687 209113
rect 10715 209085 10749 209113
rect 10777 209085 10811 209113
rect 10839 209085 10887 209113
rect 10577 209051 10887 209085
rect 10577 209023 10625 209051
rect 10653 209023 10687 209051
rect 10715 209023 10749 209051
rect 10777 209023 10811 209051
rect 10839 209023 10887 209051
rect 10577 208989 10887 209023
rect 10577 208961 10625 208989
rect 10653 208961 10687 208989
rect 10715 208961 10749 208989
rect 10777 208961 10811 208989
rect 10839 208961 10887 208989
rect 10577 200175 10887 208961
rect 10577 200147 10625 200175
rect 10653 200147 10687 200175
rect 10715 200147 10749 200175
rect 10777 200147 10811 200175
rect 10839 200147 10887 200175
rect 10577 200113 10887 200147
rect 10577 200085 10625 200113
rect 10653 200085 10687 200113
rect 10715 200085 10749 200113
rect 10777 200085 10811 200113
rect 10839 200085 10887 200113
rect 10577 200051 10887 200085
rect 10577 200023 10625 200051
rect 10653 200023 10687 200051
rect 10715 200023 10749 200051
rect 10777 200023 10811 200051
rect 10839 200023 10887 200051
rect 10577 199989 10887 200023
rect 10577 199961 10625 199989
rect 10653 199961 10687 199989
rect 10715 199961 10749 199989
rect 10777 199961 10811 199989
rect 10839 199961 10887 199989
rect 10577 191175 10887 199961
rect 10577 191147 10625 191175
rect 10653 191147 10687 191175
rect 10715 191147 10749 191175
rect 10777 191147 10811 191175
rect 10839 191147 10887 191175
rect 10577 191113 10887 191147
rect 10577 191085 10625 191113
rect 10653 191085 10687 191113
rect 10715 191085 10749 191113
rect 10777 191085 10811 191113
rect 10839 191085 10887 191113
rect 10577 191051 10887 191085
rect 10577 191023 10625 191051
rect 10653 191023 10687 191051
rect 10715 191023 10749 191051
rect 10777 191023 10811 191051
rect 10839 191023 10887 191051
rect 10577 190989 10887 191023
rect 10577 190961 10625 190989
rect 10653 190961 10687 190989
rect 10715 190961 10749 190989
rect 10777 190961 10811 190989
rect 10839 190961 10887 190989
rect 10577 182175 10887 190961
rect 10577 182147 10625 182175
rect 10653 182147 10687 182175
rect 10715 182147 10749 182175
rect 10777 182147 10811 182175
rect 10839 182147 10887 182175
rect 10577 182113 10887 182147
rect 10577 182085 10625 182113
rect 10653 182085 10687 182113
rect 10715 182085 10749 182113
rect 10777 182085 10811 182113
rect 10839 182085 10887 182113
rect 10577 182051 10887 182085
rect 10577 182023 10625 182051
rect 10653 182023 10687 182051
rect 10715 182023 10749 182051
rect 10777 182023 10811 182051
rect 10839 182023 10887 182051
rect 10577 181989 10887 182023
rect 10577 181961 10625 181989
rect 10653 181961 10687 181989
rect 10715 181961 10749 181989
rect 10777 181961 10811 181989
rect 10839 181961 10887 181989
rect 10577 173175 10887 181961
rect 10577 173147 10625 173175
rect 10653 173147 10687 173175
rect 10715 173147 10749 173175
rect 10777 173147 10811 173175
rect 10839 173147 10887 173175
rect 10577 173113 10887 173147
rect 10577 173085 10625 173113
rect 10653 173085 10687 173113
rect 10715 173085 10749 173113
rect 10777 173085 10811 173113
rect 10839 173085 10887 173113
rect 10577 173051 10887 173085
rect 10577 173023 10625 173051
rect 10653 173023 10687 173051
rect 10715 173023 10749 173051
rect 10777 173023 10811 173051
rect 10839 173023 10887 173051
rect 10577 172989 10887 173023
rect 10577 172961 10625 172989
rect 10653 172961 10687 172989
rect 10715 172961 10749 172989
rect 10777 172961 10811 172989
rect 10839 172961 10887 172989
rect 10577 164175 10887 172961
rect 10577 164147 10625 164175
rect 10653 164147 10687 164175
rect 10715 164147 10749 164175
rect 10777 164147 10811 164175
rect 10839 164147 10887 164175
rect 10577 164113 10887 164147
rect 10577 164085 10625 164113
rect 10653 164085 10687 164113
rect 10715 164085 10749 164113
rect 10777 164085 10811 164113
rect 10839 164085 10887 164113
rect 10577 164051 10887 164085
rect 10577 164023 10625 164051
rect 10653 164023 10687 164051
rect 10715 164023 10749 164051
rect 10777 164023 10811 164051
rect 10839 164023 10887 164051
rect 10577 163989 10887 164023
rect 10577 163961 10625 163989
rect 10653 163961 10687 163989
rect 10715 163961 10749 163989
rect 10777 163961 10811 163989
rect 10839 163961 10887 163989
rect 10577 155175 10887 163961
rect 10577 155147 10625 155175
rect 10653 155147 10687 155175
rect 10715 155147 10749 155175
rect 10777 155147 10811 155175
rect 10839 155147 10887 155175
rect 10577 155113 10887 155147
rect 10577 155085 10625 155113
rect 10653 155085 10687 155113
rect 10715 155085 10749 155113
rect 10777 155085 10811 155113
rect 10839 155085 10887 155113
rect 10577 155051 10887 155085
rect 10577 155023 10625 155051
rect 10653 155023 10687 155051
rect 10715 155023 10749 155051
rect 10777 155023 10811 155051
rect 10839 155023 10887 155051
rect 10577 154989 10887 155023
rect 10577 154961 10625 154989
rect 10653 154961 10687 154989
rect 10715 154961 10749 154989
rect 10777 154961 10811 154989
rect 10839 154961 10887 154989
rect 10577 146175 10887 154961
rect 10577 146147 10625 146175
rect 10653 146147 10687 146175
rect 10715 146147 10749 146175
rect 10777 146147 10811 146175
rect 10839 146147 10887 146175
rect 10577 146113 10887 146147
rect 10577 146085 10625 146113
rect 10653 146085 10687 146113
rect 10715 146085 10749 146113
rect 10777 146085 10811 146113
rect 10839 146085 10887 146113
rect 10577 146051 10887 146085
rect 10577 146023 10625 146051
rect 10653 146023 10687 146051
rect 10715 146023 10749 146051
rect 10777 146023 10811 146051
rect 10839 146023 10887 146051
rect 10577 145989 10887 146023
rect 10577 145961 10625 145989
rect 10653 145961 10687 145989
rect 10715 145961 10749 145989
rect 10777 145961 10811 145989
rect 10839 145961 10887 145989
rect 10577 137175 10887 145961
rect 10577 137147 10625 137175
rect 10653 137147 10687 137175
rect 10715 137147 10749 137175
rect 10777 137147 10811 137175
rect 10839 137147 10887 137175
rect 10577 137113 10887 137147
rect 10577 137085 10625 137113
rect 10653 137085 10687 137113
rect 10715 137085 10749 137113
rect 10777 137085 10811 137113
rect 10839 137085 10887 137113
rect 10577 137051 10887 137085
rect 10577 137023 10625 137051
rect 10653 137023 10687 137051
rect 10715 137023 10749 137051
rect 10777 137023 10811 137051
rect 10839 137023 10887 137051
rect 10577 136989 10887 137023
rect 10577 136961 10625 136989
rect 10653 136961 10687 136989
rect 10715 136961 10749 136989
rect 10777 136961 10811 136989
rect 10839 136961 10887 136989
rect 10577 128175 10887 136961
rect 10577 128147 10625 128175
rect 10653 128147 10687 128175
rect 10715 128147 10749 128175
rect 10777 128147 10811 128175
rect 10839 128147 10887 128175
rect 10577 128113 10887 128147
rect 10577 128085 10625 128113
rect 10653 128085 10687 128113
rect 10715 128085 10749 128113
rect 10777 128085 10811 128113
rect 10839 128085 10887 128113
rect 10577 128051 10887 128085
rect 10577 128023 10625 128051
rect 10653 128023 10687 128051
rect 10715 128023 10749 128051
rect 10777 128023 10811 128051
rect 10839 128023 10887 128051
rect 10577 127989 10887 128023
rect 10577 127961 10625 127989
rect 10653 127961 10687 127989
rect 10715 127961 10749 127989
rect 10777 127961 10811 127989
rect 10839 127961 10887 127989
rect 10577 119175 10887 127961
rect 10577 119147 10625 119175
rect 10653 119147 10687 119175
rect 10715 119147 10749 119175
rect 10777 119147 10811 119175
rect 10839 119147 10887 119175
rect 10577 119113 10887 119147
rect 10577 119085 10625 119113
rect 10653 119085 10687 119113
rect 10715 119085 10749 119113
rect 10777 119085 10811 119113
rect 10839 119085 10887 119113
rect 10577 119051 10887 119085
rect 10577 119023 10625 119051
rect 10653 119023 10687 119051
rect 10715 119023 10749 119051
rect 10777 119023 10811 119051
rect 10839 119023 10887 119051
rect 10577 118989 10887 119023
rect 10577 118961 10625 118989
rect 10653 118961 10687 118989
rect 10715 118961 10749 118989
rect 10777 118961 10811 118989
rect 10839 118961 10887 118989
rect 10577 110175 10887 118961
rect 10577 110147 10625 110175
rect 10653 110147 10687 110175
rect 10715 110147 10749 110175
rect 10777 110147 10811 110175
rect 10839 110147 10887 110175
rect 10577 110113 10887 110147
rect 10577 110085 10625 110113
rect 10653 110085 10687 110113
rect 10715 110085 10749 110113
rect 10777 110085 10811 110113
rect 10839 110085 10887 110113
rect 10577 110051 10887 110085
rect 10577 110023 10625 110051
rect 10653 110023 10687 110051
rect 10715 110023 10749 110051
rect 10777 110023 10811 110051
rect 10839 110023 10887 110051
rect 10577 109989 10887 110023
rect 10577 109961 10625 109989
rect 10653 109961 10687 109989
rect 10715 109961 10749 109989
rect 10777 109961 10811 109989
rect 10839 109961 10887 109989
rect 10577 101175 10887 109961
rect 10577 101147 10625 101175
rect 10653 101147 10687 101175
rect 10715 101147 10749 101175
rect 10777 101147 10811 101175
rect 10839 101147 10887 101175
rect 10577 101113 10887 101147
rect 10577 101085 10625 101113
rect 10653 101085 10687 101113
rect 10715 101085 10749 101113
rect 10777 101085 10811 101113
rect 10839 101085 10887 101113
rect 10577 101051 10887 101085
rect 10577 101023 10625 101051
rect 10653 101023 10687 101051
rect 10715 101023 10749 101051
rect 10777 101023 10811 101051
rect 10839 101023 10887 101051
rect 10577 100989 10887 101023
rect 10577 100961 10625 100989
rect 10653 100961 10687 100989
rect 10715 100961 10749 100989
rect 10777 100961 10811 100989
rect 10839 100961 10887 100989
rect 10577 92175 10887 100961
rect 10577 92147 10625 92175
rect 10653 92147 10687 92175
rect 10715 92147 10749 92175
rect 10777 92147 10811 92175
rect 10839 92147 10887 92175
rect 10577 92113 10887 92147
rect 10577 92085 10625 92113
rect 10653 92085 10687 92113
rect 10715 92085 10749 92113
rect 10777 92085 10811 92113
rect 10839 92085 10887 92113
rect 10577 92051 10887 92085
rect 10577 92023 10625 92051
rect 10653 92023 10687 92051
rect 10715 92023 10749 92051
rect 10777 92023 10811 92051
rect 10839 92023 10887 92051
rect 10577 91989 10887 92023
rect 10577 91961 10625 91989
rect 10653 91961 10687 91989
rect 10715 91961 10749 91989
rect 10777 91961 10811 91989
rect 10839 91961 10887 91989
rect 10577 83175 10887 91961
rect 10577 83147 10625 83175
rect 10653 83147 10687 83175
rect 10715 83147 10749 83175
rect 10777 83147 10811 83175
rect 10839 83147 10887 83175
rect 10577 83113 10887 83147
rect 10577 83085 10625 83113
rect 10653 83085 10687 83113
rect 10715 83085 10749 83113
rect 10777 83085 10811 83113
rect 10839 83085 10887 83113
rect 10577 83051 10887 83085
rect 10577 83023 10625 83051
rect 10653 83023 10687 83051
rect 10715 83023 10749 83051
rect 10777 83023 10811 83051
rect 10839 83023 10887 83051
rect 10577 82989 10887 83023
rect 10577 82961 10625 82989
rect 10653 82961 10687 82989
rect 10715 82961 10749 82989
rect 10777 82961 10811 82989
rect 10839 82961 10887 82989
rect 10577 74175 10887 82961
rect 10577 74147 10625 74175
rect 10653 74147 10687 74175
rect 10715 74147 10749 74175
rect 10777 74147 10811 74175
rect 10839 74147 10887 74175
rect 10577 74113 10887 74147
rect 10577 74085 10625 74113
rect 10653 74085 10687 74113
rect 10715 74085 10749 74113
rect 10777 74085 10811 74113
rect 10839 74085 10887 74113
rect 10577 74051 10887 74085
rect 10577 74023 10625 74051
rect 10653 74023 10687 74051
rect 10715 74023 10749 74051
rect 10777 74023 10811 74051
rect 10839 74023 10887 74051
rect 10577 73989 10887 74023
rect 10577 73961 10625 73989
rect 10653 73961 10687 73989
rect 10715 73961 10749 73989
rect 10777 73961 10811 73989
rect 10839 73961 10887 73989
rect 10577 65175 10887 73961
rect 10577 65147 10625 65175
rect 10653 65147 10687 65175
rect 10715 65147 10749 65175
rect 10777 65147 10811 65175
rect 10839 65147 10887 65175
rect 10577 65113 10887 65147
rect 10577 65085 10625 65113
rect 10653 65085 10687 65113
rect 10715 65085 10749 65113
rect 10777 65085 10811 65113
rect 10839 65085 10887 65113
rect 10577 65051 10887 65085
rect 10577 65023 10625 65051
rect 10653 65023 10687 65051
rect 10715 65023 10749 65051
rect 10777 65023 10811 65051
rect 10839 65023 10887 65051
rect 10577 64989 10887 65023
rect 10577 64961 10625 64989
rect 10653 64961 10687 64989
rect 10715 64961 10749 64989
rect 10777 64961 10811 64989
rect 10839 64961 10887 64989
rect 10577 56175 10887 64961
rect 10577 56147 10625 56175
rect 10653 56147 10687 56175
rect 10715 56147 10749 56175
rect 10777 56147 10811 56175
rect 10839 56147 10887 56175
rect 10577 56113 10887 56147
rect 10577 56085 10625 56113
rect 10653 56085 10687 56113
rect 10715 56085 10749 56113
rect 10777 56085 10811 56113
rect 10839 56085 10887 56113
rect 10577 56051 10887 56085
rect 10577 56023 10625 56051
rect 10653 56023 10687 56051
rect 10715 56023 10749 56051
rect 10777 56023 10811 56051
rect 10839 56023 10887 56051
rect 10577 55989 10887 56023
rect 10577 55961 10625 55989
rect 10653 55961 10687 55989
rect 10715 55961 10749 55989
rect 10777 55961 10811 55989
rect 10839 55961 10887 55989
rect 10577 47175 10887 55961
rect 10577 47147 10625 47175
rect 10653 47147 10687 47175
rect 10715 47147 10749 47175
rect 10777 47147 10811 47175
rect 10839 47147 10887 47175
rect 10577 47113 10887 47147
rect 10577 47085 10625 47113
rect 10653 47085 10687 47113
rect 10715 47085 10749 47113
rect 10777 47085 10811 47113
rect 10839 47085 10887 47113
rect 10577 47051 10887 47085
rect 10577 47023 10625 47051
rect 10653 47023 10687 47051
rect 10715 47023 10749 47051
rect 10777 47023 10811 47051
rect 10839 47023 10887 47051
rect 10577 46989 10887 47023
rect 10577 46961 10625 46989
rect 10653 46961 10687 46989
rect 10715 46961 10749 46989
rect 10777 46961 10811 46989
rect 10839 46961 10887 46989
rect 10577 38175 10887 46961
rect 10577 38147 10625 38175
rect 10653 38147 10687 38175
rect 10715 38147 10749 38175
rect 10777 38147 10811 38175
rect 10839 38147 10887 38175
rect 10577 38113 10887 38147
rect 10577 38085 10625 38113
rect 10653 38085 10687 38113
rect 10715 38085 10749 38113
rect 10777 38085 10811 38113
rect 10839 38085 10887 38113
rect 10577 38051 10887 38085
rect 10577 38023 10625 38051
rect 10653 38023 10687 38051
rect 10715 38023 10749 38051
rect 10777 38023 10811 38051
rect 10839 38023 10887 38051
rect 10577 37989 10887 38023
rect 10577 37961 10625 37989
rect 10653 37961 10687 37989
rect 10715 37961 10749 37989
rect 10777 37961 10811 37989
rect 10839 37961 10887 37989
rect 10577 29175 10887 37961
rect 10577 29147 10625 29175
rect 10653 29147 10687 29175
rect 10715 29147 10749 29175
rect 10777 29147 10811 29175
rect 10839 29147 10887 29175
rect 10577 29113 10887 29147
rect 10577 29085 10625 29113
rect 10653 29085 10687 29113
rect 10715 29085 10749 29113
rect 10777 29085 10811 29113
rect 10839 29085 10887 29113
rect 10577 29051 10887 29085
rect 10577 29023 10625 29051
rect 10653 29023 10687 29051
rect 10715 29023 10749 29051
rect 10777 29023 10811 29051
rect 10839 29023 10887 29051
rect 10577 28989 10887 29023
rect 10577 28961 10625 28989
rect 10653 28961 10687 28989
rect 10715 28961 10749 28989
rect 10777 28961 10811 28989
rect 10839 28961 10887 28989
rect 10577 20175 10887 28961
rect 10577 20147 10625 20175
rect 10653 20147 10687 20175
rect 10715 20147 10749 20175
rect 10777 20147 10811 20175
rect 10839 20147 10887 20175
rect 10577 20113 10887 20147
rect 10577 20085 10625 20113
rect 10653 20085 10687 20113
rect 10715 20085 10749 20113
rect 10777 20085 10811 20113
rect 10839 20085 10887 20113
rect 10577 20051 10887 20085
rect 10577 20023 10625 20051
rect 10653 20023 10687 20051
rect 10715 20023 10749 20051
rect 10777 20023 10811 20051
rect 10839 20023 10887 20051
rect 10577 19989 10887 20023
rect 10577 19961 10625 19989
rect 10653 19961 10687 19989
rect 10715 19961 10749 19989
rect 10777 19961 10811 19989
rect 10839 19961 10887 19989
rect 10577 11175 10887 19961
rect 10577 11147 10625 11175
rect 10653 11147 10687 11175
rect 10715 11147 10749 11175
rect 10777 11147 10811 11175
rect 10839 11147 10887 11175
rect 10577 11113 10887 11147
rect 10577 11085 10625 11113
rect 10653 11085 10687 11113
rect 10715 11085 10749 11113
rect 10777 11085 10811 11113
rect 10839 11085 10887 11113
rect 10577 11051 10887 11085
rect 10577 11023 10625 11051
rect 10653 11023 10687 11051
rect 10715 11023 10749 11051
rect 10777 11023 10811 11051
rect 10839 11023 10887 11051
rect 10577 10989 10887 11023
rect 10577 10961 10625 10989
rect 10653 10961 10687 10989
rect 10715 10961 10749 10989
rect 10777 10961 10811 10989
rect 10839 10961 10887 10989
rect 10577 2175 10887 10961
rect 10577 2147 10625 2175
rect 10653 2147 10687 2175
rect 10715 2147 10749 2175
rect 10777 2147 10811 2175
rect 10839 2147 10887 2175
rect 10577 2113 10887 2147
rect 10577 2085 10625 2113
rect 10653 2085 10687 2113
rect 10715 2085 10749 2113
rect 10777 2085 10811 2113
rect 10839 2085 10887 2113
rect 10577 2051 10887 2085
rect 10577 2023 10625 2051
rect 10653 2023 10687 2051
rect 10715 2023 10749 2051
rect 10777 2023 10811 2051
rect 10839 2023 10887 2051
rect 10577 1989 10887 2023
rect 10577 1961 10625 1989
rect 10653 1961 10687 1989
rect 10715 1961 10749 1989
rect 10777 1961 10811 1989
rect 10839 1961 10887 1989
rect 10577 -80 10887 1961
rect 10577 -108 10625 -80
rect 10653 -108 10687 -80
rect 10715 -108 10749 -80
rect 10777 -108 10811 -80
rect 10839 -108 10887 -80
rect 10577 -142 10887 -108
rect 10577 -170 10625 -142
rect 10653 -170 10687 -142
rect 10715 -170 10749 -142
rect 10777 -170 10811 -142
rect 10839 -170 10887 -142
rect 10577 -204 10887 -170
rect 10577 -232 10625 -204
rect 10653 -232 10687 -204
rect 10715 -232 10749 -204
rect 10777 -232 10811 -204
rect 10839 -232 10887 -204
rect 10577 -266 10887 -232
rect 10577 -294 10625 -266
rect 10653 -294 10687 -266
rect 10715 -294 10749 -266
rect 10777 -294 10811 -266
rect 10839 -294 10887 -266
rect 10577 -822 10887 -294
rect 12437 299086 12747 299134
rect 12437 299058 12485 299086
rect 12513 299058 12547 299086
rect 12575 299058 12609 299086
rect 12637 299058 12671 299086
rect 12699 299058 12747 299086
rect 12437 299024 12747 299058
rect 12437 298996 12485 299024
rect 12513 298996 12547 299024
rect 12575 298996 12609 299024
rect 12637 298996 12671 299024
rect 12699 298996 12747 299024
rect 12437 298962 12747 298996
rect 12437 298934 12485 298962
rect 12513 298934 12547 298962
rect 12575 298934 12609 298962
rect 12637 298934 12671 298962
rect 12699 298934 12747 298962
rect 12437 298900 12747 298934
rect 12437 298872 12485 298900
rect 12513 298872 12547 298900
rect 12575 298872 12609 298900
rect 12637 298872 12671 298900
rect 12699 298872 12747 298900
rect 12437 293175 12747 298872
rect 12437 293147 12485 293175
rect 12513 293147 12547 293175
rect 12575 293147 12609 293175
rect 12637 293147 12671 293175
rect 12699 293147 12747 293175
rect 12437 293113 12747 293147
rect 12437 293085 12485 293113
rect 12513 293085 12547 293113
rect 12575 293085 12609 293113
rect 12637 293085 12671 293113
rect 12699 293085 12747 293113
rect 12437 293051 12747 293085
rect 12437 293023 12485 293051
rect 12513 293023 12547 293051
rect 12575 293023 12609 293051
rect 12637 293023 12671 293051
rect 12699 293023 12747 293051
rect 12437 292989 12747 293023
rect 12437 292961 12485 292989
rect 12513 292961 12547 292989
rect 12575 292961 12609 292989
rect 12637 292961 12671 292989
rect 12699 292961 12747 292989
rect 12437 284175 12747 292961
rect 12437 284147 12485 284175
rect 12513 284147 12547 284175
rect 12575 284147 12609 284175
rect 12637 284147 12671 284175
rect 12699 284147 12747 284175
rect 12437 284113 12747 284147
rect 12437 284085 12485 284113
rect 12513 284085 12547 284113
rect 12575 284085 12609 284113
rect 12637 284085 12671 284113
rect 12699 284085 12747 284113
rect 12437 284051 12747 284085
rect 12437 284023 12485 284051
rect 12513 284023 12547 284051
rect 12575 284023 12609 284051
rect 12637 284023 12671 284051
rect 12699 284023 12747 284051
rect 12437 283989 12747 284023
rect 12437 283961 12485 283989
rect 12513 283961 12547 283989
rect 12575 283961 12609 283989
rect 12637 283961 12671 283989
rect 12699 283961 12747 283989
rect 12437 275175 12747 283961
rect 12437 275147 12485 275175
rect 12513 275147 12547 275175
rect 12575 275147 12609 275175
rect 12637 275147 12671 275175
rect 12699 275147 12747 275175
rect 12437 275113 12747 275147
rect 12437 275085 12485 275113
rect 12513 275085 12547 275113
rect 12575 275085 12609 275113
rect 12637 275085 12671 275113
rect 12699 275085 12747 275113
rect 12437 275051 12747 275085
rect 12437 275023 12485 275051
rect 12513 275023 12547 275051
rect 12575 275023 12609 275051
rect 12637 275023 12671 275051
rect 12699 275023 12747 275051
rect 12437 274989 12747 275023
rect 12437 274961 12485 274989
rect 12513 274961 12547 274989
rect 12575 274961 12609 274989
rect 12637 274961 12671 274989
rect 12699 274961 12747 274989
rect 12437 266175 12747 274961
rect 12437 266147 12485 266175
rect 12513 266147 12547 266175
rect 12575 266147 12609 266175
rect 12637 266147 12671 266175
rect 12699 266147 12747 266175
rect 12437 266113 12747 266147
rect 12437 266085 12485 266113
rect 12513 266085 12547 266113
rect 12575 266085 12609 266113
rect 12637 266085 12671 266113
rect 12699 266085 12747 266113
rect 12437 266051 12747 266085
rect 12437 266023 12485 266051
rect 12513 266023 12547 266051
rect 12575 266023 12609 266051
rect 12637 266023 12671 266051
rect 12699 266023 12747 266051
rect 12437 265989 12747 266023
rect 12437 265961 12485 265989
rect 12513 265961 12547 265989
rect 12575 265961 12609 265989
rect 12637 265961 12671 265989
rect 12699 265961 12747 265989
rect 12437 257175 12747 265961
rect 12437 257147 12485 257175
rect 12513 257147 12547 257175
rect 12575 257147 12609 257175
rect 12637 257147 12671 257175
rect 12699 257147 12747 257175
rect 12437 257113 12747 257147
rect 12437 257085 12485 257113
rect 12513 257085 12547 257113
rect 12575 257085 12609 257113
rect 12637 257085 12671 257113
rect 12699 257085 12747 257113
rect 12437 257051 12747 257085
rect 12437 257023 12485 257051
rect 12513 257023 12547 257051
rect 12575 257023 12609 257051
rect 12637 257023 12671 257051
rect 12699 257023 12747 257051
rect 12437 256989 12747 257023
rect 12437 256961 12485 256989
rect 12513 256961 12547 256989
rect 12575 256961 12609 256989
rect 12637 256961 12671 256989
rect 12699 256961 12747 256989
rect 12437 248175 12747 256961
rect 12437 248147 12485 248175
rect 12513 248147 12547 248175
rect 12575 248147 12609 248175
rect 12637 248147 12671 248175
rect 12699 248147 12747 248175
rect 12437 248113 12747 248147
rect 12437 248085 12485 248113
rect 12513 248085 12547 248113
rect 12575 248085 12609 248113
rect 12637 248085 12671 248113
rect 12699 248085 12747 248113
rect 12437 248051 12747 248085
rect 12437 248023 12485 248051
rect 12513 248023 12547 248051
rect 12575 248023 12609 248051
rect 12637 248023 12671 248051
rect 12699 248023 12747 248051
rect 12437 247989 12747 248023
rect 12437 247961 12485 247989
rect 12513 247961 12547 247989
rect 12575 247961 12609 247989
rect 12637 247961 12671 247989
rect 12699 247961 12747 247989
rect 12437 239175 12747 247961
rect 12437 239147 12485 239175
rect 12513 239147 12547 239175
rect 12575 239147 12609 239175
rect 12637 239147 12671 239175
rect 12699 239147 12747 239175
rect 12437 239113 12747 239147
rect 12437 239085 12485 239113
rect 12513 239085 12547 239113
rect 12575 239085 12609 239113
rect 12637 239085 12671 239113
rect 12699 239085 12747 239113
rect 12437 239051 12747 239085
rect 12437 239023 12485 239051
rect 12513 239023 12547 239051
rect 12575 239023 12609 239051
rect 12637 239023 12671 239051
rect 12699 239023 12747 239051
rect 12437 238989 12747 239023
rect 12437 238961 12485 238989
rect 12513 238961 12547 238989
rect 12575 238961 12609 238989
rect 12637 238961 12671 238989
rect 12699 238961 12747 238989
rect 12437 230175 12747 238961
rect 12437 230147 12485 230175
rect 12513 230147 12547 230175
rect 12575 230147 12609 230175
rect 12637 230147 12671 230175
rect 12699 230147 12747 230175
rect 12437 230113 12747 230147
rect 12437 230085 12485 230113
rect 12513 230085 12547 230113
rect 12575 230085 12609 230113
rect 12637 230085 12671 230113
rect 12699 230085 12747 230113
rect 12437 230051 12747 230085
rect 12437 230023 12485 230051
rect 12513 230023 12547 230051
rect 12575 230023 12609 230051
rect 12637 230023 12671 230051
rect 12699 230023 12747 230051
rect 12437 229989 12747 230023
rect 12437 229961 12485 229989
rect 12513 229961 12547 229989
rect 12575 229961 12609 229989
rect 12637 229961 12671 229989
rect 12699 229961 12747 229989
rect 12437 221175 12747 229961
rect 12437 221147 12485 221175
rect 12513 221147 12547 221175
rect 12575 221147 12609 221175
rect 12637 221147 12671 221175
rect 12699 221147 12747 221175
rect 12437 221113 12747 221147
rect 12437 221085 12485 221113
rect 12513 221085 12547 221113
rect 12575 221085 12609 221113
rect 12637 221085 12671 221113
rect 12699 221085 12747 221113
rect 12437 221051 12747 221085
rect 12437 221023 12485 221051
rect 12513 221023 12547 221051
rect 12575 221023 12609 221051
rect 12637 221023 12671 221051
rect 12699 221023 12747 221051
rect 12437 220989 12747 221023
rect 12437 220961 12485 220989
rect 12513 220961 12547 220989
rect 12575 220961 12609 220989
rect 12637 220961 12671 220989
rect 12699 220961 12747 220989
rect 12437 212175 12747 220961
rect 12437 212147 12485 212175
rect 12513 212147 12547 212175
rect 12575 212147 12609 212175
rect 12637 212147 12671 212175
rect 12699 212147 12747 212175
rect 12437 212113 12747 212147
rect 12437 212085 12485 212113
rect 12513 212085 12547 212113
rect 12575 212085 12609 212113
rect 12637 212085 12671 212113
rect 12699 212085 12747 212113
rect 12437 212051 12747 212085
rect 12437 212023 12485 212051
rect 12513 212023 12547 212051
rect 12575 212023 12609 212051
rect 12637 212023 12671 212051
rect 12699 212023 12747 212051
rect 12437 211989 12747 212023
rect 12437 211961 12485 211989
rect 12513 211961 12547 211989
rect 12575 211961 12609 211989
rect 12637 211961 12671 211989
rect 12699 211961 12747 211989
rect 12437 203175 12747 211961
rect 12437 203147 12485 203175
rect 12513 203147 12547 203175
rect 12575 203147 12609 203175
rect 12637 203147 12671 203175
rect 12699 203147 12747 203175
rect 12437 203113 12747 203147
rect 12437 203085 12485 203113
rect 12513 203085 12547 203113
rect 12575 203085 12609 203113
rect 12637 203085 12671 203113
rect 12699 203085 12747 203113
rect 12437 203051 12747 203085
rect 12437 203023 12485 203051
rect 12513 203023 12547 203051
rect 12575 203023 12609 203051
rect 12637 203023 12671 203051
rect 12699 203023 12747 203051
rect 12437 202989 12747 203023
rect 12437 202961 12485 202989
rect 12513 202961 12547 202989
rect 12575 202961 12609 202989
rect 12637 202961 12671 202989
rect 12699 202961 12747 202989
rect 12437 194175 12747 202961
rect 12437 194147 12485 194175
rect 12513 194147 12547 194175
rect 12575 194147 12609 194175
rect 12637 194147 12671 194175
rect 12699 194147 12747 194175
rect 12437 194113 12747 194147
rect 12437 194085 12485 194113
rect 12513 194085 12547 194113
rect 12575 194085 12609 194113
rect 12637 194085 12671 194113
rect 12699 194085 12747 194113
rect 12437 194051 12747 194085
rect 12437 194023 12485 194051
rect 12513 194023 12547 194051
rect 12575 194023 12609 194051
rect 12637 194023 12671 194051
rect 12699 194023 12747 194051
rect 12437 193989 12747 194023
rect 12437 193961 12485 193989
rect 12513 193961 12547 193989
rect 12575 193961 12609 193989
rect 12637 193961 12671 193989
rect 12699 193961 12747 193989
rect 12437 185175 12747 193961
rect 12437 185147 12485 185175
rect 12513 185147 12547 185175
rect 12575 185147 12609 185175
rect 12637 185147 12671 185175
rect 12699 185147 12747 185175
rect 12437 185113 12747 185147
rect 12437 185085 12485 185113
rect 12513 185085 12547 185113
rect 12575 185085 12609 185113
rect 12637 185085 12671 185113
rect 12699 185085 12747 185113
rect 12437 185051 12747 185085
rect 12437 185023 12485 185051
rect 12513 185023 12547 185051
rect 12575 185023 12609 185051
rect 12637 185023 12671 185051
rect 12699 185023 12747 185051
rect 12437 184989 12747 185023
rect 12437 184961 12485 184989
rect 12513 184961 12547 184989
rect 12575 184961 12609 184989
rect 12637 184961 12671 184989
rect 12699 184961 12747 184989
rect 12437 176175 12747 184961
rect 12437 176147 12485 176175
rect 12513 176147 12547 176175
rect 12575 176147 12609 176175
rect 12637 176147 12671 176175
rect 12699 176147 12747 176175
rect 12437 176113 12747 176147
rect 12437 176085 12485 176113
rect 12513 176085 12547 176113
rect 12575 176085 12609 176113
rect 12637 176085 12671 176113
rect 12699 176085 12747 176113
rect 12437 176051 12747 176085
rect 12437 176023 12485 176051
rect 12513 176023 12547 176051
rect 12575 176023 12609 176051
rect 12637 176023 12671 176051
rect 12699 176023 12747 176051
rect 12437 175989 12747 176023
rect 12437 175961 12485 175989
rect 12513 175961 12547 175989
rect 12575 175961 12609 175989
rect 12637 175961 12671 175989
rect 12699 175961 12747 175989
rect 12437 167175 12747 175961
rect 12437 167147 12485 167175
rect 12513 167147 12547 167175
rect 12575 167147 12609 167175
rect 12637 167147 12671 167175
rect 12699 167147 12747 167175
rect 12437 167113 12747 167147
rect 12437 167085 12485 167113
rect 12513 167085 12547 167113
rect 12575 167085 12609 167113
rect 12637 167085 12671 167113
rect 12699 167085 12747 167113
rect 12437 167051 12747 167085
rect 12437 167023 12485 167051
rect 12513 167023 12547 167051
rect 12575 167023 12609 167051
rect 12637 167023 12671 167051
rect 12699 167023 12747 167051
rect 12437 166989 12747 167023
rect 12437 166961 12485 166989
rect 12513 166961 12547 166989
rect 12575 166961 12609 166989
rect 12637 166961 12671 166989
rect 12699 166961 12747 166989
rect 12437 158175 12747 166961
rect 12437 158147 12485 158175
rect 12513 158147 12547 158175
rect 12575 158147 12609 158175
rect 12637 158147 12671 158175
rect 12699 158147 12747 158175
rect 12437 158113 12747 158147
rect 12437 158085 12485 158113
rect 12513 158085 12547 158113
rect 12575 158085 12609 158113
rect 12637 158085 12671 158113
rect 12699 158085 12747 158113
rect 12437 158051 12747 158085
rect 12437 158023 12485 158051
rect 12513 158023 12547 158051
rect 12575 158023 12609 158051
rect 12637 158023 12671 158051
rect 12699 158023 12747 158051
rect 12437 157989 12747 158023
rect 12437 157961 12485 157989
rect 12513 157961 12547 157989
rect 12575 157961 12609 157989
rect 12637 157961 12671 157989
rect 12699 157961 12747 157989
rect 12437 149175 12747 157961
rect 12437 149147 12485 149175
rect 12513 149147 12547 149175
rect 12575 149147 12609 149175
rect 12637 149147 12671 149175
rect 12699 149147 12747 149175
rect 12437 149113 12747 149147
rect 12437 149085 12485 149113
rect 12513 149085 12547 149113
rect 12575 149085 12609 149113
rect 12637 149085 12671 149113
rect 12699 149085 12747 149113
rect 12437 149051 12747 149085
rect 12437 149023 12485 149051
rect 12513 149023 12547 149051
rect 12575 149023 12609 149051
rect 12637 149023 12671 149051
rect 12699 149023 12747 149051
rect 12437 148989 12747 149023
rect 12437 148961 12485 148989
rect 12513 148961 12547 148989
rect 12575 148961 12609 148989
rect 12637 148961 12671 148989
rect 12699 148961 12747 148989
rect 12437 140175 12747 148961
rect 12437 140147 12485 140175
rect 12513 140147 12547 140175
rect 12575 140147 12609 140175
rect 12637 140147 12671 140175
rect 12699 140147 12747 140175
rect 12437 140113 12747 140147
rect 12437 140085 12485 140113
rect 12513 140085 12547 140113
rect 12575 140085 12609 140113
rect 12637 140085 12671 140113
rect 12699 140085 12747 140113
rect 12437 140051 12747 140085
rect 12437 140023 12485 140051
rect 12513 140023 12547 140051
rect 12575 140023 12609 140051
rect 12637 140023 12671 140051
rect 12699 140023 12747 140051
rect 12437 139989 12747 140023
rect 12437 139961 12485 139989
rect 12513 139961 12547 139989
rect 12575 139961 12609 139989
rect 12637 139961 12671 139989
rect 12699 139961 12747 139989
rect 12437 131175 12747 139961
rect 12437 131147 12485 131175
rect 12513 131147 12547 131175
rect 12575 131147 12609 131175
rect 12637 131147 12671 131175
rect 12699 131147 12747 131175
rect 12437 131113 12747 131147
rect 12437 131085 12485 131113
rect 12513 131085 12547 131113
rect 12575 131085 12609 131113
rect 12637 131085 12671 131113
rect 12699 131085 12747 131113
rect 12437 131051 12747 131085
rect 12437 131023 12485 131051
rect 12513 131023 12547 131051
rect 12575 131023 12609 131051
rect 12637 131023 12671 131051
rect 12699 131023 12747 131051
rect 12437 130989 12747 131023
rect 12437 130961 12485 130989
rect 12513 130961 12547 130989
rect 12575 130961 12609 130989
rect 12637 130961 12671 130989
rect 12699 130961 12747 130989
rect 12437 122175 12747 130961
rect 12437 122147 12485 122175
rect 12513 122147 12547 122175
rect 12575 122147 12609 122175
rect 12637 122147 12671 122175
rect 12699 122147 12747 122175
rect 12437 122113 12747 122147
rect 12437 122085 12485 122113
rect 12513 122085 12547 122113
rect 12575 122085 12609 122113
rect 12637 122085 12671 122113
rect 12699 122085 12747 122113
rect 12437 122051 12747 122085
rect 12437 122023 12485 122051
rect 12513 122023 12547 122051
rect 12575 122023 12609 122051
rect 12637 122023 12671 122051
rect 12699 122023 12747 122051
rect 12437 121989 12747 122023
rect 12437 121961 12485 121989
rect 12513 121961 12547 121989
rect 12575 121961 12609 121989
rect 12637 121961 12671 121989
rect 12699 121961 12747 121989
rect 12437 113175 12747 121961
rect 12437 113147 12485 113175
rect 12513 113147 12547 113175
rect 12575 113147 12609 113175
rect 12637 113147 12671 113175
rect 12699 113147 12747 113175
rect 12437 113113 12747 113147
rect 12437 113085 12485 113113
rect 12513 113085 12547 113113
rect 12575 113085 12609 113113
rect 12637 113085 12671 113113
rect 12699 113085 12747 113113
rect 12437 113051 12747 113085
rect 12437 113023 12485 113051
rect 12513 113023 12547 113051
rect 12575 113023 12609 113051
rect 12637 113023 12671 113051
rect 12699 113023 12747 113051
rect 12437 112989 12747 113023
rect 12437 112961 12485 112989
rect 12513 112961 12547 112989
rect 12575 112961 12609 112989
rect 12637 112961 12671 112989
rect 12699 112961 12747 112989
rect 12437 104175 12747 112961
rect 12437 104147 12485 104175
rect 12513 104147 12547 104175
rect 12575 104147 12609 104175
rect 12637 104147 12671 104175
rect 12699 104147 12747 104175
rect 12437 104113 12747 104147
rect 12437 104085 12485 104113
rect 12513 104085 12547 104113
rect 12575 104085 12609 104113
rect 12637 104085 12671 104113
rect 12699 104085 12747 104113
rect 12437 104051 12747 104085
rect 12437 104023 12485 104051
rect 12513 104023 12547 104051
rect 12575 104023 12609 104051
rect 12637 104023 12671 104051
rect 12699 104023 12747 104051
rect 12437 103989 12747 104023
rect 12437 103961 12485 103989
rect 12513 103961 12547 103989
rect 12575 103961 12609 103989
rect 12637 103961 12671 103989
rect 12699 103961 12747 103989
rect 12437 95175 12747 103961
rect 12437 95147 12485 95175
rect 12513 95147 12547 95175
rect 12575 95147 12609 95175
rect 12637 95147 12671 95175
rect 12699 95147 12747 95175
rect 12437 95113 12747 95147
rect 12437 95085 12485 95113
rect 12513 95085 12547 95113
rect 12575 95085 12609 95113
rect 12637 95085 12671 95113
rect 12699 95085 12747 95113
rect 12437 95051 12747 95085
rect 12437 95023 12485 95051
rect 12513 95023 12547 95051
rect 12575 95023 12609 95051
rect 12637 95023 12671 95051
rect 12699 95023 12747 95051
rect 12437 94989 12747 95023
rect 12437 94961 12485 94989
rect 12513 94961 12547 94989
rect 12575 94961 12609 94989
rect 12637 94961 12671 94989
rect 12699 94961 12747 94989
rect 12437 86175 12747 94961
rect 12437 86147 12485 86175
rect 12513 86147 12547 86175
rect 12575 86147 12609 86175
rect 12637 86147 12671 86175
rect 12699 86147 12747 86175
rect 12437 86113 12747 86147
rect 12437 86085 12485 86113
rect 12513 86085 12547 86113
rect 12575 86085 12609 86113
rect 12637 86085 12671 86113
rect 12699 86085 12747 86113
rect 12437 86051 12747 86085
rect 12437 86023 12485 86051
rect 12513 86023 12547 86051
rect 12575 86023 12609 86051
rect 12637 86023 12671 86051
rect 12699 86023 12747 86051
rect 12437 85989 12747 86023
rect 12437 85961 12485 85989
rect 12513 85961 12547 85989
rect 12575 85961 12609 85989
rect 12637 85961 12671 85989
rect 12699 85961 12747 85989
rect 12437 77175 12747 85961
rect 12437 77147 12485 77175
rect 12513 77147 12547 77175
rect 12575 77147 12609 77175
rect 12637 77147 12671 77175
rect 12699 77147 12747 77175
rect 12437 77113 12747 77147
rect 12437 77085 12485 77113
rect 12513 77085 12547 77113
rect 12575 77085 12609 77113
rect 12637 77085 12671 77113
rect 12699 77085 12747 77113
rect 12437 77051 12747 77085
rect 12437 77023 12485 77051
rect 12513 77023 12547 77051
rect 12575 77023 12609 77051
rect 12637 77023 12671 77051
rect 12699 77023 12747 77051
rect 12437 76989 12747 77023
rect 12437 76961 12485 76989
rect 12513 76961 12547 76989
rect 12575 76961 12609 76989
rect 12637 76961 12671 76989
rect 12699 76961 12747 76989
rect 12437 68175 12747 76961
rect 12437 68147 12485 68175
rect 12513 68147 12547 68175
rect 12575 68147 12609 68175
rect 12637 68147 12671 68175
rect 12699 68147 12747 68175
rect 12437 68113 12747 68147
rect 12437 68085 12485 68113
rect 12513 68085 12547 68113
rect 12575 68085 12609 68113
rect 12637 68085 12671 68113
rect 12699 68085 12747 68113
rect 12437 68051 12747 68085
rect 12437 68023 12485 68051
rect 12513 68023 12547 68051
rect 12575 68023 12609 68051
rect 12637 68023 12671 68051
rect 12699 68023 12747 68051
rect 12437 67989 12747 68023
rect 12437 67961 12485 67989
rect 12513 67961 12547 67989
rect 12575 67961 12609 67989
rect 12637 67961 12671 67989
rect 12699 67961 12747 67989
rect 12437 59175 12747 67961
rect 12437 59147 12485 59175
rect 12513 59147 12547 59175
rect 12575 59147 12609 59175
rect 12637 59147 12671 59175
rect 12699 59147 12747 59175
rect 12437 59113 12747 59147
rect 12437 59085 12485 59113
rect 12513 59085 12547 59113
rect 12575 59085 12609 59113
rect 12637 59085 12671 59113
rect 12699 59085 12747 59113
rect 12437 59051 12747 59085
rect 12437 59023 12485 59051
rect 12513 59023 12547 59051
rect 12575 59023 12609 59051
rect 12637 59023 12671 59051
rect 12699 59023 12747 59051
rect 12437 58989 12747 59023
rect 12437 58961 12485 58989
rect 12513 58961 12547 58989
rect 12575 58961 12609 58989
rect 12637 58961 12671 58989
rect 12699 58961 12747 58989
rect 12437 50175 12747 58961
rect 12437 50147 12485 50175
rect 12513 50147 12547 50175
rect 12575 50147 12609 50175
rect 12637 50147 12671 50175
rect 12699 50147 12747 50175
rect 12437 50113 12747 50147
rect 12437 50085 12485 50113
rect 12513 50085 12547 50113
rect 12575 50085 12609 50113
rect 12637 50085 12671 50113
rect 12699 50085 12747 50113
rect 12437 50051 12747 50085
rect 12437 50023 12485 50051
rect 12513 50023 12547 50051
rect 12575 50023 12609 50051
rect 12637 50023 12671 50051
rect 12699 50023 12747 50051
rect 12437 49989 12747 50023
rect 12437 49961 12485 49989
rect 12513 49961 12547 49989
rect 12575 49961 12609 49989
rect 12637 49961 12671 49989
rect 12699 49961 12747 49989
rect 12437 41175 12747 49961
rect 12437 41147 12485 41175
rect 12513 41147 12547 41175
rect 12575 41147 12609 41175
rect 12637 41147 12671 41175
rect 12699 41147 12747 41175
rect 12437 41113 12747 41147
rect 12437 41085 12485 41113
rect 12513 41085 12547 41113
rect 12575 41085 12609 41113
rect 12637 41085 12671 41113
rect 12699 41085 12747 41113
rect 12437 41051 12747 41085
rect 12437 41023 12485 41051
rect 12513 41023 12547 41051
rect 12575 41023 12609 41051
rect 12637 41023 12671 41051
rect 12699 41023 12747 41051
rect 12437 40989 12747 41023
rect 12437 40961 12485 40989
rect 12513 40961 12547 40989
rect 12575 40961 12609 40989
rect 12637 40961 12671 40989
rect 12699 40961 12747 40989
rect 12437 32175 12747 40961
rect 12437 32147 12485 32175
rect 12513 32147 12547 32175
rect 12575 32147 12609 32175
rect 12637 32147 12671 32175
rect 12699 32147 12747 32175
rect 12437 32113 12747 32147
rect 12437 32085 12485 32113
rect 12513 32085 12547 32113
rect 12575 32085 12609 32113
rect 12637 32085 12671 32113
rect 12699 32085 12747 32113
rect 12437 32051 12747 32085
rect 12437 32023 12485 32051
rect 12513 32023 12547 32051
rect 12575 32023 12609 32051
rect 12637 32023 12671 32051
rect 12699 32023 12747 32051
rect 12437 31989 12747 32023
rect 12437 31961 12485 31989
rect 12513 31961 12547 31989
rect 12575 31961 12609 31989
rect 12637 31961 12671 31989
rect 12699 31961 12747 31989
rect 12437 23175 12747 31961
rect 12437 23147 12485 23175
rect 12513 23147 12547 23175
rect 12575 23147 12609 23175
rect 12637 23147 12671 23175
rect 12699 23147 12747 23175
rect 12437 23113 12747 23147
rect 12437 23085 12485 23113
rect 12513 23085 12547 23113
rect 12575 23085 12609 23113
rect 12637 23085 12671 23113
rect 12699 23085 12747 23113
rect 12437 23051 12747 23085
rect 12437 23023 12485 23051
rect 12513 23023 12547 23051
rect 12575 23023 12609 23051
rect 12637 23023 12671 23051
rect 12699 23023 12747 23051
rect 12437 22989 12747 23023
rect 12437 22961 12485 22989
rect 12513 22961 12547 22989
rect 12575 22961 12609 22989
rect 12637 22961 12671 22989
rect 12699 22961 12747 22989
rect 12437 14175 12747 22961
rect 12437 14147 12485 14175
rect 12513 14147 12547 14175
rect 12575 14147 12609 14175
rect 12637 14147 12671 14175
rect 12699 14147 12747 14175
rect 12437 14113 12747 14147
rect 12437 14085 12485 14113
rect 12513 14085 12547 14113
rect 12575 14085 12609 14113
rect 12637 14085 12671 14113
rect 12699 14085 12747 14113
rect 12437 14051 12747 14085
rect 12437 14023 12485 14051
rect 12513 14023 12547 14051
rect 12575 14023 12609 14051
rect 12637 14023 12671 14051
rect 12699 14023 12747 14051
rect 12437 13989 12747 14023
rect 12437 13961 12485 13989
rect 12513 13961 12547 13989
rect 12575 13961 12609 13989
rect 12637 13961 12671 13989
rect 12699 13961 12747 13989
rect 12437 5175 12747 13961
rect 12437 5147 12485 5175
rect 12513 5147 12547 5175
rect 12575 5147 12609 5175
rect 12637 5147 12671 5175
rect 12699 5147 12747 5175
rect 12437 5113 12747 5147
rect 12437 5085 12485 5113
rect 12513 5085 12547 5113
rect 12575 5085 12609 5113
rect 12637 5085 12671 5113
rect 12699 5085 12747 5113
rect 12437 5051 12747 5085
rect 12437 5023 12485 5051
rect 12513 5023 12547 5051
rect 12575 5023 12609 5051
rect 12637 5023 12671 5051
rect 12699 5023 12747 5051
rect 12437 4989 12747 5023
rect 12437 4961 12485 4989
rect 12513 4961 12547 4989
rect 12575 4961 12609 4989
rect 12637 4961 12671 4989
rect 12699 4961 12747 4989
rect 12437 -560 12747 4961
rect 12437 -588 12485 -560
rect 12513 -588 12547 -560
rect 12575 -588 12609 -560
rect 12637 -588 12671 -560
rect 12699 -588 12747 -560
rect 12437 -622 12747 -588
rect 12437 -650 12485 -622
rect 12513 -650 12547 -622
rect 12575 -650 12609 -622
rect 12637 -650 12671 -622
rect 12699 -650 12747 -622
rect 12437 -684 12747 -650
rect 12437 -712 12485 -684
rect 12513 -712 12547 -684
rect 12575 -712 12609 -684
rect 12637 -712 12671 -684
rect 12699 -712 12747 -684
rect 12437 -746 12747 -712
rect 12437 -774 12485 -746
rect 12513 -774 12547 -746
rect 12575 -774 12609 -746
rect 12637 -774 12671 -746
rect 12699 -774 12747 -746
rect 12437 -822 12747 -774
rect 19577 298606 19887 299134
rect 19577 298578 19625 298606
rect 19653 298578 19687 298606
rect 19715 298578 19749 298606
rect 19777 298578 19811 298606
rect 19839 298578 19887 298606
rect 19577 298544 19887 298578
rect 19577 298516 19625 298544
rect 19653 298516 19687 298544
rect 19715 298516 19749 298544
rect 19777 298516 19811 298544
rect 19839 298516 19887 298544
rect 19577 298482 19887 298516
rect 19577 298454 19625 298482
rect 19653 298454 19687 298482
rect 19715 298454 19749 298482
rect 19777 298454 19811 298482
rect 19839 298454 19887 298482
rect 19577 298420 19887 298454
rect 19577 298392 19625 298420
rect 19653 298392 19687 298420
rect 19715 298392 19749 298420
rect 19777 298392 19811 298420
rect 19839 298392 19887 298420
rect 19577 290175 19887 298392
rect 19577 290147 19625 290175
rect 19653 290147 19687 290175
rect 19715 290147 19749 290175
rect 19777 290147 19811 290175
rect 19839 290147 19887 290175
rect 19577 290113 19887 290147
rect 19577 290085 19625 290113
rect 19653 290085 19687 290113
rect 19715 290085 19749 290113
rect 19777 290085 19811 290113
rect 19839 290085 19887 290113
rect 19577 290051 19887 290085
rect 19577 290023 19625 290051
rect 19653 290023 19687 290051
rect 19715 290023 19749 290051
rect 19777 290023 19811 290051
rect 19839 290023 19887 290051
rect 19577 289989 19887 290023
rect 19577 289961 19625 289989
rect 19653 289961 19687 289989
rect 19715 289961 19749 289989
rect 19777 289961 19811 289989
rect 19839 289961 19887 289989
rect 19577 281175 19887 289961
rect 19577 281147 19625 281175
rect 19653 281147 19687 281175
rect 19715 281147 19749 281175
rect 19777 281147 19811 281175
rect 19839 281147 19887 281175
rect 19577 281113 19887 281147
rect 19577 281085 19625 281113
rect 19653 281085 19687 281113
rect 19715 281085 19749 281113
rect 19777 281085 19811 281113
rect 19839 281085 19887 281113
rect 19577 281051 19887 281085
rect 19577 281023 19625 281051
rect 19653 281023 19687 281051
rect 19715 281023 19749 281051
rect 19777 281023 19811 281051
rect 19839 281023 19887 281051
rect 19577 280989 19887 281023
rect 19577 280961 19625 280989
rect 19653 280961 19687 280989
rect 19715 280961 19749 280989
rect 19777 280961 19811 280989
rect 19839 280961 19887 280989
rect 19577 272175 19887 280961
rect 19577 272147 19625 272175
rect 19653 272147 19687 272175
rect 19715 272147 19749 272175
rect 19777 272147 19811 272175
rect 19839 272147 19887 272175
rect 19577 272113 19887 272147
rect 19577 272085 19625 272113
rect 19653 272085 19687 272113
rect 19715 272085 19749 272113
rect 19777 272085 19811 272113
rect 19839 272085 19887 272113
rect 19577 272051 19887 272085
rect 19577 272023 19625 272051
rect 19653 272023 19687 272051
rect 19715 272023 19749 272051
rect 19777 272023 19811 272051
rect 19839 272023 19887 272051
rect 19577 271989 19887 272023
rect 19577 271961 19625 271989
rect 19653 271961 19687 271989
rect 19715 271961 19749 271989
rect 19777 271961 19811 271989
rect 19839 271961 19887 271989
rect 19577 263175 19887 271961
rect 19577 263147 19625 263175
rect 19653 263147 19687 263175
rect 19715 263147 19749 263175
rect 19777 263147 19811 263175
rect 19839 263147 19887 263175
rect 19577 263113 19887 263147
rect 19577 263085 19625 263113
rect 19653 263085 19687 263113
rect 19715 263085 19749 263113
rect 19777 263085 19811 263113
rect 19839 263085 19887 263113
rect 19577 263051 19887 263085
rect 19577 263023 19625 263051
rect 19653 263023 19687 263051
rect 19715 263023 19749 263051
rect 19777 263023 19811 263051
rect 19839 263023 19887 263051
rect 19577 262989 19887 263023
rect 19577 262961 19625 262989
rect 19653 262961 19687 262989
rect 19715 262961 19749 262989
rect 19777 262961 19811 262989
rect 19839 262961 19887 262989
rect 19577 254175 19887 262961
rect 19577 254147 19625 254175
rect 19653 254147 19687 254175
rect 19715 254147 19749 254175
rect 19777 254147 19811 254175
rect 19839 254147 19887 254175
rect 19577 254113 19887 254147
rect 19577 254085 19625 254113
rect 19653 254085 19687 254113
rect 19715 254085 19749 254113
rect 19777 254085 19811 254113
rect 19839 254085 19887 254113
rect 19577 254051 19887 254085
rect 19577 254023 19625 254051
rect 19653 254023 19687 254051
rect 19715 254023 19749 254051
rect 19777 254023 19811 254051
rect 19839 254023 19887 254051
rect 19577 253989 19887 254023
rect 19577 253961 19625 253989
rect 19653 253961 19687 253989
rect 19715 253961 19749 253989
rect 19777 253961 19811 253989
rect 19839 253961 19887 253989
rect 19577 245175 19887 253961
rect 19577 245147 19625 245175
rect 19653 245147 19687 245175
rect 19715 245147 19749 245175
rect 19777 245147 19811 245175
rect 19839 245147 19887 245175
rect 19577 245113 19887 245147
rect 19577 245085 19625 245113
rect 19653 245085 19687 245113
rect 19715 245085 19749 245113
rect 19777 245085 19811 245113
rect 19839 245085 19887 245113
rect 19577 245051 19887 245085
rect 19577 245023 19625 245051
rect 19653 245023 19687 245051
rect 19715 245023 19749 245051
rect 19777 245023 19811 245051
rect 19839 245023 19887 245051
rect 19577 244989 19887 245023
rect 19577 244961 19625 244989
rect 19653 244961 19687 244989
rect 19715 244961 19749 244989
rect 19777 244961 19811 244989
rect 19839 244961 19887 244989
rect 19577 236175 19887 244961
rect 19577 236147 19625 236175
rect 19653 236147 19687 236175
rect 19715 236147 19749 236175
rect 19777 236147 19811 236175
rect 19839 236147 19887 236175
rect 19577 236113 19887 236147
rect 19577 236085 19625 236113
rect 19653 236085 19687 236113
rect 19715 236085 19749 236113
rect 19777 236085 19811 236113
rect 19839 236085 19887 236113
rect 19577 236051 19887 236085
rect 19577 236023 19625 236051
rect 19653 236023 19687 236051
rect 19715 236023 19749 236051
rect 19777 236023 19811 236051
rect 19839 236023 19887 236051
rect 19577 235989 19887 236023
rect 19577 235961 19625 235989
rect 19653 235961 19687 235989
rect 19715 235961 19749 235989
rect 19777 235961 19811 235989
rect 19839 235961 19887 235989
rect 19577 227175 19887 235961
rect 19577 227147 19625 227175
rect 19653 227147 19687 227175
rect 19715 227147 19749 227175
rect 19777 227147 19811 227175
rect 19839 227147 19887 227175
rect 19577 227113 19887 227147
rect 19577 227085 19625 227113
rect 19653 227085 19687 227113
rect 19715 227085 19749 227113
rect 19777 227085 19811 227113
rect 19839 227085 19887 227113
rect 19577 227051 19887 227085
rect 19577 227023 19625 227051
rect 19653 227023 19687 227051
rect 19715 227023 19749 227051
rect 19777 227023 19811 227051
rect 19839 227023 19887 227051
rect 19577 226989 19887 227023
rect 19577 226961 19625 226989
rect 19653 226961 19687 226989
rect 19715 226961 19749 226989
rect 19777 226961 19811 226989
rect 19839 226961 19887 226989
rect 19577 218175 19887 226961
rect 19577 218147 19625 218175
rect 19653 218147 19687 218175
rect 19715 218147 19749 218175
rect 19777 218147 19811 218175
rect 19839 218147 19887 218175
rect 19577 218113 19887 218147
rect 19577 218085 19625 218113
rect 19653 218085 19687 218113
rect 19715 218085 19749 218113
rect 19777 218085 19811 218113
rect 19839 218085 19887 218113
rect 19577 218051 19887 218085
rect 19577 218023 19625 218051
rect 19653 218023 19687 218051
rect 19715 218023 19749 218051
rect 19777 218023 19811 218051
rect 19839 218023 19887 218051
rect 19577 217989 19887 218023
rect 19577 217961 19625 217989
rect 19653 217961 19687 217989
rect 19715 217961 19749 217989
rect 19777 217961 19811 217989
rect 19839 217961 19887 217989
rect 19577 209175 19887 217961
rect 19577 209147 19625 209175
rect 19653 209147 19687 209175
rect 19715 209147 19749 209175
rect 19777 209147 19811 209175
rect 19839 209147 19887 209175
rect 19577 209113 19887 209147
rect 19577 209085 19625 209113
rect 19653 209085 19687 209113
rect 19715 209085 19749 209113
rect 19777 209085 19811 209113
rect 19839 209085 19887 209113
rect 19577 209051 19887 209085
rect 19577 209023 19625 209051
rect 19653 209023 19687 209051
rect 19715 209023 19749 209051
rect 19777 209023 19811 209051
rect 19839 209023 19887 209051
rect 19577 208989 19887 209023
rect 19577 208961 19625 208989
rect 19653 208961 19687 208989
rect 19715 208961 19749 208989
rect 19777 208961 19811 208989
rect 19839 208961 19887 208989
rect 19577 200175 19887 208961
rect 19577 200147 19625 200175
rect 19653 200147 19687 200175
rect 19715 200147 19749 200175
rect 19777 200147 19811 200175
rect 19839 200147 19887 200175
rect 19577 200113 19887 200147
rect 19577 200085 19625 200113
rect 19653 200085 19687 200113
rect 19715 200085 19749 200113
rect 19777 200085 19811 200113
rect 19839 200085 19887 200113
rect 19577 200051 19887 200085
rect 19577 200023 19625 200051
rect 19653 200023 19687 200051
rect 19715 200023 19749 200051
rect 19777 200023 19811 200051
rect 19839 200023 19887 200051
rect 19577 199989 19887 200023
rect 19577 199961 19625 199989
rect 19653 199961 19687 199989
rect 19715 199961 19749 199989
rect 19777 199961 19811 199989
rect 19839 199961 19887 199989
rect 19577 191175 19887 199961
rect 19577 191147 19625 191175
rect 19653 191147 19687 191175
rect 19715 191147 19749 191175
rect 19777 191147 19811 191175
rect 19839 191147 19887 191175
rect 19577 191113 19887 191147
rect 19577 191085 19625 191113
rect 19653 191085 19687 191113
rect 19715 191085 19749 191113
rect 19777 191085 19811 191113
rect 19839 191085 19887 191113
rect 19577 191051 19887 191085
rect 19577 191023 19625 191051
rect 19653 191023 19687 191051
rect 19715 191023 19749 191051
rect 19777 191023 19811 191051
rect 19839 191023 19887 191051
rect 19577 190989 19887 191023
rect 19577 190961 19625 190989
rect 19653 190961 19687 190989
rect 19715 190961 19749 190989
rect 19777 190961 19811 190989
rect 19839 190961 19887 190989
rect 19577 182175 19887 190961
rect 19577 182147 19625 182175
rect 19653 182147 19687 182175
rect 19715 182147 19749 182175
rect 19777 182147 19811 182175
rect 19839 182147 19887 182175
rect 19577 182113 19887 182147
rect 19577 182085 19625 182113
rect 19653 182085 19687 182113
rect 19715 182085 19749 182113
rect 19777 182085 19811 182113
rect 19839 182085 19887 182113
rect 19577 182051 19887 182085
rect 19577 182023 19625 182051
rect 19653 182023 19687 182051
rect 19715 182023 19749 182051
rect 19777 182023 19811 182051
rect 19839 182023 19887 182051
rect 19577 181989 19887 182023
rect 19577 181961 19625 181989
rect 19653 181961 19687 181989
rect 19715 181961 19749 181989
rect 19777 181961 19811 181989
rect 19839 181961 19887 181989
rect 19577 173175 19887 181961
rect 19577 173147 19625 173175
rect 19653 173147 19687 173175
rect 19715 173147 19749 173175
rect 19777 173147 19811 173175
rect 19839 173147 19887 173175
rect 19577 173113 19887 173147
rect 19577 173085 19625 173113
rect 19653 173085 19687 173113
rect 19715 173085 19749 173113
rect 19777 173085 19811 173113
rect 19839 173085 19887 173113
rect 19577 173051 19887 173085
rect 19577 173023 19625 173051
rect 19653 173023 19687 173051
rect 19715 173023 19749 173051
rect 19777 173023 19811 173051
rect 19839 173023 19887 173051
rect 19577 172989 19887 173023
rect 19577 172961 19625 172989
rect 19653 172961 19687 172989
rect 19715 172961 19749 172989
rect 19777 172961 19811 172989
rect 19839 172961 19887 172989
rect 19577 164175 19887 172961
rect 19577 164147 19625 164175
rect 19653 164147 19687 164175
rect 19715 164147 19749 164175
rect 19777 164147 19811 164175
rect 19839 164147 19887 164175
rect 19577 164113 19887 164147
rect 19577 164085 19625 164113
rect 19653 164085 19687 164113
rect 19715 164085 19749 164113
rect 19777 164085 19811 164113
rect 19839 164085 19887 164113
rect 19577 164051 19887 164085
rect 19577 164023 19625 164051
rect 19653 164023 19687 164051
rect 19715 164023 19749 164051
rect 19777 164023 19811 164051
rect 19839 164023 19887 164051
rect 19577 163989 19887 164023
rect 19577 163961 19625 163989
rect 19653 163961 19687 163989
rect 19715 163961 19749 163989
rect 19777 163961 19811 163989
rect 19839 163961 19887 163989
rect 19577 155175 19887 163961
rect 19577 155147 19625 155175
rect 19653 155147 19687 155175
rect 19715 155147 19749 155175
rect 19777 155147 19811 155175
rect 19839 155147 19887 155175
rect 19577 155113 19887 155147
rect 19577 155085 19625 155113
rect 19653 155085 19687 155113
rect 19715 155085 19749 155113
rect 19777 155085 19811 155113
rect 19839 155085 19887 155113
rect 19577 155051 19887 155085
rect 19577 155023 19625 155051
rect 19653 155023 19687 155051
rect 19715 155023 19749 155051
rect 19777 155023 19811 155051
rect 19839 155023 19887 155051
rect 19577 154989 19887 155023
rect 19577 154961 19625 154989
rect 19653 154961 19687 154989
rect 19715 154961 19749 154989
rect 19777 154961 19811 154989
rect 19839 154961 19887 154989
rect 19577 146175 19887 154961
rect 19577 146147 19625 146175
rect 19653 146147 19687 146175
rect 19715 146147 19749 146175
rect 19777 146147 19811 146175
rect 19839 146147 19887 146175
rect 19577 146113 19887 146147
rect 19577 146085 19625 146113
rect 19653 146085 19687 146113
rect 19715 146085 19749 146113
rect 19777 146085 19811 146113
rect 19839 146085 19887 146113
rect 19577 146051 19887 146085
rect 19577 146023 19625 146051
rect 19653 146023 19687 146051
rect 19715 146023 19749 146051
rect 19777 146023 19811 146051
rect 19839 146023 19887 146051
rect 19577 145989 19887 146023
rect 19577 145961 19625 145989
rect 19653 145961 19687 145989
rect 19715 145961 19749 145989
rect 19777 145961 19811 145989
rect 19839 145961 19887 145989
rect 19577 137175 19887 145961
rect 19577 137147 19625 137175
rect 19653 137147 19687 137175
rect 19715 137147 19749 137175
rect 19777 137147 19811 137175
rect 19839 137147 19887 137175
rect 19577 137113 19887 137147
rect 19577 137085 19625 137113
rect 19653 137085 19687 137113
rect 19715 137085 19749 137113
rect 19777 137085 19811 137113
rect 19839 137085 19887 137113
rect 19577 137051 19887 137085
rect 19577 137023 19625 137051
rect 19653 137023 19687 137051
rect 19715 137023 19749 137051
rect 19777 137023 19811 137051
rect 19839 137023 19887 137051
rect 19577 136989 19887 137023
rect 19577 136961 19625 136989
rect 19653 136961 19687 136989
rect 19715 136961 19749 136989
rect 19777 136961 19811 136989
rect 19839 136961 19887 136989
rect 19577 128175 19887 136961
rect 19577 128147 19625 128175
rect 19653 128147 19687 128175
rect 19715 128147 19749 128175
rect 19777 128147 19811 128175
rect 19839 128147 19887 128175
rect 19577 128113 19887 128147
rect 19577 128085 19625 128113
rect 19653 128085 19687 128113
rect 19715 128085 19749 128113
rect 19777 128085 19811 128113
rect 19839 128085 19887 128113
rect 19577 128051 19887 128085
rect 19577 128023 19625 128051
rect 19653 128023 19687 128051
rect 19715 128023 19749 128051
rect 19777 128023 19811 128051
rect 19839 128023 19887 128051
rect 19577 127989 19887 128023
rect 19577 127961 19625 127989
rect 19653 127961 19687 127989
rect 19715 127961 19749 127989
rect 19777 127961 19811 127989
rect 19839 127961 19887 127989
rect 19577 119175 19887 127961
rect 19577 119147 19625 119175
rect 19653 119147 19687 119175
rect 19715 119147 19749 119175
rect 19777 119147 19811 119175
rect 19839 119147 19887 119175
rect 19577 119113 19887 119147
rect 19577 119085 19625 119113
rect 19653 119085 19687 119113
rect 19715 119085 19749 119113
rect 19777 119085 19811 119113
rect 19839 119085 19887 119113
rect 19577 119051 19887 119085
rect 19577 119023 19625 119051
rect 19653 119023 19687 119051
rect 19715 119023 19749 119051
rect 19777 119023 19811 119051
rect 19839 119023 19887 119051
rect 19577 118989 19887 119023
rect 19577 118961 19625 118989
rect 19653 118961 19687 118989
rect 19715 118961 19749 118989
rect 19777 118961 19811 118989
rect 19839 118961 19887 118989
rect 19577 110175 19887 118961
rect 19577 110147 19625 110175
rect 19653 110147 19687 110175
rect 19715 110147 19749 110175
rect 19777 110147 19811 110175
rect 19839 110147 19887 110175
rect 19577 110113 19887 110147
rect 19577 110085 19625 110113
rect 19653 110085 19687 110113
rect 19715 110085 19749 110113
rect 19777 110085 19811 110113
rect 19839 110085 19887 110113
rect 19577 110051 19887 110085
rect 19577 110023 19625 110051
rect 19653 110023 19687 110051
rect 19715 110023 19749 110051
rect 19777 110023 19811 110051
rect 19839 110023 19887 110051
rect 19577 109989 19887 110023
rect 19577 109961 19625 109989
rect 19653 109961 19687 109989
rect 19715 109961 19749 109989
rect 19777 109961 19811 109989
rect 19839 109961 19887 109989
rect 19577 101175 19887 109961
rect 19577 101147 19625 101175
rect 19653 101147 19687 101175
rect 19715 101147 19749 101175
rect 19777 101147 19811 101175
rect 19839 101147 19887 101175
rect 19577 101113 19887 101147
rect 19577 101085 19625 101113
rect 19653 101085 19687 101113
rect 19715 101085 19749 101113
rect 19777 101085 19811 101113
rect 19839 101085 19887 101113
rect 19577 101051 19887 101085
rect 19577 101023 19625 101051
rect 19653 101023 19687 101051
rect 19715 101023 19749 101051
rect 19777 101023 19811 101051
rect 19839 101023 19887 101051
rect 19577 100989 19887 101023
rect 19577 100961 19625 100989
rect 19653 100961 19687 100989
rect 19715 100961 19749 100989
rect 19777 100961 19811 100989
rect 19839 100961 19887 100989
rect 19577 92175 19887 100961
rect 19577 92147 19625 92175
rect 19653 92147 19687 92175
rect 19715 92147 19749 92175
rect 19777 92147 19811 92175
rect 19839 92147 19887 92175
rect 19577 92113 19887 92147
rect 19577 92085 19625 92113
rect 19653 92085 19687 92113
rect 19715 92085 19749 92113
rect 19777 92085 19811 92113
rect 19839 92085 19887 92113
rect 19577 92051 19887 92085
rect 19577 92023 19625 92051
rect 19653 92023 19687 92051
rect 19715 92023 19749 92051
rect 19777 92023 19811 92051
rect 19839 92023 19887 92051
rect 19577 91989 19887 92023
rect 19577 91961 19625 91989
rect 19653 91961 19687 91989
rect 19715 91961 19749 91989
rect 19777 91961 19811 91989
rect 19839 91961 19887 91989
rect 19577 83175 19887 91961
rect 19577 83147 19625 83175
rect 19653 83147 19687 83175
rect 19715 83147 19749 83175
rect 19777 83147 19811 83175
rect 19839 83147 19887 83175
rect 19577 83113 19887 83147
rect 19577 83085 19625 83113
rect 19653 83085 19687 83113
rect 19715 83085 19749 83113
rect 19777 83085 19811 83113
rect 19839 83085 19887 83113
rect 19577 83051 19887 83085
rect 19577 83023 19625 83051
rect 19653 83023 19687 83051
rect 19715 83023 19749 83051
rect 19777 83023 19811 83051
rect 19839 83023 19887 83051
rect 19577 82989 19887 83023
rect 19577 82961 19625 82989
rect 19653 82961 19687 82989
rect 19715 82961 19749 82989
rect 19777 82961 19811 82989
rect 19839 82961 19887 82989
rect 19577 74175 19887 82961
rect 19577 74147 19625 74175
rect 19653 74147 19687 74175
rect 19715 74147 19749 74175
rect 19777 74147 19811 74175
rect 19839 74147 19887 74175
rect 19577 74113 19887 74147
rect 19577 74085 19625 74113
rect 19653 74085 19687 74113
rect 19715 74085 19749 74113
rect 19777 74085 19811 74113
rect 19839 74085 19887 74113
rect 19577 74051 19887 74085
rect 19577 74023 19625 74051
rect 19653 74023 19687 74051
rect 19715 74023 19749 74051
rect 19777 74023 19811 74051
rect 19839 74023 19887 74051
rect 19577 73989 19887 74023
rect 19577 73961 19625 73989
rect 19653 73961 19687 73989
rect 19715 73961 19749 73989
rect 19777 73961 19811 73989
rect 19839 73961 19887 73989
rect 19577 65175 19887 73961
rect 19577 65147 19625 65175
rect 19653 65147 19687 65175
rect 19715 65147 19749 65175
rect 19777 65147 19811 65175
rect 19839 65147 19887 65175
rect 19577 65113 19887 65147
rect 19577 65085 19625 65113
rect 19653 65085 19687 65113
rect 19715 65085 19749 65113
rect 19777 65085 19811 65113
rect 19839 65085 19887 65113
rect 19577 65051 19887 65085
rect 19577 65023 19625 65051
rect 19653 65023 19687 65051
rect 19715 65023 19749 65051
rect 19777 65023 19811 65051
rect 19839 65023 19887 65051
rect 19577 64989 19887 65023
rect 19577 64961 19625 64989
rect 19653 64961 19687 64989
rect 19715 64961 19749 64989
rect 19777 64961 19811 64989
rect 19839 64961 19887 64989
rect 19577 56175 19887 64961
rect 19577 56147 19625 56175
rect 19653 56147 19687 56175
rect 19715 56147 19749 56175
rect 19777 56147 19811 56175
rect 19839 56147 19887 56175
rect 19577 56113 19887 56147
rect 19577 56085 19625 56113
rect 19653 56085 19687 56113
rect 19715 56085 19749 56113
rect 19777 56085 19811 56113
rect 19839 56085 19887 56113
rect 19577 56051 19887 56085
rect 19577 56023 19625 56051
rect 19653 56023 19687 56051
rect 19715 56023 19749 56051
rect 19777 56023 19811 56051
rect 19839 56023 19887 56051
rect 19577 55989 19887 56023
rect 19577 55961 19625 55989
rect 19653 55961 19687 55989
rect 19715 55961 19749 55989
rect 19777 55961 19811 55989
rect 19839 55961 19887 55989
rect 19577 47175 19887 55961
rect 19577 47147 19625 47175
rect 19653 47147 19687 47175
rect 19715 47147 19749 47175
rect 19777 47147 19811 47175
rect 19839 47147 19887 47175
rect 19577 47113 19887 47147
rect 19577 47085 19625 47113
rect 19653 47085 19687 47113
rect 19715 47085 19749 47113
rect 19777 47085 19811 47113
rect 19839 47085 19887 47113
rect 19577 47051 19887 47085
rect 19577 47023 19625 47051
rect 19653 47023 19687 47051
rect 19715 47023 19749 47051
rect 19777 47023 19811 47051
rect 19839 47023 19887 47051
rect 19577 46989 19887 47023
rect 19577 46961 19625 46989
rect 19653 46961 19687 46989
rect 19715 46961 19749 46989
rect 19777 46961 19811 46989
rect 19839 46961 19887 46989
rect 19577 38175 19887 46961
rect 19577 38147 19625 38175
rect 19653 38147 19687 38175
rect 19715 38147 19749 38175
rect 19777 38147 19811 38175
rect 19839 38147 19887 38175
rect 19577 38113 19887 38147
rect 19577 38085 19625 38113
rect 19653 38085 19687 38113
rect 19715 38085 19749 38113
rect 19777 38085 19811 38113
rect 19839 38085 19887 38113
rect 19577 38051 19887 38085
rect 19577 38023 19625 38051
rect 19653 38023 19687 38051
rect 19715 38023 19749 38051
rect 19777 38023 19811 38051
rect 19839 38023 19887 38051
rect 19577 37989 19887 38023
rect 19577 37961 19625 37989
rect 19653 37961 19687 37989
rect 19715 37961 19749 37989
rect 19777 37961 19811 37989
rect 19839 37961 19887 37989
rect 19577 29175 19887 37961
rect 19577 29147 19625 29175
rect 19653 29147 19687 29175
rect 19715 29147 19749 29175
rect 19777 29147 19811 29175
rect 19839 29147 19887 29175
rect 19577 29113 19887 29147
rect 19577 29085 19625 29113
rect 19653 29085 19687 29113
rect 19715 29085 19749 29113
rect 19777 29085 19811 29113
rect 19839 29085 19887 29113
rect 19577 29051 19887 29085
rect 19577 29023 19625 29051
rect 19653 29023 19687 29051
rect 19715 29023 19749 29051
rect 19777 29023 19811 29051
rect 19839 29023 19887 29051
rect 19577 28989 19887 29023
rect 19577 28961 19625 28989
rect 19653 28961 19687 28989
rect 19715 28961 19749 28989
rect 19777 28961 19811 28989
rect 19839 28961 19887 28989
rect 19577 20175 19887 28961
rect 19577 20147 19625 20175
rect 19653 20147 19687 20175
rect 19715 20147 19749 20175
rect 19777 20147 19811 20175
rect 19839 20147 19887 20175
rect 19577 20113 19887 20147
rect 19577 20085 19625 20113
rect 19653 20085 19687 20113
rect 19715 20085 19749 20113
rect 19777 20085 19811 20113
rect 19839 20085 19887 20113
rect 19577 20051 19887 20085
rect 19577 20023 19625 20051
rect 19653 20023 19687 20051
rect 19715 20023 19749 20051
rect 19777 20023 19811 20051
rect 19839 20023 19887 20051
rect 19577 19989 19887 20023
rect 19577 19961 19625 19989
rect 19653 19961 19687 19989
rect 19715 19961 19749 19989
rect 19777 19961 19811 19989
rect 19839 19961 19887 19989
rect 19577 11175 19887 19961
rect 19577 11147 19625 11175
rect 19653 11147 19687 11175
rect 19715 11147 19749 11175
rect 19777 11147 19811 11175
rect 19839 11147 19887 11175
rect 19577 11113 19887 11147
rect 19577 11085 19625 11113
rect 19653 11085 19687 11113
rect 19715 11085 19749 11113
rect 19777 11085 19811 11113
rect 19839 11085 19887 11113
rect 19577 11051 19887 11085
rect 19577 11023 19625 11051
rect 19653 11023 19687 11051
rect 19715 11023 19749 11051
rect 19777 11023 19811 11051
rect 19839 11023 19887 11051
rect 19577 10989 19887 11023
rect 19577 10961 19625 10989
rect 19653 10961 19687 10989
rect 19715 10961 19749 10989
rect 19777 10961 19811 10989
rect 19839 10961 19887 10989
rect 19577 2175 19887 10961
rect 19577 2147 19625 2175
rect 19653 2147 19687 2175
rect 19715 2147 19749 2175
rect 19777 2147 19811 2175
rect 19839 2147 19887 2175
rect 19577 2113 19887 2147
rect 19577 2085 19625 2113
rect 19653 2085 19687 2113
rect 19715 2085 19749 2113
rect 19777 2085 19811 2113
rect 19839 2085 19887 2113
rect 19577 2051 19887 2085
rect 19577 2023 19625 2051
rect 19653 2023 19687 2051
rect 19715 2023 19749 2051
rect 19777 2023 19811 2051
rect 19839 2023 19887 2051
rect 19577 1989 19887 2023
rect 19577 1961 19625 1989
rect 19653 1961 19687 1989
rect 19715 1961 19749 1989
rect 19777 1961 19811 1989
rect 19839 1961 19887 1989
rect 19577 -80 19887 1961
rect 19577 -108 19625 -80
rect 19653 -108 19687 -80
rect 19715 -108 19749 -80
rect 19777 -108 19811 -80
rect 19839 -108 19887 -80
rect 19577 -142 19887 -108
rect 19577 -170 19625 -142
rect 19653 -170 19687 -142
rect 19715 -170 19749 -142
rect 19777 -170 19811 -142
rect 19839 -170 19887 -142
rect 19577 -204 19887 -170
rect 19577 -232 19625 -204
rect 19653 -232 19687 -204
rect 19715 -232 19749 -204
rect 19777 -232 19811 -204
rect 19839 -232 19887 -204
rect 19577 -266 19887 -232
rect 19577 -294 19625 -266
rect 19653 -294 19687 -266
rect 19715 -294 19749 -266
rect 19777 -294 19811 -266
rect 19839 -294 19887 -266
rect 19577 -822 19887 -294
rect 21437 299086 21747 299134
rect 21437 299058 21485 299086
rect 21513 299058 21547 299086
rect 21575 299058 21609 299086
rect 21637 299058 21671 299086
rect 21699 299058 21747 299086
rect 21437 299024 21747 299058
rect 21437 298996 21485 299024
rect 21513 298996 21547 299024
rect 21575 298996 21609 299024
rect 21637 298996 21671 299024
rect 21699 298996 21747 299024
rect 21437 298962 21747 298996
rect 21437 298934 21485 298962
rect 21513 298934 21547 298962
rect 21575 298934 21609 298962
rect 21637 298934 21671 298962
rect 21699 298934 21747 298962
rect 21437 298900 21747 298934
rect 21437 298872 21485 298900
rect 21513 298872 21547 298900
rect 21575 298872 21609 298900
rect 21637 298872 21671 298900
rect 21699 298872 21747 298900
rect 21437 293175 21747 298872
rect 21437 293147 21485 293175
rect 21513 293147 21547 293175
rect 21575 293147 21609 293175
rect 21637 293147 21671 293175
rect 21699 293147 21747 293175
rect 21437 293113 21747 293147
rect 21437 293085 21485 293113
rect 21513 293085 21547 293113
rect 21575 293085 21609 293113
rect 21637 293085 21671 293113
rect 21699 293085 21747 293113
rect 21437 293051 21747 293085
rect 21437 293023 21485 293051
rect 21513 293023 21547 293051
rect 21575 293023 21609 293051
rect 21637 293023 21671 293051
rect 21699 293023 21747 293051
rect 21437 292989 21747 293023
rect 21437 292961 21485 292989
rect 21513 292961 21547 292989
rect 21575 292961 21609 292989
rect 21637 292961 21671 292989
rect 21699 292961 21747 292989
rect 21437 284175 21747 292961
rect 21437 284147 21485 284175
rect 21513 284147 21547 284175
rect 21575 284147 21609 284175
rect 21637 284147 21671 284175
rect 21699 284147 21747 284175
rect 21437 284113 21747 284147
rect 21437 284085 21485 284113
rect 21513 284085 21547 284113
rect 21575 284085 21609 284113
rect 21637 284085 21671 284113
rect 21699 284085 21747 284113
rect 21437 284051 21747 284085
rect 21437 284023 21485 284051
rect 21513 284023 21547 284051
rect 21575 284023 21609 284051
rect 21637 284023 21671 284051
rect 21699 284023 21747 284051
rect 21437 283989 21747 284023
rect 21437 283961 21485 283989
rect 21513 283961 21547 283989
rect 21575 283961 21609 283989
rect 21637 283961 21671 283989
rect 21699 283961 21747 283989
rect 21437 275175 21747 283961
rect 21437 275147 21485 275175
rect 21513 275147 21547 275175
rect 21575 275147 21609 275175
rect 21637 275147 21671 275175
rect 21699 275147 21747 275175
rect 21437 275113 21747 275147
rect 21437 275085 21485 275113
rect 21513 275085 21547 275113
rect 21575 275085 21609 275113
rect 21637 275085 21671 275113
rect 21699 275085 21747 275113
rect 21437 275051 21747 275085
rect 21437 275023 21485 275051
rect 21513 275023 21547 275051
rect 21575 275023 21609 275051
rect 21637 275023 21671 275051
rect 21699 275023 21747 275051
rect 21437 274989 21747 275023
rect 21437 274961 21485 274989
rect 21513 274961 21547 274989
rect 21575 274961 21609 274989
rect 21637 274961 21671 274989
rect 21699 274961 21747 274989
rect 21437 266175 21747 274961
rect 21437 266147 21485 266175
rect 21513 266147 21547 266175
rect 21575 266147 21609 266175
rect 21637 266147 21671 266175
rect 21699 266147 21747 266175
rect 21437 266113 21747 266147
rect 21437 266085 21485 266113
rect 21513 266085 21547 266113
rect 21575 266085 21609 266113
rect 21637 266085 21671 266113
rect 21699 266085 21747 266113
rect 21437 266051 21747 266085
rect 21437 266023 21485 266051
rect 21513 266023 21547 266051
rect 21575 266023 21609 266051
rect 21637 266023 21671 266051
rect 21699 266023 21747 266051
rect 21437 265989 21747 266023
rect 21437 265961 21485 265989
rect 21513 265961 21547 265989
rect 21575 265961 21609 265989
rect 21637 265961 21671 265989
rect 21699 265961 21747 265989
rect 21437 257175 21747 265961
rect 21437 257147 21485 257175
rect 21513 257147 21547 257175
rect 21575 257147 21609 257175
rect 21637 257147 21671 257175
rect 21699 257147 21747 257175
rect 21437 257113 21747 257147
rect 21437 257085 21485 257113
rect 21513 257085 21547 257113
rect 21575 257085 21609 257113
rect 21637 257085 21671 257113
rect 21699 257085 21747 257113
rect 21437 257051 21747 257085
rect 21437 257023 21485 257051
rect 21513 257023 21547 257051
rect 21575 257023 21609 257051
rect 21637 257023 21671 257051
rect 21699 257023 21747 257051
rect 21437 256989 21747 257023
rect 21437 256961 21485 256989
rect 21513 256961 21547 256989
rect 21575 256961 21609 256989
rect 21637 256961 21671 256989
rect 21699 256961 21747 256989
rect 21437 248175 21747 256961
rect 21437 248147 21485 248175
rect 21513 248147 21547 248175
rect 21575 248147 21609 248175
rect 21637 248147 21671 248175
rect 21699 248147 21747 248175
rect 21437 248113 21747 248147
rect 21437 248085 21485 248113
rect 21513 248085 21547 248113
rect 21575 248085 21609 248113
rect 21637 248085 21671 248113
rect 21699 248085 21747 248113
rect 21437 248051 21747 248085
rect 21437 248023 21485 248051
rect 21513 248023 21547 248051
rect 21575 248023 21609 248051
rect 21637 248023 21671 248051
rect 21699 248023 21747 248051
rect 21437 247989 21747 248023
rect 21437 247961 21485 247989
rect 21513 247961 21547 247989
rect 21575 247961 21609 247989
rect 21637 247961 21671 247989
rect 21699 247961 21747 247989
rect 21437 239175 21747 247961
rect 21437 239147 21485 239175
rect 21513 239147 21547 239175
rect 21575 239147 21609 239175
rect 21637 239147 21671 239175
rect 21699 239147 21747 239175
rect 21437 239113 21747 239147
rect 21437 239085 21485 239113
rect 21513 239085 21547 239113
rect 21575 239085 21609 239113
rect 21637 239085 21671 239113
rect 21699 239085 21747 239113
rect 21437 239051 21747 239085
rect 21437 239023 21485 239051
rect 21513 239023 21547 239051
rect 21575 239023 21609 239051
rect 21637 239023 21671 239051
rect 21699 239023 21747 239051
rect 21437 238989 21747 239023
rect 21437 238961 21485 238989
rect 21513 238961 21547 238989
rect 21575 238961 21609 238989
rect 21637 238961 21671 238989
rect 21699 238961 21747 238989
rect 21437 230175 21747 238961
rect 21437 230147 21485 230175
rect 21513 230147 21547 230175
rect 21575 230147 21609 230175
rect 21637 230147 21671 230175
rect 21699 230147 21747 230175
rect 21437 230113 21747 230147
rect 21437 230085 21485 230113
rect 21513 230085 21547 230113
rect 21575 230085 21609 230113
rect 21637 230085 21671 230113
rect 21699 230085 21747 230113
rect 21437 230051 21747 230085
rect 21437 230023 21485 230051
rect 21513 230023 21547 230051
rect 21575 230023 21609 230051
rect 21637 230023 21671 230051
rect 21699 230023 21747 230051
rect 21437 229989 21747 230023
rect 21437 229961 21485 229989
rect 21513 229961 21547 229989
rect 21575 229961 21609 229989
rect 21637 229961 21671 229989
rect 21699 229961 21747 229989
rect 21437 221175 21747 229961
rect 21437 221147 21485 221175
rect 21513 221147 21547 221175
rect 21575 221147 21609 221175
rect 21637 221147 21671 221175
rect 21699 221147 21747 221175
rect 21437 221113 21747 221147
rect 21437 221085 21485 221113
rect 21513 221085 21547 221113
rect 21575 221085 21609 221113
rect 21637 221085 21671 221113
rect 21699 221085 21747 221113
rect 21437 221051 21747 221085
rect 21437 221023 21485 221051
rect 21513 221023 21547 221051
rect 21575 221023 21609 221051
rect 21637 221023 21671 221051
rect 21699 221023 21747 221051
rect 21437 220989 21747 221023
rect 21437 220961 21485 220989
rect 21513 220961 21547 220989
rect 21575 220961 21609 220989
rect 21637 220961 21671 220989
rect 21699 220961 21747 220989
rect 21437 212175 21747 220961
rect 21437 212147 21485 212175
rect 21513 212147 21547 212175
rect 21575 212147 21609 212175
rect 21637 212147 21671 212175
rect 21699 212147 21747 212175
rect 21437 212113 21747 212147
rect 21437 212085 21485 212113
rect 21513 212085 21547 212113
rect 21575 212085 21609 212113
rect 21637 212085 21671 212113
rect 21699 212085 21747 212113
rect 21437 212051 21747 212085
rect 21437 212023 21485 212051
rect 21513 212023 21547 212051
rect 21575 212023 21609 212051
rect 21637 212023 21671 212051
rect 21699 212023 21747 212051
rect 21437 211989 21747 212023
rect 21437 211961 21485 211989
rect 21513 211961 21547 211989
rect 21575 211961 21609 211989
rect 21637 211961 21671 211989
rect 21699 211961 21747 211989
rect 21437 203175 21747 211961
rect 21437 203147 21485 203175
rect 21513 203147 21547 203175
rect 21575 203147 21609 203175
rect 21637 203147 21671 203175
rect 21699 203147 21747 203175
rect 21437 203113 21747 203147
rect 21437 203085 21485 203113
rect 21513 203085 21547 203113
rect 21575 203085 21609 203113
rect 21637 203085 21671 203113
rect 21699 203085 21747 203113
rect 21437 203051 21747 203085
rect 21437 203023 21485 203051
rect 21513 203023 21547 203051
rect 21575 203023 21609 203051
rect 21637 203023 21671 203051
rect 21699 203023 21747 203051
rect 21437 202989 21747 203023
rect 21437 202961 21485 202989
rect 21513 202961 21547 202989
rect 21575 202961 21609 202989
rect 21637 202961 21671 202989
rect 21699 202961 21747 202989
rect 21437 194175 21747 202961
rect 21437 194147 21485 194175
rect 21513 194147 21547 194175
rect 21575 194147 21609 194175
rect 21637 194147 21671 194175
rect 21699 194147 21747 194175
rect 21437 194113 21747 194147
rect 21437 194085 21485 194113
rect 21513 194085 21547 194113
rect 21575 194085 21609 194113
rect 21637 194085 21671 194113
rect 21699 194085 21747 194113
rect 21437 194051 21747 194085
rect 21437 194023 21485 194051
rect 21513 194023 21547 194051
rect 21575 194023 21609 194051
rect 21637 194023 21671 194051
rect 21699 194023 21747 194051
rect 21437 193989 21747 194023
rect 21437 193961 21485 193989
rect 21513 193961 21547 193989
rect 21575 193961 21609 193989
rect 21637 193961 21671 193989
rect 21699 193961 21747 193989
rect 21437 185175 21747 193961
rect 21437 185147 21485 185175
rect 21513 185147 21547 185175
rect 21575 185147 21609 185175
rect 21637 185147 21671 185175
rect 21699 185147 21747 185175
rect 21437 185113 21747 185147
rect 21437 185085 21485 185113
rect 21513 185085 21547 185113
rect 21575 185085 21609 185113
rect 21637 185085 21671 185113
rect 21699 185085 21747 185113
rect 21437 185051 21747 185085
rect 21437 185023 21485 185051
rect 21513 185023 21547 185051
rect 21575 185023 21609 185051
rect 21637 185023 21671 185051
rect 21699 185023 21747 185051
rect 21437 184989 21747 185023
rect 21437 184961 21485 184989
rect 21513 184961 21547 184989
rect 21575 184961 21609 184989
rect 21637 184961 21671 184989
rect 21699 184961 21747 184989
rect 21437 176175 21747 184961
rect 21437 176147 21485 176175
rect 21513 176147 21547 176175
rect 21575 176147 21609 176175
rect 21637 176147 21671 176175
rect 21699 176147 21747 176175
rect 21437 176113 21747 176147
rect 21437 176085 21485 176113
rect 21513 176085 21547 176113
rect 21575 176085 21609 176113
rect 21637 176085 21671 176113
rect 21699 176085 21747 176113
rect 21437 176051 21747 176085
rect 21437 176023 21485 176051
rect 21513 176023 21547 176051
rect 21575 176023 21609 176051
rect 21637 176023 21671 176051
rect 21699 176023 21747 176051
rect 21437 175989 21747 176023
rect 21437 175961 21485 175989
rect 21513 175961 21547 175989
rect 21575 175961 21609 175989
rect 21637 175961 21671 175989
rect 21699 175961 21747 175989
rect 21437 167175 21747 175961
rect 21437 167147 21485 167175
rect 21513 167147 21547 167175
rect 21575 167147 21609 167175
rect 21637 167147 21671 167175
rect 21699 167147 21747 167175
rect 21437 167113 21747 167147
rect 21437 167085 21485 167113
rect 21513 167085 21547 167113
rect 21575 167085 21609 167113
rect 21637 167085 21671 167113
rect 21699 167085 21747 167113
rect 21437 167051 21747 167085
rect 21437 167023 21485 167051
rect 21513 167023 21547 167051
rect 21575 167023 21609 167051
rect 21637 167023 21671 167051
rect 21699 167023 21747 167051
rect 21437 166989 21747 167023
rect 21437 166961 21485 166989
rect 21513 166961 21547 166989
rect 21575 166961 21609 166989
rect 21637 166961 21671 166989
rect 21699 166961 21747 166989
rect 21437 158175 21747 166961
rect 21437 158147 21485 158175
rect 21513 158147 21547 158175
rect 21575 158147 21609 158175
rect 21637 158147 21671 158175
rect 21699 158147 21747 158175
rect 21437 158113 21747 158147
rect 21437 158085 21485 158113
rect 21513 158085 21547 158113
rect 21575 158085 21609 158113
rect 21637 158085 21671 158113
rect 21699 158085 21747 158113
rect 21437 158051 21747 158085
rect 21437 158023 21485 158051
rect 21513 158023 21547 158051
rect 21575 158023 21609 158051
rect 21637 158023 21671 158051
rect 21699 158023 21747 158051
rect 21437 157989 21747 158023
rect 21437 157961 21485 157989
rect 21513 157961 21547 157989
rect 21575 157961 21609 157989
rect 21637 157961 21671 157989
rect 21699 157961 21747 157989
rect 21437 149175 21747 157961
rect 21437 149147 21485 149175
rect 21513 149147 21547 149175
rect 21575 149147 21609 149175
rect 21637 149147 21671 149175
rect 21699 149147 21747 149175
rect 21437 149113 21747 149147
rect 21437 149085 21485 149113
rect 21513 149085 21547 149113
rect 21575 149085 21609 149113
rect 21637 149085 21671 149113
rect 21699 149085 21747 149113
rect 21437 149051 21747 149085
rect 21437 149023 21485 149051
rect 21513 149023 21547 149051
rect 21575 149023 21609 149051
rect 21637 149023 21671 149051
rect 21699 149023 21747 149051
rect 21437 148989 21747 149023
rect 21437 148961 21485 148989
rect 21513 148961 21547 148989
rect 21575 148961 21609 148989
rect 21637 148961 21671 148989
rect 21699 148961 21747 148989
rect 21437 140175 21747 148961
rect 21437 140147 21485 140175
rect 21513 140147 21547 140175
rect 21575 140147 21609 140175
rect 21637 140147 21671 140175
rect 21699 140147 21747 140175
rect 21437 140113 21747 140147
rect 21437 140085 21485 140113
rect 21513 140085 21547 140113
rect 21575 140085 21609 140113
rect 21637 140085 21671 140113
rect 21699 140085 21747 140113
rect 21437 140051 21747 140085
rect 21437 140023 21485 140051
rect 21513 140023 21547 140051
rect 21575 140023 21609 140051
rect 21637 140023 21671 140051
rect 21699 140023 21747 140051
rect 21437 139989 21747 140023
rect 21437 139961 21485 139989
rect 21513 139961 21547 139989
rect 21575 139961 21609 139989
rect 21637 139961 21671 139989
rect 21699 139961 21747 139989
rect 21437 131175 21747 139961
rect 21437 131147 21485 131175
rect 21513 131147 21547 131175
rect 21575 131147 21609 131175
rect 21637 131147 21671 131175
rect 21699 131147 21747 131175
rect 21437 131113 21747 131147
rect 21437 131085 21485 131113
rect 21513 131085 21547 131113
rect 21575 131085 21609 131113
rect 21637 131085 21671 131113
rect 21699 131085 21747 131113
rect 21437 131051 21747 131085
rect 21437 131023 21485 131051
rect 21513 131023 21547 131051
rect 21575 131023 21609 131051
rect 21637 131023 21671 131051
rect 21699 131023 21747 131051
rect 21437 130989 21747 131023
rect 21437 130961 21485 130989
rect 21513 130961 21547 130989
rect 21575 130961 21609 130989
rect 21637 130961 21671 130989
rect 21699 130961 21747 130989
rect 21437 122175 21747 130961
rect 21437 122147 21485 122175
rect 21513 122147 21547 122175
rect 21575 122147 21609 122175
rect 21637 122147 21671 122175
rect 21699 122147 21747 122175
rect 21437 122113 21747 122147
rect 21437 122085 21485 122113
rect 21513 122085 21547 122113
rect 21575 122085 21609 122113
rect 21637 122085 21671 122113
rect 21699 122085 21747 122113
rect 21437 122051 21747 122085
rect 21437 122023 21485 122051
rect 21513 122023 21547 122051
rect 21575 122023 21609 122051
rect 21637 122023 21671 122051
rect 21699 122023 21747 122051
rect 21437 121989 21747 122023
rect 21437 121961 21485 121989
rect 21513 121961 21547 121989
rect 21575 121961 21609 121989
rect 21637 121961 21671 121989
rect 21699 121961 21747 121989
rect 21437 113175 21747 121961
rect 21437 113147 21485 113175
rect 21513 113147 21547 113175
rect 21575 113147 21609 113175
rect 21637 113147 21671 113175
rect 21699 113147 21747 113175
rect 21437 113113 21747 113147
rect 21437 113085 21485 113113
rect 21513 113085 21547 113113
rect 21575 113085 21609 113113
rect 21637 113085 21671 113113
rect 21699 113085 21747 113113
rect 21437 113051 21747 113085
rect 21437 113023 21485 113051
rect 21513 113023 21547 113051
rect 21575 113023 21609 113051
rect 21637 113023 21671 113051
rect 21699 113023 21747 113051
rect 21437 112989 21747 113023
rect 21437 112961 21485 112989
rect 21513 112961 21547 112989
rect 21575 112961 21609 112989
rect 21637 112961 21671 112989
rect 21699 112961 21747 112989
rect 21437 104175 21747 112961
rect 21437 104147 21485 104175
rect 21513 104147 21547 104175
rect 21575 104147 21609 104175
rect 21637 104147 21671 104175
rect 21699 104147 21747 104175
rect 21437 104113 21747 104147
rect 21437 104085 21485 104113
rect 21513 104085 21547 104113
rect 21575 104085 21609 104113
rect 21637 104085 21671 104113
rect 21699 104085 21747 104113
rect 21437 104051 21747 104085
rect 21437 104023 21485 104051
rect 21513 104023 21547 104051
rect 21575 104023 21609 104051
rect 21637 104023 21671 104051
rect 21699 104023 21747 104051
rect 21437 103989 21747 104023
rect 21437 103961 21485 103989
rect 21513 103961 21547 103989
rect 21575 103961 21609 103989
rect 21637 103961 21671 103989
rect 21699 103961 21747 103989
rect 21437 95175 21747 103961
rect 21437 95147 21485 95175
rect 21513 95147 21547 95175
rect 21575 95147 21609 95175
rect 21637 95147 21671 95175
rect 21699 95147 21747 95175
rect 21437 95113 21747 95147
rect 21437 95085 21485 95113
rect 21513 95085 21547 95113
rect 21575 95085 21609 95113
rect 21637 95085 21671 95113
rect 21699 95085 21747 95113
rect 21437 95051 21747 95085
rect 21437 95023 21485 95051
rect 21513 95023 21547 95051
rect 21575 95023 21609 95051
rect 21637 95023 21671 95051
rect 21699 95023 21747 95051
rect 21437 94989 21747 95023
rect 21437 94961 21485 94989
rect 21513 94961 21547 94989
rect 21575 94961 21609 94989
rect 21637 94961 21671 94989
rect 21699 94961 21747 94989
rect 21437 86175 21747 94961
rect 21437 86147 21485 86175
rect 21513 86147 21547 86175
rect 21575 86147 21609 86175
rect 21637 86147 21671 86175
rect 21699 86147 21747 86175
rect 21437 86113 21747 86147
rect 21437 86085 21485 86113
rect 21513 86085 21547 86113
rect 21575 86085 21609 86113
rect 21637 86085 21671 86113
rect 21699 86085 21747 86113
rect 21437 86051 21747 86085
rect 21437 86023 21485 86051
rect 21513 86023 21547 86051
rect 21575 86023 21609 86051
rect 21637 86023 21671 86051
rect 21699 86023 21747 86051
rect 21437 85989 21747 86023
rect 21437 85961 21485 85989
rect 21513 85961 21547 85989
rect 21575 85961 21609 85989
rect 21637 85961 21671 85989
rect 21699 85961 21747 85989
rect 21437 77175 21747 85961
rect 21437 77147 21485 77175
rect 21513 77147 21547 77175
rect 21575 77147 21609 77175
rect 21637 77147 21671 77175
rect 21699 77147 21747 77175
rect 21437 77113 21747 77147
rect 21437 77085 21485 77113
rect 21513 77085 21547 77113
rect 21575 77085 21609 77113
rect 21637 77085 21671 77113
rect 21699 77085 21747 77113
rect 21437 77051 21747 77085
rect 21437 77023 21485 77051
rect 21513 77023 21547 77051
rect 21575 77023 21609 77051
rect 21637 77023 21671 77051
rect 21699 77023 21747 77051
rect 21437 76989 21747 77023
rect 21437 76961 21485 76989
rect 21513 76961 21547 76989
rect 21575 76961 21609 76989
rect 21637 76961 21671 76989
rect 21699 76961 21747 76989
rect 21437 68175 21747 76961
rect 21437 68147 21485 68175
rect 21513 68147 21547 68175
rect 21575 68147 21609 68175
rect 21637 68147 21671 68175
rect 21699 68147 21747 68175
rect 21437 68113 21747 68147
rect 21437 68085 21485 68113
rect 21513 68085 21547 68113
rect 21575 68085 21609 68113
rect 21637 68085 21671 68113
rect 21699 68085 21747 68113
rect 21437 68051 21747 68085
rect 21437 68023 21485 68051
rect 21513 68023 21547 68051
rect 21575 68023 21609 68051
rect 21637 68023 21671 68051
rect 21699 68023 21747 68051
rect 21437 67989 21747 68023
rect 21437 67961 21485 67989
rect 21513 67961 21547 67989
rect 21575 67961 21609 67989
rect 21637 67961 21671 67989
rect 21699 67961 21747 67989
rect 21437 59175 21747 67961
rect 21437 59147 21485 59175
rect 21513 59147 21547 59175
rect 21575 59147 21609 59175
rect 21637 59147 21671 59175
rect 21699 59147 21747 59175
rect 21437 59113 21747 59147
rect 21437 59085 21485 59113
rect 21513 59085 21547 59113
rect 21575 59085 21609 59113
rect 21637 59085 21671 59113
rect 21699 59085 21747 59113
rect 21437 59051 21747 59085
rect 21437 59023 21485 59051
rect 21513 59023 21547 59051
rect 21575 59023 21609 59051
rect 21637 59023 21671 59051
rect 21699 59023 21747 59051
rect 21437 58989 21747 59023
rect 21437 58961 21485 58989
rect 21513 58961 21547 58989
rect 21575 58961 21609 58989
rect 21637 58961 21671 58989
rect 21699 58961 21747 58989
rect 21437 50175 21747 58961
rect 21437 50147 21485 50175
rect 21513 50147 21547 50175
rect 21575 50147 21609 50175
rect 21637 50147 21671 50175
rect 21699 50147 21747 50175
rect 21437 50113 21747 50147
rect 21437 50085 21485 50113
rect 21513 50085 21547 50113
rect 21575 50085 21609 50113
rect 21637 50085 21671 50113
rect 21699 50085 21747 50113
rect 21437 50051 21747 50085
rect 21437 50023 21485 50051
rect 21513 50023 21547 50051
rect 21575 50023 21609 50051
rect 21637 50023 21671 50051
rect 21699 50023 21747 50051
rect 21437 49989 21747 50023
rect 21437 49961 21485 49989
rect 21513 49961 21547 49989
rect 21575 49961 21609 49989
rect 21637 49961 21671 49989
rect 21699 49961 21747 49989
rect 21437 41175 21747 49961
rect 21437 41147 21485 41175
rect 21513 41147 21547 41175
rect 21575 41147 21609 41175
rect 21637 41147 21671 41175
rect 21699 41147 21747 41175
rect 21437 41113 21747 41147
rect 21437 41085 21485 41113
rect 21513 41085 21547 41113
rect 21575 41085 21609 41113
rect 21637 41085 21671 41113
rect 21699 41085 21747 41113
rect 21437 41051 21747 41085
rect 21437 41023 21485 41051
rect 21513 41023 21547 41051
rect 21575 41023 21609 41051
rect 21637 41023 21671 41051
rect 21699 41023 21747 41051
rect 21437 40989 21747 41023
rect 21437 40961 21485 40989
rect 21513 40961 21547 40989
rect 21575 40961 21609 40989
rect 21637 40961 21671 40989
rect 21699 40961 21747 40989
rect 21437 32175 21747 40961
rect 21437 32147 21485 32175
rect 21513 32147 21547 32175
rect 21575 32147 21609 32175
rect 21637 32147 21671 32175
rect 21699 32147 21747 32175
rect 21437 32113 21747 32147
rect 21437 32085 21485 32113
rect 21513 32085 21547 32113
rect 21575 32085 21609 32113
rect 21637 32085 21671 32113
rect 21699 32085 21747 32113
rect 21437 32051 21747 32085
rect 21437 32023 21485 32051
rect 21513 32023 21547 32051
rect 21575 32023 21609 32051
rect 21637 32023 21671 32051
rect 21699 32023 21747 32051
rect 21437 31989 21747 32023
rect 21437 31961 21485 31989
rect 21513 31961 21547 31989
rect 21575 31961 21609 31989
rect 21637 31961 21671 31989
rect 21699 31961 21747 31989
rect 21437 23175 21747 31961
rect 21437 23147 21485 23175
rect 21513 23147 21547 23175
rect 21575 23147 21609 23175
rect 21637 23147 21671 23175
rect 21699 23147 21747 23175
rect 21437 23113 21747 23147
rect 21437 23085 21485 23113
rect 21513 23085 21547 23113
rect 21575 23085 21609 23113
rect 21637 23085 21671 23113
rect 21699 23085 21747 23113
rect 21437 23051 21747 23085
rect 21437 23023 21485 23051
rect 21513 23023 21547 23051
rect 21575 23023 21609 23051
rect 21637 23023 21671 23051
rect 21699 23023 21747 23051
rect 21437 22989 21747 23023
rect 21437 22961 21485 22989
rect 21513 22961 21547 22989
rect 21575 22961 21609 22989
rect 21637 22961 21671 22989
rect 21699 22961 21747 22989
rect 21437 14175 21747 22961
rect 21437 14147 21485 14175
rect 21513 14147 21547 14175
rect 21575 14147 21609 14175
rect 21637 14147 21671 14175
rect 21699 14147 21747 14175
rect 21437 14113 21747 14147
rect 21437 14085 21485 14113
rect 21513 14085 21547 14113
rect 21575 14085 21609 14113
rect 21637 14085 21671 14113
rect 21699 14085 21747 14113
rect 21437 14051 21747 14085
rect 21437 14023 21485 14051
rect 21513 14023 21547 14051
rect 21575 14023 21609 14051
rect 21637 14023 21671 14051
rect 21699 14023 21747 14051
rect 21437 13989 21747 14023
rect 21437 13961 21485 13989
rect 21513 13961 21547 13989
rect 21575 13961 21609 13989
rect 21637 13961 21671 13989
rect 21699 13961 21747 13989
rect 21437 5175 21747 13961
rect 21437 5147 21485 5175
rect 21513 5147 21547 5175
rect 21575 5147 21609 5175
rect 21637 5147 21671 5175
rect 21699 5147 21747 5175
rect 21437 5113 21747 5147
rect 21437 5085 21485 5113
rect 21513 5085 21547 5113
rect 21575 5085 21609 5113
rect 21637 5085 21671 5113
rect 21699 5085 21747 5113
rect 21437 5051 21747 5085
rect 21437 5023 21485 5051
rect 21513 5023 21547 5051
rect 21575 5023 21609 5051
rect 21637 5023 21671 5051
rect 21699 5023 21747 5051
rect 21437 4989 21747 5023
rect 21437 4961 21485 4989
rect 21513 4961 21547 4989
rect 21575 4961 21609 4989
rect 21637 4961 21671 4989
rect 21699 4961 21747 4989
rect 21437 -560 21747 4961
rect 21437 -588 21485 -560
rect 21513 -588 21547 -560
rect 21575 -588 21609 -560
rect 21637 -588 21671 -560
rect 21699 -588 21747 -560
rect 21437 -622 21747 -588
rect 21437 -650 21485 -622
rect 21513 -650 21547 -622
rect 21575 -650 21609 -622
rect 21637 -650 21671 -622
rect 21699 -650 21747 -622
rect 21437 -684 21747 -650
rect 21437 -712 21485 -684
rect 21513 -712 21547 -684
rect 21575 -712 21609 -684
rect 21637 -712 21671 -684
rect 21699 -712 21747 -684
rect 21437 -746 21747 -712
rect 21437 -774 21485 -746
rect 21513 -774 21547 -746
rect 21575 -774 21609 -746
rect 21637 -774 21671 -746
rect 21699 -774 21747 -746
rect 21437 -822 21747 -774
rect 28577 298606 28887 299134
rect 28577 298578 28625 298606
rect 28653 298578 28687 298606
rect 28715 298578 28749 298606
rect 28777 298578 28811 298606
rect 28839 298578 28887 298606
rect 28577 298544 28887 298578
rect 28577 298516 28625 298544
rect 28653 298516 28687 298544
rect 28715 298516 28749 298544
rect 28777 298516 28811 298544
rect 28839 298516 28887 298544
rect 28577 298482 28887 298516
rect 28577 298454 28625 298482
rect 28653 298454 28687 298482
rect 28715 298454 28749 298482
rect 28777 298454 28811 298482
rect 28839 298454 28887 298482
rect 28577 298420 28887 298454
rect 28577 298392 28625 298420
rect 28653 298392 28687 298420
rect 28715 298392 28749 298420
rect 28777 298392 28811 298420
rect 28839 298392 28887 298420
rect 28577 290175 28887 298392
rect 28577 290147 28625 290175
rect 28653 290147 28687 290175
rect 28715 290147 28749 290175
rect 28777 290147 28811 290175
rect 28839 290147 28887 290175
rect 28577 290113 28887 290147
rect 28577 290085 28625 290113
rect 28653 290085 28687 290113
rect 28715 290085 28749 290113
rect 28777 290085 28811 290113
rect 28839 290085 28887 290113
rect 28577 290051 28887 290085
rect 28577 290023 28625 290051
rect 28653 290023 28687 290051
rect 28715 290023 28749 290051
rect 28777 290023 28811 290051
rect 28839 290023 28887 290051
rect 28577 289989 28887 290023
rect 28577 289961 28625 289989
rect 28653 289961 28687 289989
rect 28715 289961 28749 289989
rect 28777 289961 28811 289989
rect 28839 289961 28887 289989
rect 28577 281175 28887 289961
rect 28577 281147 28625 281175
rect 28653 281147 28687 281175
rect 28715 281147 28749 281175
rect 28777 281147 28811 281175
rect 28839 281147 28887 281175
rect 28577 281113 28887 281147
rect 28577 281085 28625 281113
rect 28653 281085 28687 281113
rect 28715 281085 28749 281113
rect 28777 281085 28811 281113
rect 28839 281085 28887 281113
rect 28577 281051 28887 281085
rect 28577 281023 28625 281051
rect 28653 281023 28687 281051
rect 28715 281023 28749 281051
rect 28777 281023 28811 281051
rect 28839 281023 28887 281051
rect 28577 280989 28887 281023
rect 28577 280961 28625 280989
rect 28653 280961 28687 280989
rect 28715 280961 28749 280989
rect 28777 280961 28811 280989
rect 28839 280961 28887 280989
rect 28577 272175 28887 280961
rect 28577 272147 28625 272175
rect 28653 272147 28687 272175
rect 28715 272147 28749 272175
rect 28777 272147 28811 272175
rect 28839 272147 28887 272175
rect 28577 272113 28887 272147
rect 28577 272085 28625 272113
rect 28653 272085 28687 272113
rect 28715 272085 28749 272113
rect 28777 272085 28811 272113
rect 28839 272085 28887 272113
rect 28577 272051 28887 272085
rect 28577 272023 28625 272051
rect 28653 272023 28687 272051
rect 28715 272023 28749 272051
rect 28777 272023 28811 272051
rect 28839 272023 28887 272051
rect 28577 271989 28887 272023
rect 28577 271961 28625 271989
rect 28653 271961 28687 271989
rect 28715 271961 28749 271989
rect 28777 271961 28811 271989
rect 28839 271961 28887 271989
rect 28577 263175 28887 271961
rect 28577 263147 28625 263175
rect 28653 263147 28687 263175
rect 28715 263147 28749 263175
rect 28777 263147 28811 263175
rect 28839 263147 28887 263175
rect 28577 263113 28887 263147
rect 28577 263085 28625 263113
rect 28653 263085 28687 263113
rect 28715 263085 28749 263113
rect 28777 263085 28811 263113
rect 28839 263085 28887 263113
rect 28577 263051 28887 263085
rect 28577 263023 28625 263051
rect 28653 263023 28687 263051
rect 28715 263023 28749 263051
rect 28777 263023 28811 263051
rect 28839 263023 28887 263051
rect 28577 262989 28887 263023
rect 28577 262961 28625 262989
rect 28653 262961 28687 262989
rect 28715 262961 28749 262989
rect 28777 262961 28811 262989
rect 28839 262961 28887 262989
rect 28577 254175 28887 262961
rect 28577 254147 28625 254175
rect 28653 254147 28687 254175
rect 28715 254147 28749 254175
rect 28777 254147 28811 254175
rect 28839 254147 28887 254175
rect 28577 254113 28887 254147
rect 28577 254085 28625 254113
rect 28653 254085 28687 254113
rect 28715 254085 28749 254113
rect 28777 254085 28811 254113
rect 28839 254085 28887 254113
rect 28577 254051 28887 254085
rect 28577 254023 28625 254051
rect 28653 254023 28687 254051
rect 28715 254023 28749 254051
rect 28777 254023 28811 254051
rect 28839 254023 28887 254051
rect 28577 253989 28887 254023
rect 28577 253961 28625 253989
rect 28653 253961 28687 253989
rect 28715 253961 28749 253989
rect 28777 253961 28811 253989
rect 28839 253961 28887 253989
rect 28577 245175 28887 253961
rect 28577 245147 28625 245175
rect 28653 245147 28687 245175
rect 28715 245147 28749 245175
rect 28777 245147 28811 245175
rect 28839 245147 28887 245175
rect 28577 245113 28887 245147
rect 28577 245085 28625 245113
rect 28653 245085 28687 245113
rect 28715 245085 28749 245113
rect 28777 245085 28811 245113
rect 28839 245085 28887 245113
rect 28577 245051 28887 245085
rect 28577 245023 28625 245051
rect 28653 245023 28687 245051
rect 28715 245023 28749 245051
rect 28777 245023 28811 245051
rect 28839 245023 28887 245051
rect 28577 244989 28887 245023
rect 28577 244961 28625 244989
rect 28653 244961 28687 244989
rect 28715 244961 28749 244989
rect 28777 244961 28811 244989
rect 28839 244961 28887 244989
rect 28577 236175 28887 244961
rect 28577 236147 28625 236175
rect 28653 236147 28687 236175
rect 28715 236147 28749 236175
rect 28777 236147 28811 236175
rect 28839 236147 28887 236175
rect 28577 236113 28887 236147
rect 28577 236085 28625 236113
rect 28653 236085 28687 236113
rect 28715 236085 28749 236113
rect 28777 236085 28811 236113
rect 28839 236085 28887 236113
rect 28577 236051 28887 236085
rect 28577 236023 28625 236051
rect 28653 236023 28687 236051
rect 28715 236023 28749 236051
rect 28777 236023 28811 236051
rect 28839 236023 28887 236051
rect 28577 235989 28887 236023
rect 28577 235961 28625 235989
rect 28653 235961 28687 235989
rect 28715 235961 28749 235989
rect 28777 235961 28811 235989
rect 28839 235961 28887 235989
rect 28577 227175 28887 235961
rect 28577 227147 28625 227175
rect 28653 227147 28687 227175
rect 28715 227147 28749 227175
rect 28777 227147 28811 227175
rect 28839 227147 28887 227175
rect 28577 227113 28887 227147
rect 28577 227085 28625 227113
rect 28653 227085 28687 227113
rect 28715 227085 28749 227113
rect 28777 227085 28811 227113
rect 28839 227085 28887 227113
rect 28577 227051 28887 227085
rect 28577 227023 28625 227051
rect 28653 227023 28687 227051
rect 28715 227023 28749 227051
rect 28777 227023 28811 227051
rect 28839 227023 28887 227051
rect 28577 226989 28887 227023
rect 28577 226961 28625 226989
rect 28653 226961 28687 226989
rect 28715 226961 28749 226989
rect 28777 226961 28811 226989
rect 28839 226961 28887 226989
rect 28577 218175 28887 226961
rect 28577 218147 28625 218175
rect 28653 218147 28687 218175
rect 28715 218147 28749 218175
rect 28777 218147 28811 218175
rect 28839 218147 28887 218175
rect 28577 218113 28887 218147
rect 28577 218085 28625 218113
rect 28653 218085 28687 218113
rect 28715 218085 28749 218113
rect 28777 218085 28811 218113
rect 28839 218085 28887 218113
rect 28577 218051 28887 218085
rect 28577 218023 28625 218051
rect 28653 218023 28687 218051
rect 28715 218023 28749 218051
rect 28777 218023 28811 218051
rect 28839 218023 28887 218051
rect 28577 217989 28887 218023
rect 28577 217961 28625 217989
rect 28653 217961 28687 217989
rect 28715 217961 28749 217989
rect 28777 217961 28811 217989
rect 28839 217961 28887 217989
rect 28577 209175 28887 217961
rect 28577 209147 28625 209175
rect 28653 209147 28687 209175
rect 28715 209147 28749 209175
rect 28777 209147 28811 209175
rect 28839 209147 28887 209175
rect 28577 209113 28887 209147
rect 28577 209085 28625 209113
rect 28653 209085 28687 209113
rect 28715 209085 28749 209113
rect 28777 209085 28811 209113
rect 28839 209085 28887 209113
rect 28577 209051 28887 209085
rect 28577 209023 28625 209051
rect 28653 209023 28687 209051
rect 28715 209023 28749 209051
rect 28777 209023 28811 209051
rect 28839 209023 28887 209051
rect 28577 208989 28887 209023
rect 28577 208961 28625 208989
rect 28653 208961 28687 208989
rect 28715 208961 28749 208989
rect 28777 208961 28811 208989
rect 28839 208961 28887 208989
rect 28577 200175 28887 208961
rect 28577 200147 28625 200175
rect 28653 200147 28687 200175
rect 28715 200147 28749 200175
rect 28777 200147 28811 200175
rect 28839 200147 28887 200175
rect 28577 200113 28887 200147
rect 28577 200085 28625 200113
rect 28653 200085 28687 200113
rect 28715 200085 28749 200113
rect 28777 200085 28811 200113
rect 28839 200085 28887 200113
rect 28577 200051 28887 200085
rect 28577 200023 28625 200051
rect 28653 200023 28687 200051
rect 28715 200023 28749 200051
rect 28777 200023 28811 200051
rect 28839 200023 28887 200051
rect 28577 199989 28887 200023
rect 28577 199961 28625 199989
rect 28653 199961 28687 199989
rect 28715 199961 28749 199989
rect 28777 199961 28811 199989
rect 28839 199961 28887 199989
rect 28577 191175 28887 199961
rect 28577 191147 28625 191175
rect 28653 191147 28687 191175
rect 28715 191147 28749 191175
rect 28777 191147 28811 191175
rect 28839 191147 28887 191175
rect 28577 191113 28887 191147
rect 28577 191085 28625 191113
rect 28653 191085 28687 191113
rect 28715 191085 28749 191113
rect 28777 191085 28811 191113
rect 28839 191085 28887 191113
rect 28577 191051 28887 191085
rect 28577 191023 28625 191051
rect 28653 191023 28687 191051
rect 28715 191023 28749 191051
rect 28777 191023 28811 191051
rect 28839 191023 28887 191051
rect 28577 190989 28887 191023
rect 28577 190961 28625 190989
rect 28653 190961 28687 190989
rect 28715 190961 28749 190989
rect 28777 190961 28811 190989
rect 28839 190961 28887 190989
rect 28577 182175 28887 190961
rect 28577 182147 28625 182175
rect 28653 182147 28687 182175
rect 28715 182147 28749 182175
rect 28777 182147 28811 182175
rect 28839 182147 28887 182175
rect 28577 182113 28887 182147
rect 28577 182085 28625 182113
rect 28653 182085 28687 182113
rect 28715 182085 28749 182113
rect 28777 182085 28811 182113
rect 28839 182085 28887 182113
rect 28577 182051 28887 182085
rect 28577 182023 28625 182051
rect 28653 182023 28687 182051
rect 28715 182023 28749 182051
rect 28777 182023 28811 182051
rect 28839 182023 28887 182051
rect 28577 181989 28887 182023
rect 28577 181961 28625 181989
rect 28653 181961 28687 181989
rect 28715 181961 28749 181989
rect 28777 181961 28811 181989
rect 28839 181961 28887 181989
rect 28577 173175 28887 181961
rect 28577 173147 28625 173175
rect 28653 173147 28687 173175
rect 28715 173147 28749 173175
rect 28777 173147 28811 173175
rect 28839 173147 28887 173175
rect 28577 173113 28887 173147
rect 28577 173085 28625 173113
rect 28653 173085 28687 173113
rect 28715 173085 28749 173113
rect 28777 173085 28811 173113
rect 28839 173085 28887 173113
rect 28577 173051 28887 173085
rect 28577 173023 28625 173051
rect 28653 173023 28687 173051
rect 28715 173023 28749 173051
rect 28777 173023 28811 173051
rect 28839 173023 28887 173051
rect 28577 172989 28887 173023
rect 28577 172961 28625 172989
rect 28653 172961 28687 172989
rect 28715 172961 28749 172989
rect 28777 172961 28811 172989
rect 28839 172961 28887 172989
rect 28577 164175 28887 172961
rect 28577 164147 28625 164175
rect 28653 164147 28687 164175
rect 28715 164147 28749 164175
rect 28777 164147 28811 164175
rect 28839 164147 28887 164175
rect 28577 164113 28887 164147
rect 28577 164085 28625 164113
rect 28653 164085 28687 164113
rect 28715 164085 28749 164113
rect 28777 164085 28811 164113
rect 28839 164085 28887 164113
rect 28577 164051 28887 164085
rect 28577 164023 28625 164051
rect 28653 164023 28687 164051
rect 28715 164023 28749 164051
rect 28777 164023 28811 164051
rect 28839 164023 28887 164051
rect 28577 163989 28887 164023
rect 28577 163961 28625 163989
rect 28653 163961 28687 163989
rect 28715 163961 28749 163989
rect 28777 163961 28811 163989
rect 28839 163961 28887 163989
rect 28577 155175 28887 163961
rect 28577 155147 28625 155175
rect 28653 155147 28687 155175
rect 28715 155147 28749 155175
rect 28777 155147 28811 155175
rect 28839 155147 28887 155175
rect 28577 155113 28887 155147
rect 28577 155085 28625 155113
rect 28653 155085 28687 155113
rect 28715 155085 28749 155113
rect 28777 155085 28811 155113
rect 28839 155085 28887 155113
rect 28577 155051 28887 155085
rect 28577 155023 28625 155051
rect 28653 155023 28687 155051
rect 28715 155023 28749 155051
rect 28777 155023 28811 155051
rect 28839 155023 28887 155051
rect 28577 154989 28887 155023
rect 28577 154961 28625 154989
rect 28653 154961 28687 154989
rect 28715 154961 28749 154989
rect 28777 154961 28811 154989
rect 28839 154961 28887 154989
rect 28577 146175 28887 154961
rect 28577 146147 28625 146175
rect 28653 146147 28687 146175
rect 28715 146147 28749 146175
rect 28777 146147 28811 146175
rect 28839 146147 28887 146175
rect 28577 146113 28887 146147
rect 28577 146085 28625 146113
rect 28653 146085 28687 146113
rect 28715 146085 28749 146113
rect 28777 146085 28811 146113
rect 28839 146085 28887 146113
rect 28577 146051 28887 146085
rect 28577 146023 28625 146051
rect 28653 146023 28687 146051
rect 28715 146023 28749 146051
rect 28777 146023 28811 146051
rect 28839 146023 28887 146051
rect 28577 145989 28887 146023
rect 28577 145961 28625 145989
rect 28653 145961 28687 145989
rect 28715 145961 28749 145989
rect 28777 145961 28811 145989
rect 28839 145961 28887 145989
rect 28577 137175 28887 145961
rect 28577 137147 28625 137175
rect 28653 137147 28687 137175
rect 28715 137147 28749 137175
rect 28777 137147 28811 137175
rect 28839 137147 28887 137175
rect 28577 137113 28887 137147
rect 28577 137085 28625 137113
rect 28653 137085 28687 137113
rect 28715 137085 28749 137113
rect 28777 137085 28811 137113
rect 28839 137085 28887 137113
rect 28577 137051 28887 137085
rect 28577 137023 28625 137051
rect 28653 137023 28687 137051
rect 28715 137023 28749 137051
rect 28777 137023 28811 137051
rect 28839 137023 28887 137051
rect 28577 136989 28887 137023
rect 28577 136961 28625 136989
rect 28653 136961 28687 136989
rect 28715 136961 28749 136989
rect 28777 136961 28811 136989
rect 28839 136961 28887 136989
rect 28577 128175 28887 136961
rect 28577 128147 28625 128175
rect 28653 128147 28687 128175
rect 28715 128147 28749 128175
rect 28777 128147 28811 128175
rect 28839 128147 28887 128175
rect 28577 128113 28887 128147
rect 28577 128085 28625 128113
rect 28653 128085 28687 128113
rect 28715 128085 28749 128113
rect 28777 128085 28811 128113
rect 28839 128085 28887 128113
rect 28577 128051 28887 128085
rect 28577 128023 28625 128051
rect 28653 128023 28687 128051
rect 28715 128023 28749 128051
rect 28777 128023 28811 128051
rect 28839 128023 28887 128051
rect 28577 127989 28887 128023
rect 28577 127961 28625 127989
rect 28653 127961 28687 127989
rect 28715 127961 28749 127989
rect 28777 127961 28811 127989
rect 28839 127961 28887 127989
rect 28577 119175 28887 127961
rect 28577 119147 28625 119175
rect 28653 119147 28687 119175
rect 28715 119147 28749 119175
rect 28777 119147 28811 119175
rect 28839 119147 28887 119175
rect 28577 119113 28887 119147
rect 28577 119085 28625 119113
rect 28653 119085 28687 119113
rect 28715 119085 28749 119113
rect 28777 119085 28811 119113
rect 28839 119085 28887 119113
rect 28577 119051 28887 119085
rect 28577 119023 28625 119051
rect 28653 119023 28687 119051
rect 28715 119023 28749 119051
rect 28777 119023 28811 119051
rect 28839 119023 28887 119051
rect 28577 118989 28887 119023
rect 28577 118961 28625 118989
rect 28653 118961 28687 118989
rect 28715 118961 28749 118989
rect 28777 118961 28811 118989
rect 28839 118961 28887 118989
rect 28577 110175 28887 118961
rect 28577 110147 28625 110175
rect 28653 110147 28687 110175
rect 28715 110147 28749 110175
rect 28777 110147 28811 110175
rect 28839 110147 28887 110175
rect 28577 110113 28887 110147
rect 28577 110085 28625 110113
rect 28653 110085 28687 110113
rect 28715 110085 28749 110113
rect 28777 110085 28811 110113
rect 28839 110085 28887 110113
rect 28577 110051 28887 110085
rect 28577 110023 28625 110051
rect 28653 110023 28687 110051
rect 28715 110023 28749 110051
rect 28777 110023 28811 110051
rect 28839 110023 28887 110051
rect 28577 109989 28887 110023
rect 28577 109961 28625 109989
rect 28653 109961 28687 109989
rect 28715 109961 28749 109989
rect 28777 109961 28811 109989
rect 28839 109961 28887 109989
rect 28577 101175 28887 109961
rect 28577 101147 28625 101175
rect 28653 101147 28687 101175
rect 28715 101147 28749 101175
rect 28777 101147 28811 101175
rect 28839 101147 28887 101175
rect 28577 101113 28887 101147
rect 28577 101085 28625 101113
rect 28653 101085 28687 101113
rect 28715 101085 28749 101113
rect 28777 101085 28811 101113
rect 28839 101085 28887 101113
rect 28577 101051 28887 101085
rect 28577 101023 28625 101051
rect 28653 101023 28687 101051
rect 28715 101023 28749 101051
rect 28777 101023 28811 101051
rect 28839 101023 28887 101051
rect 28577 100989 28887 101023
rect 28577 100961 28625 100989
rect 28653 100961 28687 100989
rect 28715 100961 28749 100989
rect 28777 100961 28811 100989
rect 28839 100961 28887 100989
rect 28577 92175 28887 100961
rect 28577 92147 28625 92175
rect 28653 92147 28687 92175
rect 28715 92147 28749 92175
rect 28777 92147 28811 92175
rect 28839 92147 28887 92175
rect 28577 92113 28887 92147
rect 28577 92085 28625 92113
rect 28653 92085 28687 92113
rect 28715 92085 28749 92113
rect 28777 92085 28811 92113
rect 28839 92085 28887 92113
rect 28577 92051 28887 92085
rect 28577 92023 28625 92051
rect 28653 92023 28687 92051
rect 28715 92023 28749 92051
rect 28777 92023 28811 92051
rect 28839 92023 28887 92051
rect 28577 91989 28887 92023
rect 28577 91961 28625 91989
rect 28653 91961 28687 91989
rect 28715 91961 28749 91989
rect 28777 91961 28811 91989
rect 28839 91961 28887 91989
rect 28577 83175 28887 91961
rect 28577 83147 28625 83175
rect 28653 83147 28687 83175
rect 28715 83147 28749 83175
rect 28777 83147 28811 83175
rect 28839 83147 28887 83175
rect 28577 83113 28887 83147
rect 28577 83085 28625 83113
rect 28653 83085 28687 83113
rect 28715 83085 28749 83113
rect 28777 83085 28811 83113
rect 28839 83085 28887 83113
rect 28577 83051 28887 83085
rect 28577 83023 28625 83051
rect 28653 83023 28687 83051
rect 28715 83023 28749 83051
rect 28777 83023 28811 83051
rect 28839 83023 28887 83051
rect 28577 82989 28887 83023
rect 28577 82961 28625 82989
rect 28653 82961 28687 82989
rect 28715 82961 28749 82989
rect 28777 82961 28811 82989
rect 28839 82961 28887 82989
rect 28577 74175 28887 82961
rect 28577 74147 28625 74175
rect 28653 74147 28687 74175
rect 28715 74147 28749 74175
rect 28777 74147 28811 74175
rect 28839 74147 28887 74175
rect 28577 74113 28887 74147
rect 28577 74085 28625 74113
rect 28653 74085 28687 74113
rect 28715 74085 28749 74113
rect 28777 74085 28811 74113
rect 28839 74085 28887 74113
rect 28577 74051 28887 74085
rect 28577 74023 28625 74051
rect 28653 74023 28687 74051
rect 28715 74023 28749 74051
rect 28777 74023 28811 74051
rect 28839 74023 28887 74051
rect 28577 73989 28887 74023
rect 28577 73961 28625 73989
rect 28653 73961 28687 73989
rect 28715 73961 28749 73989
rect 28777 73961 28811 73989
rect 28839 73961 28887 73989
rect 28577 65175 28887 73961
rect 28577 65147 28625 65175
rect 28653 65147 28687 65175
rect 28715 65147 28749 65175
rect 28777 65147 28811 65175
rect 28839 65147 28887 65175
rect 28577 65113 28887 65147
rect 28577 65085 28625 65113
rect 28653 65085 28687 65113
rect 28715 65085 28749 65113
rect 28777 65085 28811 65113
rect 28839 65085 28887 65113
rect 28577 65051 28887 65085
rect 28577 65023 28625 65051
rect 28653 65023 28687 65051
rect 28715 65023 28749 65051
rect 28777 65023 28811 65051
rect 28839 65023 28887 65051
rect 28577 64989 28887 65023
rect 28577 64961 28625 64989
rect 28653 64961 28687 64989
rect 28715 64961 28749 64989
rect 28777 64961 28811 64989
rect 28839 64961 28887 64989
rect 28577 56175 28887 64961
rect 28577 56147 28625 56175
rect 28653 56147 28687 56175
rect 28715 56147 28749 56175
rect 28777 56147 28811 56175
rect 28839 56147 28887 56175
rect 28577 56113 28887 56147
rect 28577 56085 28625 56113
rect 28653 56085 28687 56113
rect 28715 56085 28749 56113
rect 28777 56085 28811 56113
rect 28839 56085 28887 56113
rect 28577 56051 28887 56085
rect 28577 56023 28625 56051
rect 28653 56023 28687 56051
rect 28715 56023 28749 56051
rect 28777 56023 28811 56051
rect 28839 56023 28887 56051
rect 28577 55989 28887 56023
rect 28577 55961 28625 55989
rect 28653 55961 28687 55989
rect 28715 55961 28749 55989
rect 28777 55961 28811 55989
rect 28839 55961 28887 55989
rect 28577 47175 28887 55961
rect 28577 47147 28625 47175
rect 28653 47147 28687 47175
rect 28715 47147 28749 47175
rect 28777 47147 28811 47175
rect 28839 47147 28887 47175
rect 28577 47113 28887 47147
rect 28577 47085 28625 47113
rect 28653 47085 28687 47113
rect 28715 47085 28749 47113
rect 28777 47085 28811 47113
rect 28839 47085 28887 47113
rect 28577 47051 28887 47085
rect 28577 47023 28625 47051
rect 28653 47023 28687 47051
rect 28715 47023 28749 47051
rect 28777 47023 28811 47051
rect 28839 47023 28887 47051
rect 28577 46989 28887 47023
rect 28577 46961 28625 46989
rect 28653 46961 28687 46989
rect 28715 46961 28749 46989
rect 28777 46961 28811 46989
rect 28839 46961 28887 46989
rect 28577 38175 28887 46961
rect 28577 38147 28625 38175
rect 28653 38147 28687 38175
rect 28715 38147 28749 38175
rect 28777 38147 28811 38175
rect 28839 38147 28887 38175
rect 28577 38113 28887 38147
rect 28577 38085 28625 38113
rect 28653 38085 28687 38113
rect 28715 38085 28749 38113
rect 28777 38085 28811 38113
rect 28839 38085 28887 38113
rect 28577 38051 28887 38085
rect 28577 38023 28625 38051
rect 28653 38023 28687 38051
rect 28715 38023 28749 38051
rect 28777 38023 28811 38051
rect 28839 38023 28887 38051
rect 28577 37989 28887 38023
rect 28577 37961 28625 37989
rect 28653 37961 28687 37989
rect 28715 37961 28749 37989
rect 28777 37961 28811 37989
rect 28839 37961 28887 37989
rect 28577 29175 28887 37961
rect 28577 29147 28625 29175
rect 28653 29147 28687 29175
rect 28715 29147 28749 29175
rect 28777 29147 28811 29175
rect 28839 29147 28887 29175
rect 28577 29113 28887 29147
rect 28577 29085 28625 29113
rect 28653 29085 28687 29113
rect 28715 29085 28749 29113
rect 28777 29085 28811 29113
rect 28839 29085 28887 29113
rect 28577 29051 28887 29085
rect 28577 29023 28625 29051
rect 28653 29023 28687 29051
rect 28715 29023 28749 29051
rect 28777 29023 28811 29051
rect 28839 29023 28887 29051
rect 28577 28989 28887 29023
rect 28577 28961 28625 28989
rect 28653 28961 28687 28989
rect 28715 28961 28749 28989
rect 28777 28961 28811 28989
rect 28839 28961 28887 28989
rect 28577 20175 28887 28961
rect 28577 20147 28625 20175
rect 28653 20147 28687 20175
rect 28715 20147 28749 20175
rect 28777 20147 28811 20175
rect 28839 20147 28887 20175
rect 28577 20113 28887 20147
rect 28577 20085 28625 20113
rect 28653 20085 28687 20113
rect 28715 20085 28749 20113
rect 28777 20085 28811 20113
rect 28839 20085 28887 20113
rect 28577 20051 28887 20085
rect 28577 20023 28625 20051
rect 28653 20023 28687 20051
rect 28715 20023 28749 20051
rect 28777 20023 28811 20051
rect 28839 20023 28887 20051
rect 28577 19989 28887 20023
rect 28577 19961 28625 19989
rect 28653 19961 28687 19989
rect 28715 19961 28749 19989
rect 28777 19961 28811 19989
rect 28839 19961 28887 19989
rect 28577 11175 28887 19961
rect 28577 11147 28625 11175
rect 28653 11147 28687 11175
rect 28715 11147 28749 11175
rect 28777 11147 28811 11175
rect 28839 11147 28887 11175
rect 28577 11113 28887 11147
rect 28577 11085 28625 11113
rect 28653 11085 28687 11113
rect 28715 11085 28749 11113
rect 28777 11085 28811 11113
rect 28839 11085 28887 11113
rect 28577 11051 28887 11085
rect 28577 11023 28625 11051
rect 28653 11023 28687 11051
rect 28715 11023 28749 11051
rect 28777 11023 28811 11051
rect 28839 11023 28887 11051
rect 28577 10989 28887 11023
rect 28577 10961 28625 10989
rect 28653 10961 28687 10989
rect 28715 10961 28749 10989
rect 28777 10961 28811 10989
rect 28839 10961 28887 10989
rect 28577 2175 28887 10961
rect 28577 2147 28625 2175
rect 28653 2147 28687 2175
rect 28715 2147 28749 2175
rect 28777 2147 28811 2175
rect 28839 2147 28887 2175
rect 28577 2113 28887 2147
rect 28577 2085 28625 2113
rect 28653 2085 28687 2113
rect 28715 2085 28749 2113
rect 28777 2085 28811 2113
rect 28839 2085 28887 2113
rect 28577 2051 28887 2085
rect 28577 2023 28625 2051
rect 28653 2023 28687 2051
rect 28715 2023 28749 2051
rect 28777 2023 28811 2051
rect 28839 2023 28887 2051
rect 28577 1989 28887 2023
rect 28577 1961 28625 1989
rect 28653 1961 28687 1989
rect 28715 1961 28749 1989
rect 28777 1961 28811 1989
rect 28839 1961 28887 1989
rect 28577 -80 28887 1961
rect 28577 -108 28625 -80
rect 28653 -108 28687 -80
rect 28715 -108 28749 -80
rect 28777 -108 28811 -80
rect 28839 -108 28887 -80
rect 28577 -142 28887 -108
rect 28577 -170 28625 -142
rect 28653 -170 28687 -142
rect 28715 -170 28749 -142
rect 28777 -170 28811 -142
rect 28839 -170 28887 -142
rect 28577 -204 28887 -170
rect 28577 -232 28625 -204
rect 28653 -232 28687 -204
rect 28715 -232 28749 -204
rect 28777 -232 28811 -204
rect 28839 -232 28887 -204
rect 28577 -266 28887 -232
rect 28577 -294 28625 -266
rect 28653 -294 28687 -266
rect 28715 -294 28749 -266
rect 28777 -294 28811 -266
rect 28839 -294 28887 -266
rect 28577 -822 28887 -294
rect 30437 299086 30747 299134
rect 30437 299058 30485 299086
rect 30513 299058 30547 299086
rect 30575 299058 30609 299086
rect 30637 299058 30671 299086
rect 30699 299058 30747 299086
rect 30437 299024 30747 299058
rect 30437 298996 30485 299024
rect 30513 298996 30547 299024
rect 30575 298996 30609 299024
rect 30637 298996 30671 299024
rect 30699 298996 30747 299024
rect 30437 298962 30747 298996
rect 30437 298934 30485 298962
rect 30513 298934 30547 298962
rect 30575 298934 30609 298962
rect 30637 298934 30671 298962
rect 30699 298934 30747 298962
rect 30437 298900 30747 298934
rect 30437 298872 30485 298900
rect 30513 298872 30547 298900
rect 30575 298872 30609 298900
rect 30637 298872 30671 298900
rect 30699 298872 30747 298900
rect 30437 293175 30747 298872
rect 30437 293147 30485 293175
rect 30513 293147 30547 293175
rect 30575 293147 30609 293175
rect 30637 293147 30671 293175
rect 30699 293147 30747 293175
rect 30437 293113 30747 293147
rect 30437 293085 30485 293113
rect 30513 293085 30547 293113
rect 30575 293085 30609 293113
rect 30637 293085 30671 293113
rect 30699 293085 30747 293113
rect 30437 293051 30747 293085
rect 30437 293023 30485 293051
rect 30513 293023 30547 293051
rect 30575 293023 30609 293051
rect 30637 293023 30671 293051
rect 30699 293023 30747 293051
rect 30437 292989 30747 293023
rect 30437 292961 30485 292989
rect 30513 292961 30547 292989
rect 30575 292961 30609 292989
rect 30637 292961 30671 292989
rect 30699 292961 30747 292989
rect 30437 284175 30747 292961
rect 30437 284147 30485 284175
rect 30513 284147 30547 284175
rect 30575 284147 30609 284175
rect 30637 284147 30671 284175
rect 30699 284147 30747 284175
rect 30437 284113 30747 284147
rect 30437 284085 30485 284113
rect 30513 284085 30547 284113
rect 30575 284085 30609 284113
rect 30637 284085 30671 284113
rect 30699 284085 30747 284113
rect 30437 284051 30747 284085
rect 30437 284023 30485 284051
rect 30513 284023 30547 284051
rect 30575 284023 30609 284051
rect 30637 284023 30671 284051
rect 30699 284023 30747 284051
rect 30437 283989 30747 284023
rect 30437 283961 30485 283989
rect 30513 283961 30547 283989
rect 30575 283961 30609 283989
rect 30637 283961 30671 283989
rect 30699 283961 30747 283989
rect 30437 275175 30747 283961
rect 30437 275147 30485 275175
rect 30513 275147 30547 275175
rect 30575 275147 30609 275175
rect 30637 275147 30671 275175
rect 30699 275147 30747 275175
rect 30437 275113 30747 275147
rect 30437 275085 30485 275113
rect 30513 275085 30547 275113
rect 30575 275085 30609 275113
rect 30637 275085 30671 275113
rect 30699 275085 30747 275113
rect 30437 275051 30747 275085
rect 30437 275023 30485 275051
rect 30513 275023 30547 275051
rect 30575 275023 30609 275051
rect 30637 275023 30671 275051
rect 30699 275023 30747 275051
rect 30437 274989 30747 275023
rect 30437 274961 30485 274989
rect 30513 274961 30547 274989
rect 30575 274961 30609 274989
rect 30637 274961 30671 274989
rect 30699 274961 30747 274989
rect 30437 266175 30747 274961
rect 30437 266147 30485 266175
rect 30513 266147 30547 266175
rect 30575 266147 30609 266175
rect 30637 266147 30671 266175
rect 30699 266147 30747 266175
rect 30437 266113 30747 266147
rect 30437 266085 30485 266113
rect 30513 266085 30547 266113
rect 30575 266085 30609 266113
rect 30637 266085 30671 266113
rect 30699 266085 30747 266113
rect 30437 266051 30747 266085
rect 30437 266023 30485 266051
rect 30513 266023 30547 266051
rect 30575 266023 30609 266051
rect 30637 266023 30671 266051
rect 30699 266023 30747 266051
rect 30437 265989 30747 266023
rect 30437 265961 30485 265989
rect 30513 265961 30547 265989
rect 30575 265961 30609 265989
rect 30637 265961 30671 265989
rect 30699 265961 30747 265989
rect 30437 257175 30747 265961
rect 30437 257147 30485 257175
rect 30513 257147 30547 257175
rect 30575 257147 30609 257175
rect 30637 257147 30671 257175
rect 30699 257147 30747 257175
rect 30437 257113 30747 257147
rect 30437 257085 30485 257113
rect 30513 257085 30547 257113
rect 30575 257085 30609 257113
rect 30637 257085 30671 257113
rect 30699 257085 30747 257113
rect 30437 257051 30747 257085
rect 30437 257023 30485 257051
rect 30513 257023 30547 257051
rect 30575 257023 30609 257051
rect 30637 257023 30671 257051
rect 30699 257023 30747 257051
rect 30437 256989 30747 257023
rect 30437 256961 30485 256989
rect 30513 256961 30547 256989
rect 30575 256961 30609 256989
rect 30637 256961 30671 256989
rect 30699 256961 30747 256989
rect 30437 248175 30747 256961
rect 30437 248147 30485 248175
rect 30513 248147 30547 248175
rect 30575 248147 30609 248175
rect 30637 248147 30671 248175
rect 30699 248147 30747 248175
rect 30437 248113 30747 248147
rect 30437 248085 30485 248113
rect 30513 248085 30547 248113
rect 30575 248085 30609 248113
rect 30637 248085 30671 248113
rect 30699 248085 30747 248113
rect 30437 248051 30747 248085
rect 30437 248023 30485 248051
rect 30513 248023 30547 248051
rect 30575 248023 30609 248051
rect 30637 248023 30671 248051
rect 30699 248023 30747 248051
rect 30437 247989 30747 248023
rect 30437 247961 30485 247989
rect 30513 247961 30547 247989
rect 30575 247961 30609 247989
rect 30637 247961 30671 247989
rect 30699 247961 30747 247989
rect 30437 239175 30747 247961
rect 30437 239147 30485 239175
rect 30513 239147 30547 239175
rect 30575 239147 30609 239175
rect 30637 239147 30671 239175
rect 30699 239147 30747 239175
rect 30437 239113 30747 239147
rect 30437 239085 30485 239113
rect 30513 239085 30547 239113
rect 30575 239085 30609 239113
rect 30637 239085 30671 239113
rect 30699 239085 30747 239113
rect 30437 239051 30747 239085
rect 30437 239023 30485 239051
rect 30513 239023 30547 239051
rect 30575 239023 30609 239051
rect 30637 239023 30671 239051
rect 30699 239023 30747 239051
rect 30437 238989 30747 239023
rect 30437 238961 30485 238989
rect 30513 238961 30547 238989
rect 30575 238961 30609 238989
rect 30637 238961 30671 238989
rect 30699 238961 30747 238989
rect 30437 230175 30747 238961
rect 30437 230147 30485 230175
rect 30513 230147 30547 230175
rect 30575 230147 30609 230175
rect 30637 230147 30671 230175
rect 30699 230147 30747 230175
rect 30437 230113 30747 230147
rect 30437 230085 30485 230113
rect 30513 230085 30547 230113
rect 30575 230085 30609 230113
rect 30637 230085 30671 230113
rect 30699 230085 30747 230113
rect 30437 230051 30747 230085
rect 30437 230023 30485 230051
rect 30513 230023 30547 230051
rect 30575 230023 30609 230051
rect 30637 230023 30671 230051
rect 30699 230023 30747 230051
rect 30437 229989 30747 230023
rect 30437 229961 30485 229989
rect 30513 229961 30547 229989
rect 30575 229961 30609 229989
rect 30637 229961 30671 229989
rect 30699 229961 30747 229989
rect 30437 221175 30747 229961
rect 30437 221147 30485 221175
rect 30513 221147 30547 221175
rect 30575 221147 30609 221175
rect 30637 221147 30671 221175
rect 30699 221147 30747 221175
rect 30437 221113 30747 221147
rect 30437 221085 30485 221113
rect 30513 221085 30547 221113
rect 30575 221085 30609 221113
rect 30637 221085 30671 221113
rect 30699 221085 30747 221113
rect 30437 221051 30747 221085
rect 30437 221023 30485 221051
rect 30513 221023 30547 221051
rect 30575 221023 30609 221051
rect 30637 221023 30671 221051
rect 30699 221023 30747 221051
rect 30437 220989 30747 221023
rect 30437 220961 30485 220989
rect 30513 220961 30547 220989
rect 30575 220961 30609 220989
rect 30637 220961 30671 220989
rect 30699 220961 30747 220989
rect 30437 212175 30747 220961
rect 30437 212147 30485 212175
rect 30513 212147 30547 212175
rect 30575 212147 30609 212175
rect 30637 212147 30671 212175
rect 30699 212147 30747 212175
rect 30437 212113 30747 212147
rect 30437 212085 30485 212113
rect 30513 212085 30547 212113
rect 30575 212085 30609 212113
rect 30637 212085 30671 212113
rect 30699 212085 30747 212113
rect 30437 212051 30747 212085
rect 30437 212023 30485 212051
rect 30513 212023 30547 212051
rect 30575 212023 30609 212051
rect 30637 212023 30671 212051
rect 30699 212023 30747 212051
rect 30437 211989 30747 212023
rect 30437 211961 30485 211989
rect 30513 211961 30547 211989
rect 30575 211961 30609 211989
rect 30637 211961 30671 211989
rect 30699 211961 30747 211989
rect 30437 203175 30747 211961
rect 30437 203147 30485 203175
rect 30513 203147 30547 203175
rect 30575 203147 30609 203175
rect 30637 203147 30671 203175
rect 30699 203147 30747 203175
rect 30437 203113 30747 203147
rect 30437 203085 30485 203113
rect 30513 203085 30547 203113
rect 30575 203085 30609 203113
rect 30637 203085 30671 203113
rect 30699 203085 30747 203113
rect 30437 203051 30747 203085
rect 30437 203023 30485 203051
rect 30513 203023 30547 203051
rect 30575 203023 30609 203051
rect 30637 203023 30671 203051
rect 30699 203023 30747 203051
rect 30437 202989 30747 203023
rect 30437 202961 30485 202989
rect 30513 202961 30547 202989
rect 30575 202961 30609 202989
rect 30637 202961 30671 202989
rect 30699 202961 30747 202989
rect 30437 194175 30747 202961
rect 30437 194147 30485 194175
rect 30513 194147 30547 194175
rect 30575 194147 30609 194175
rect 30637 194147 30671 194175
rect 30699 194147 30747 194175
rect 30437 194113 30747 194147
rect 30437 194085 30485 194113
rect 30513 194085 30547 194113
rect 30575 194085 30609 194113
rect 30637 194085 30671 194113
rect 30699 194085 30747 194113
rect 30437 194051 30747 194085
rect 30437 194023 30485 194051
rect 30513 194023 30547 194051
rect 30575 194023 30609 194051
rect 30637 194023 30671 194051
rect 30699 194023 30747 194051
rect 30437 193989 30747 194023
rect 30437 193961 30485 193989
rect 30513 193961 30547 193989
rect 30575 193961 30609 193989
rect 30637 193961 30671 193989
rect 30699 193961 30747 193989
rect 30437 185175 30747 193961
rect 30437 185147 30485 185175
rect 30513 185147 30547 185175
rect 30575 185147 30609 185175
rect 30637 185147 30671 185175
rect 30699 185147 30747 185175
rect 30437 185113 30747 185147
rect 30437 185085 30485 185113
rect 30513 185085 30547 185113
rect 30575 185085 30609 185113
rect 30637 185085 30671 185113
rect 30699 185085 30747 185113
rect 30437 185051 30747 185085
rect 30437 185023 30485 185051
rect 30513 185023 30547 185051
rect 30575 185023 30609 185051
rect 30637 185023 30671 185051
rect 30699 185023 30747 185051
rect 30437 184989 30747 185023
rect 30437 184961 30485 184989
rect 30513 184961 30547 184989
rect 30575 184961 30609 184989
rect 30637 184961 30671 184989
rect 30699 184961 30747 184989
rect 30437 176175 30747 184961
rect 30437 176147 30485 176175
rect 30513 176147 30547 176175
rect 30575 176147 30609 176175
rect 30637 176147 30671 176175
rect 30699 176147 30747 176175
rect 30437 176113 30747 176147
rect 30437 176085 30485 176113
rect 30513 176085 30547 176113
rect 30575 176085 30609 176113
rect 30637 176085 30671 176113
rect 30699 176085 30747 176113
rect 30437 176051 30747 176085
rect 30437 176023 30485 176051
rect 30513 176023 30547 176051
rect 30575 176023 30609 176051
rect 30637 176023 30671 176051
rect 30699 176023 30747 176051
rect 30437 175989 30747 176023
rect 30437 175961 30485 175989
rect 30513 175961 30547 175989
rect 30575 175961 30609 175989
rect 30637 175961 30671 175989
rect 30699 175961 30747 175989
rect 30437 167175 30747 175961
rect 30437 167147 30485 167175
rect 30513 167147 30547 167175
rect 30575 167147 30609 167175
rect 30637 167147 30671 167175
rect 30699 167147 30747 167175
rect 30437 167113 30747 167147
rect 30437 167085 30485 167113
rect 30513 167085 30547 167113
rect 30575 167085 30609 167113
rect 30637 167085 30671 167113
rect 30699 167085 30747 167113
rect 30437 167051 30747 167085
rect 30437 167023 30485 167051
rect 30513 167023 30547 167051
rect 30575 167023 30609 167051
rect 30637 167023 30671 167051
rect 30699 167023 30747 167051
rect 30437 166989 30747 167023
rect 30437 166961 30485 166989
rect 30513 166961 30547 166989
rect 30575 166961 30609 166989
rect 30637 166961 30671 166989
rect 30699 166961 30747 166989
rect 30437 158175 30747 166961
rect 30437 158147 30485 158175
rect 30513 158147 30547 158175
rect 30575 158147 30609 158175
rect 30637 158147 30671 158175
rect 30699 158147 30747 158175
rect 30437 158113 30747 158147
rect 30437 158085 30485 158113
rect 30513 158085 30547 158113
rect 30575 158085 30609 158113
rect 30637 158085 30671 158113
rect 30699 158085 30747 158113
rect 30437 158051 30747 158085
rect 30437 158023 30485 158051
rect 30513 158023 30547 158051
rect 30575 158023 30609 158051
rect 30637 158023 30671 158051
rect 30699 158023 30747 158051
rect 30437 157989 30747 158023
rect 30437 157961 30485 157989
rect 30513 157961 30547 157989
rect 30575 157961 30609 157989
rect 30637 157961 30671 157989
rect 30699 157961 30747 157989
rect 30437 149175 30747 157961
rect 30437 149147 30485 149175
rect 30513 149147 30547 149175
rect 30575 149147 30609 149175
rect 30637 149147 30671 149175
rect 30699 149147 30747 149175
rect 30437 149113 30747 149147
rect 30437 149085 30485 149113
rect 30513 149085 30547 149113
rect 30575 149085 30609 149113
rect 30637 149085 30671 149113
rect 30699 149085 30747 149113
rect 30437 149051 30747 149085
rect 30437 149023 30485 149051
rect 30513 149023 30547 149051
rect 30575 149023 30609 149051
rect 30637 149023 30671 149051
rect 30699 149023 30747 149051
rect 30437 148989 30747 149023
rect 30437 148961 30485 148989
rect 30513 148961 30547 148989
rect 30575 148961 30609 148989
rect 30637 148961 30671 148989
rect 30699 148961 30747 148989
rect 30437 140175 30747 148961
rect 30437 140147 30485 140175
rect 30513 140147 30547 140175
rect 30575 140147 30609 140175
rect 30637 140147 30671 140175
rect 30699 140147 30747 140175
rect 30437 140113 30747 140147
rect 30437 140085 30485 140113
rect 30513 140085 30547 140113
rect 30575 140085 30609 140113
rect 30637 140085 30671 140113
rect 30699 140085 30747 140113
rect 30437 140051 30747 140085
rect 30437 140023 30485 140051
rect 30513 140023 30547 140051
rect 30575 140023 30609 140051
rect 30637 140023 30671 140051
rect 30699 140023 30747 140051
rect 30437 139989 30747 140023
rect 30437 139961 30485 139989
rect 30513 139961 30547 139989
rect 30575 139961 30609 139989
rect 30637 139961 30671 139989
rect 30699 139961 30747 139989
rect 30437 131175 30747 139961
rect 30437 131147 30485 131175
rect 30513 131147 30547 131175
rect 30575 131147 30609 131175
rect 30637 131147 30671 131175
rect 30699 131147 30747 131175
rect 30437 131113 30747 131147
rect 30437 131085 30485 131113
rect 30513 131085 30547 131113
rect 30575 131085 30609 131113
rect 30637 131085 30671 131113
rect 30699 131085 30747 131113
rect 30437 131051 30747 131085
rect 30437 131023 30485 131051
rect 30513 131023 30547 131051
rect 30575 131023 30609 131051
rect 30637 131023 30671 131051
rect 30699 131023 30747 131051
rect 30437 130989 30747 131023
rect 30437 130961 30485 130989
rect 30513 130961 30547 130989
rect 30575 130961 30609 130989
rect 30637 130961 30671 130989
rect 30699 130961 30747 130989
rect 30437 122175 30747 130961
rect 30437 122147 30485 122175
rect 30513 122147 30547 122175
rect 30575 122147 30609 122175
rect 30637 122147 30671 122175
rect 30699 122147 30747 122175
rect 30437 122113 30747 122147
rect 30437 122085 30485 122113
rect 30513 122085 30547 122113
rect 30575 122085 30609 122113
rect 30637 122085 30671 122113
rect 30699 122085 30747 122113
rect 30437 122051 30747 122085
rect 30437 122023 30485 122051
rect 30513 122023 30547 122051
rect 30575 122023 30609 122051
rect 30637 122023 30671 122051
rect 30699 122023 30747 122051
rect 30437 121989 30747 122023
rect 30437 121961 30485 121989
rect 30513 121961 30547 121989
rect 30575 121961 30609 121989
rect 30637 121961 30671 121989
rect 30699 121961 30747 121989
rect 30437 113175 30747 121961
rect 30437 113147 30485 113175
rect 30513 113147 30547 113175
rect 30575 113147 30609 113175
rect 30637 113147 30671 113175
rect 30699 113147 30747 113175
rect 30437 113113 30747 113147
rect 30437 113085 30485 113113
rect 30513 113085 30547 113113
rect 30575 113085 30609 113113
rect 30637 113085 30671 113113
rect 30699 113085 30747 113113
rect 30437 113051 30747 113085
rect 30437 113023 30485 113051
rect 30513 113023 30547 113051
rect 30575 113023 30609 113051
rect 30637 113023 30671 113051
rect 30699 113023 30747 113051
rect 30437 112989 30747 113023
rect 30437 112961 30485 112989
rect 30513 112961 30547 112989
rect 30575 112961 30609 112989
rect 30637 112961 30671 112989
rect 30699 112961 30747 112989
rect 30437 104175 30747 112961
rect 30437 104147 30485 104175
rect 30513 104147 30547 104175
rect 30575 104147 30609 104175
rect 30637 104147 30671 104175
rect 30699 104147 30747 104175
rect 30437 104113 30747 104147
rect 30437 104085 30485 104113
rect 30513 104085 30547 104113
rect 30575 104085 30609 104113
rect 30637 104085 30671 104113
rect 30699 104085 30747 104113
rect 30437 104051 30747 104085
rect 30437 104023 30485 104051
rect 30513 104023 30547 104051
rect 30575 104023 30609 104051
rect 30637 104023 30671 104051
rect 30699 104023 30747 104051
rect 30437 103989 30747 104023
rect 30437 103961 30485 103989
rect 30513 103961 30547 103989
rect 30575 103961 30609 103989
rect 30637 103961 30671 103989
rect 30699 103961 30747 103989
rect 30437 95175 30747 103961
rect 30437 95147 30485 95175
rect 30513 95147 30547 95175
rect 30575 95147 30609 95175
rect 30637 95147 30671 95175
rect 30699 95147 30747 95175
rect 30437 95113 30747 95147
rect 30437 95085 30485 95113
rect 30513 95085 30547 95113
rect 30575 95085 30609 95113
rect 30637 95085 30671 95113
rect 30699 95085 30747 95113
rect 30437 95051 30747 95085
rect 30437 95023 30485 95051
rect 30513 95023 30547 95051
rect 30575 95023 30609 95051
rect 30637 95023 30671 95051
rect 30699 95023 30747 95051
rect 30437 94989 30747 95023
rect 30437 94961 30485 94989
rect 30513 94961 30547 94989
rect 30575 94961 30609 94989
rect 30637 94961 30671 94989
rect 30699 94961 30747 94989
rect 30437 86175 30747 94961
rect 30437 86147 30485 86175
rect 30513 86147 30547 86175
rect 30575 86147 30609 86175
rect 30637 86147 30671 86175
rect 30699 86147 30747 86175
rect 30437 86113 30747 86147
rect 30437 86085 30485 86113
rect 30513 86085 30547 86113
rect 30575 86085 30609 86113
rect 30637 86085 30671 86113
rect 30699 86085 30747 86113
rect 30437 86051 30747 86085
rect 30437 86023 30485 86051
rect 30513 86023 30547 86051
rect 30575 86023 30609 86051
rect 30637 86023 30671 86051
rect 30699 86023 30747 86051
rect 30437 85989 30747 86023
rect 30437 85961 30485 85989
rect 30513 85961 30547 85989
rect 30575 85961 30609 85989
rect 30637 85961 30671 85989
rect 30699 85961 30747 85989
rect 30437 77175 30747 85961
rect 30437 77147 30485 77175
rect 30513 77147 30547 77175
rect 30575 77147 30609 77175
rect 30637 77147 30671 77175
rect 30699 77147 30747 77175
rect 30437 77113 30747 77147
rect 30437 77085 30485 77113
rect 30513 77085 30547 77113
rect 30575 77085 30609 77113
rect 30637 77085 30671 77113
rect 30699 77085 30747 77113
rect 30437 77051 30747 77085
rect 30437 77023 30485 77051
rect 30513 77023 30547 77051
rect 30575 77023 30609 77051
rect 30637 77023 30671 77051
rect 30699 77023 30747 77051
rect 30437 76989 30747 77023
rect 30437 76961 30485 76989
rect 30513 76961 30547 76989
rect 30575 76961 30609 76989
rect 30637 76961 30671 76989
rect 30699 76961 30747 76989
rect 30437 68175 30747 76961
rect 30437 68147 30485 68175
rect 30513 68147 30547 68175
rect 30575 68147 30609 68175
rect 30637 68147 30671 68175
rect 30699 68147 30747 68175
rect 30437 68113 30747 68147
rect 30437 68085 30485 68113
rect 30513 68085 30547 68113
rect 30575 68085 30609 68113
rect 30637 68085 30671 68113
rect 30699 68085 30747 68113
rect 30437 68051 30747 68085
rect 30437 68023 30485 68051
rect 30513 68023 30547 68051
rect 30575 68023 30609 68051
rect 30637 68023 30671 68051
rect 30699 68023 30747 68051
rect 30437 67989 30747 68023
rect 30437 67961 30485 67989
rect 30513 67961 30547 67989
rect 30575 67961 30609 67989
rect 30637 67961 30671 67989
rect 30699 67961 30747 67989
rect 30437 59175 30747 67961
rect 30437 59147 30485 59175
rect 30513 59147 30547 59175
rect 30575 59147 30609 59175
rect 30637 59147 30671 59175
rect 30699 59147 30747 59175
rect 30437 59113 30747 59147
rect 30437 59085 30485 59113
rect 30513 59085 30547 59113
rect 30575 59085 30609 59113
rect 30637 59085 30671 59113
rect 30699 59085 30747 59113
rect 30437 59051 30747 59085
rect 30437 59023 30485 59051
rect 30513 59023 30547 59051
rect 30575 59023 30609 59051
rect 30637 59023 30671 59051
rect 30699 59023 30747 59051
rect 30437 58989 30747 59023
rect 30437 58961 30485 58989
rect 30513 58961 30547 58989
rect 30575 58961 30609 58989
rect 30637 58961 30671 58989
rect 30699 58961 30747 58989
rect 30437 50175 30747 58961
rect 30437 50147 30485 50175
rect 30513 50147 30547 50175
rect 30575 50147 30609 50175
rect 30637 50147 30671 50175
rect 30699 50147 30747 50175
rect 30437 50113 30747 50147
rect 30437 50085 30485 50113
rect 30513 50085 30547 50113
rect 30575 50085 30609 50113
rect 30637 50085 30671 50113
rect 30699 50085 30747 50113
rect 30437 50051 30747 50085
rect 30437 50023 30485 50051
rect 30513 50023 30547 50051
rect 30575 50023 30609 50051
rect 30637 50023 30671 50051
rect 30699 50023 30747 50051
rect 30437 49989 30747 50023
rect 30437 49961 30485 49989
rect 30513 49961 30547 49989
rect 30575 49961 30609 49989
rect 30637 49961 30671 49989
rect 30699 49961 30747 49989
rect 30437 41175 30747 49961
rect 30437 41147 30485 41175
rect 30513 41147 30547 41175
rect 30575 41147 30609 41175
rect 30637 41147 30671 41175
rect 30699 41147 30747 41175
rect 30437 41113 30747 41147
rect 30437 41085 30485 41113
rect 30513 41085 30547 41113
rect 30575 41085 30609 41113
rect 30637 41085 30671 41113
rect 30699 41085 30747 41113
rect 30437 41051 30747 41085
rect 30437 41023 30485 41051
rect 30513 41023 30547 41051
rect 30575 41023 30609 41051
rect 30637 41023 30671 41051
rect 30699 41023 30747 41051
rect 30437 40989 30747 41023
rect 30437 40961 30485 40989
rect 30513 40961 30547 40989
rect 30575 40961 30609 40989
rect 30637 40961 30671 40989
rect 30699 40961 30747 40989
rect 30437 32175 30747 40961
rect 30437 32147 30485 32175
rect 30513 32147 30547 32175
rect 30575 32147 30609 32175
rect 30637 32147 30671 32175
rect 30699 32147 30747 32175
rect 30437 32113 30747 32147
rect 30437 32085 30485 32113
rect 30513 32085 30547 32113
rect 30575 32085 30609 32113
rect 30637 32085 30671 32113
rect 30699 32085 30747 32113
rect 30437 32051 30747 32085
rect 30437 32023 30485 32051
rect 30513 32023 30547 32051
rect 30575 32023 30609 32051
rect 30637 32023 30671 32051
rect 30699 32023 30747 32051
rect 30437 31989 30747 32023
rect 30437 31961 30485 31989
rect 30513 31961 30547 31989
rect 30575 31961 30609 31989
rect 30637 31961 30671 31989
rect 30699 31961 30747 31989
rect 30437 23175 30747 31961
rect 30437 23147 30485 23175
rect 30513 23147 30547 23175
rect 30575 23147 30609 23175
rect 30637 23147 30671 23175
rect 30699 23147 30747 23175
rect 30437 23113 30747 23147
rect 30437 23085 30485 23113
rect 30513 23085 30547 23113
rect 30575 23085 30609 23113
rect 30637 23085 30671 23113
rect 30699 23085 30747 23113
rect 30437 23051 30747 23085
rect 30437 23023 30485 23051
rect 30513 23023 30547 23051
rect 30575 23023 30609 23051
rect 30637 23023 30671 23051
rect 30699 23023 30747 23051
rect 30437 22989 30747 23023
rect 30437 22961 30485 22989
rect 30513 22961 30547 22989
rect 30575 22961 30609 22989
rect 30637 22961 30671 22989
rect 30699 22961 30747 22989
rect 30437 14175 30747 22961
rect 30437 14147 30485 14175
rect 30513 14147 30547 14175
rect 30575 14147 30609 14175
rect 30637 14147 30671 14175
rect 30699 14147 30747 14175
rect 30437 14113 30747 14147
rect 30437 14085 30485 14113
rect 30513 14085 30547 14113
rect 30575 14085 30609 14113
rect 30637 14085 30671 14113
rect 30699 14085 30747 14113
rect 30437 14051 30747 14085
rect 30437 14023 30485 14051
rect 30513 14023 30547 14051
rect 30575 14023 30609 14051
rect 30637 14023 30671 14051
rect 30699 14023 30747 14051
rect 30437 13989 30747 14023
rect 30437 13961 30485 13989
rect 30513 13961 30547 13989
rect 30575 13961 30609 13989
rect 30637 13961 30671 13989
rect 30699 13961 30747 13989
rect 30437 5175 30747 13961
rect 30437 5147 30485 5175
rect 30513 5147 30547 5175
rect 30575 5147 30609 5175
rect 30637 5147 30671 5175
rect 30699 5147 30747 5175
rect 30437 5113 30747 5147
rect 30437 5085 30485 5113
rect 30513 5085 30547 5113
rect 30575 5085 30609 5113
rect 30637 5085 30671 5113
rect 30699 5085 30747 5113
rect 30437 5051 30747 5085
rect 30437 5023 30485 5051
rect 30513 5023 30547 5051
rect 30575 5023 30609 5051
rect 30637 5023 30671 5051
rect 30699 5023 30747 5051
rect 30437 4989 30747 5023
rect 30437 4961 30485 4989
rect 30513 4961 30547 4989
rect 30575 4961 30609 4989
rect 30637 4961 30671 4989
rect 30699 4961 30747 4989
rect 30437 -560 30747 4961
rect 30437 -588 30485 -560
rect 30513 -588 30547 -560
rect 30575 -588 30609 -560
rect 30637 -588 30671 -560
rect 30699 -588 30747 -560
rect 30437 -622 30747 -588
rect 30437 -650 30485 -622
rect 30513 -650 30547 -622
rect 30575 -650 30609 -622
rect 30637 -650 30671 -622
rect 30699 -650 30747 -622
rect 30437 -684 30747 -650
rect 30437 -712 30485 -684
rect 30513 -712 30547 -684
rect 30575 -712 30609 -684
rect 30637 -712 30671 -684
rect 30699 -712 30747 -684
rect 30437 -746 30747 -712
rect 30437 -774 30485 -746
rect 30513 -774 30547 -746
rect 30575 -774 30609 -746
rect 30637 -774 30671 -746
rect 30699 -774 30747 -746
rect 30437 -822 30747 -774
rect 37577 298606 37887 299134
rect 37577 298578 37625 298606
rect 37653 298578 37687 298606
rect 37715 298578 37749 298606
rect 37777 298578 37811 298606
rect 37839 298578 37887 298606
rect 37577 298544 37887 298578
rect 37577 298516 37625 298544
rect 37653 298516 37687 298544
rect 37715 298516 37749 298544
rect 37777 298516 37811 298544
rect 37839 298516 37887 298544
rect 37577 298482 37887 298516
rect 37577 298454 37625 298482
rect 37653 298454 37687 298482
rect 37715 298454 37749 298482
rect 37777 298454 37811 298482
rect 37839 298454 37887 298482
rect 37577 298420 37887 298454
rect 37577 298392 37625 298420
rect 37653 298392 37687 298420
rect 37715 298392 37749 298420
rect 37777 298392 37811 298420
rect 37839 298392 37887 298420
rect 37577 290175 37887 298392
rect 37577 290147 37625 290175
rect 37653 290147 37687 290175
rect 37715 290147 37749 290175
rect 37777 290147 37811 290175
rect 37839 290147 37887 290175
rect 37577 290113 37887 290147
rect 37577 290085 37625 290113
rect 37653 290085 37687 290113
rect 37715 290085 37749 290113
rect 37777 290085 37811 290113
rect 37839 290085 37887 290113
rect 37577 290051 37887 290085
rect 37577 290023 37625 290051
rect 37653 290023 37687 290051
rect 37715 290023 37749 290051
rect 37777 290023 37811 290051
rect 37839 290023 37887 290051
rect 37577 289989 37887 290023
rect 37577 289961 37625 289989
rect 37653 289961 37687 289989
rect 37715 289961 37749 289989
rect 37777 289961 37811 289989
rect 37839 289961 37887 289989
rect 37577 281175 37887 289961
rect 37577 281147 37625 281175
rect 37653 281147 37687 281175
rect 37715 281147 37749 281175
rect 37777 281147 37811 281175
rect 37839 281147 37887 281175
rect 37577 281113 37887 281147
rect 37577 281085 37625 281113
rect 37653 281085 37687 281113
rect 37715 281085 37749 281113
rect 37777 281085 37811 281113
rect 37839 281085 37887 281113
rect 37577 281051 37887 281085
rect 37577 281023 37625 281051
rect 37653 281023 37687 281051
rect 37715 281023 37749 281051
rect 37777 281023 37811 281051
rect 37839 281023 37887 281051
rect 37577 280989 37887 281023
rect 37577 280961 37625 280989
rect 37653 280961 37687 280989
rect 37715 280961 37749 280989
rect 37777 280961 37811 280989
rect 37839 280961 37887 280989
rect 37577 272175 37887 280961
rect 37577 272147 37625 272175
rect 37653 272147 37687 272175
rect 37715 272147 37749 272175
rect 37777 272147 37811 272175
rect 37839 272147 37887 272175
rect 37577 272113 37887 272147
rect 37577 272085 37625 272113
rect 37653 272085 37687 272113
rect 37715 272085 37749 272113
rect 37777 272085 37811 272113
rect 37839 272085 37887 272113
rect 37577 272051 37887 272085
rect 37577 272023 37625 272051
rect 37653 272023 37687 272051
rect 37715 272023 37749 272051
rect 37777 272023 37811 272051
rect 37839 272023 37887 272051
rect 37577 271989 37887 272023
rect 37577 271961 37625 271989
rect 37653 271961 37687 271989
rect 37715 271961 37749 271989
rect 37777 271961 37811 271989
rect 37839 271961 37887 271989
rect 37577 263175 37887 271961
rect 37577 263147 37625 263175
rect 37653 263147 37687 263175
rect 37715 263147 37749 263175
rect 37777 263147 37811 263175
rect 37839 263147 37887 263175
rect 37577 263113 37887 263147
rect 37577 263085 37625 263113
rect 37653 263085 37687 263113
rect 37715 263085 37749 263113
rect 37777 263085 37811 263113
rect 37839 263085 37887 263113
rect 37577 263051 37887 263085
rect 37577 263023 37625 263051
rect 37653 263023 37687 263051
rect 37715 263023 37749 263051
rect 37777 263023 37811 263051
rect 37839 263023 37887 263051
rect 37577 262989 37887 263023
rect 37577 262961 37625 262989
rect 37653 262961 37687 262989
rect 37715 262961 37749 262989
rect 37777 262961 37811 262989
rect 37839 262961 37887 262989
rect 37577 254175 37887 262961
rect 37577 254147 37625 254175
rect 37653 254147 37687 254175
rect 37715 254147 37749 254175
rect 37777 254147 37811 254175
rect 37839 254147 37887 254175
rect 37577 254113 37887 254147
rect 37577 254085 37625 254113
rect 37653 254085 37687 254113
rect 37715 254085 37749 254113
rect 37777 254085 37811 254113
rect 37839 254085 37887 254113
rect 37577 254051 37887 254085
rect 37577 254023 37625 254051
rect 37653 254023 37687 254051
rect 37715 254023 37749 254051
rect 37777 254023 37811 254051
rect 37839 254023 37887 254051
rect 37577 253989 37887 254023
rect 37577 253961 37625 253989
rect 37653 253961 37687 253989
rect 37715 253961 37749 253989
rect 37777 253961 37811 253989
rect 37839 253961 37887 253989
rect 37577 245175 37887 253961
rect 37577 245147 37625 245175
rect 37653 245147 37687 245175
rect 37715 245147 37749 245175
rect 37777 245147 37811 245175
rect 37839 245147 37887 245175
rect 37577 245113 37887 245147
rect 37577 245085 37625 245113
rect 37653 245085 37687 245113
rect 37715 245085 37749 245113
rect 37777 245085 37811 245113
rect 37839 245085 37887 245113
rect 37577 245051 37887 245085
rect 37577 245023 37625 245051
rect 37653 245023 37687 245051
rect 37715 245023 37749 245051
rect 37777 245023 37811 245051
rect 37839 245023 37887 245051
rect 37577 244989 37887 245023
rect 37577 244961 37625 244989
rect 37653 244961 37687 244989
rect 37715 244961 37749 244989
rect 37777 244961 37811 244989
rect 37839 244961 37887 244989
rect 37577 236175 37887 244961
rect 37577 236147 37625 236175
rect 37653 236147 37687 236175
rect 37715 236147 37749 236175
rect 37777 236147 37811 236175
rect 37839 236147 37887 236175
rect 37577 236113 37887 236147
rect 37577 236085 37625 236113
rect 37653 236085 37687 236113
rect 37715 236085 37749 236113
rect 37777 236085 37811 236113
rect 37839 236085 37887 236113
rect 37577 236051 37887 236085
rect 37577 236023 37625 236051
rect 37653 236023 37687 236051
rect 37715 236023 37749 236051
rect 37777 236023 37811 236051
rect 37839 236023 37887 236051
rect 37577 235989 37887 236023
rect 37577 235961 37625 235989
rect 37653 235961 37687 235989
rect 37715 235961 37749 235989
rect 37777 235961 37811 235989
rect 37839 235961 37887 235989
rect 37577 227175 37887 235961
rect 37577 227147 37625 227175
rect 37653 227147 37687 227175
rect 37715 227147 37749 227175
rect 37777 227147 37811 227175
rect 37839 227147 37887 227175
rect 37577 227113 37887 227147
rect 37577 227085 37625 227113
rect 37653 227085 37687 227113
rect 37715 227085 37749 227113
rect 37777 227085 37811 227113
rect 37839 227085 37887 227113
rect 37577 227051 37887 227085
rect 37577 227023 37625 227051
rect 37653 227023 37687 227051
rect 37715 227023 37749 227051
rect 37777 227023 37811 227051
rect 37839 227023 37887 227051
rect 37577 226989 37887 227023
rect 37577 226961 37625 226989
rect 37653 226961 37687 226989
rect 37715 226961 37749 226989
rect 37777 226961 37811 226989
rect 37839 226961 37887 226989
rect 37577 218175 37887 226961
rect 37577 218147 37625 218175
rect 37653 218147 37687 218175
rect 37715 218147 37749 218175
rect 37777 218147 37811 218175
rect 37839 218147 37887 218175
rect 37577 218113 37887 218147
rect 37577 218085 37625 218113
rect 37653 218085 37687 218113
rect 37715 218085 37749 218113
rect 37777 218085 37811 218113
rect 37839 218085 37887 218113
rect 37577 218051 37887 218085
rect 37577 218023 37625 218051
rect 37653 218023 37687 218051
rect 37715 218023 37749 218051
rect 37777 218023 37811 218051
rect 37839 218023 37887 218051
rect 37577 217989 37887 218023
rect 37577 217961 37625 217989
rect 37653 217961 37687 217989
rect 37715 217961 37749 217989
rect 37777 217961 37811 217989
rect 37839 217961 37887 217989
rect 37577 209175 37887 217961
rect 37577 209147 37625 209175
rect 37653 209147 37687 209175
rect 37715 209147 37749 209175
rect 37777 209147 37811 209175
rect 37839 209147 37887 209175
rect 37577 209113 37887 209147
rect 37577 209085 37625 209113
rect 37653 209085 37687 209113
rect 37715 209085 37749 209113
rect 37777 209085 37811 209113
rect 37839 209085 37887 209113
rect 37577 209051 37887 209085
rect 37577 209023 37625 209051
rect 37653 209023 37687 209051
rect 37715 209023 37749 209051
rect 37777 209023 37811 209051
rect 37839 209023 37887 209051
rect 37577 208989 37887 209023
rect 37577 208961 37625 208989
rect 37653 208961 37687 208989
rect 37715 208961 37749 208989
rect 37777 208961 37811 208989
rect 37839 208961 37887 208989
rect 37577 200175 37887 208961
rect 37577 200147 37625 200175
rect 37653 200147 37687 200175
rect 37715 200147 37749 200175
rect 37777 200147 37811 200175
rect 37839 200147 37887 200175
rect 37577 200113 37887 200147
rect 37577 200085 37625 200113
rect 37653 200085 37687 200113
rect 37715 200085 37749 200113
rect 37777 200085 37811 200113
rect 37839 200085 37887 200113
rect 37577 200051 37887 200085
rect 37577 200023 37625 200051
rect 37653 200023 37687 200051
rect 37715 200023 37749 200051
rect 37777 200023 37811 200051
rect 37839 200023 37887 200051
rect 37577 199989 37887 200023
rect 37577 199961 37625 199989
rect 37653 199961 37687 199989
rect 37715 199961 37749 199989
rect 37777 199961 37811 199989
rect 37839 199961 37887 199989
rect 37577 191175 37887 199961
rect 37577 191147 37625 191175
rect 37653 191147 37687 191175
rect 37715 191147 37749 191175
rect 37777 191147 37811 191175
rect 37839 191147 37887 191175
rect 37577 191113 37887 191147
rect 37577 191085 37625 191113
rect 37653 191085 37687 191113
rect 37715 191085 37749 191113
rect 37777 191085 37811 191113
rect 37839 191085 37887 191113
rect 37577 191051 37887 191085
rect 37577 191023 37625 191051
rect 37653 191023 37687 191051
rect 37715 191023 37749 191051
rect 37777 191023 37811 191051
rect 37839 191023 37887 191051
rect 37577 190989 37887 191023
rect 37577 190961 37625 190989
rect 37653 190961 37687 190989
rect 37715 190961 37749 190989
rect 37777 190961 37811 190989
rect 37839 190961 37887 190989
rect 37577 182175 37887 190961
rect 37577 182147 37625 182175
rect 37653 182147 37687 182175
rect 37715 182147 37749 182175
rect 37777 182147 37811 182175
rect 37839 182147 37887 182175
rect 37577 182113 37887 182147
rect 37577 182085 37625 182113
rect 37653 182085 37687 182113
rect 37715 182085 37749 182113
rect 37777 182085 37811 182113
rect 37839 182085 37887 182113
rect 37577 182051 37887 182085
rect 37577 182023 37625 182051
rect 37653 182023 37687 182051
rect 37715 182023 37749 182051
rect 37777 182023 37811 182051
rect 37839 182023 37887 182051
rect 37577 181989 37887 182023
rect 37577 181961 37625 181989
rect 37653 181961 37687 181989
rect 37715 181961 37749 181989
rect 37777 181961 37811 181989
rect 37839 181961 37887 181989
rect 37577 173175 37887 181961
rect 37577 173147 37625 173175
rect 37653 173147 37687 173175
rect 37715 173147 37749 173175
rect 37777 173147 37811 173175
rect 37839 173147 37887 173175
rect 37577 173113 37887 173147
rect 37577 173085 37625 173113
rect 37653 173085 37687 173113
rect 37715 173085 37749 173113
rect 37777 173085 37811 173113
rect 37839 173085 37887 173113
rect 37577 173051 37887 173085
rect 37577 173023 37625 173051
rect 37653 173023 37687 173051
rect 37715 173023 37749 173051
rect 37777 173023 37811 173051
rect 37839 173023 37887 173051
rect 37577 172989 37887 173023
rect 37577 172961 37625 172989
rect 37653 172961 37687 172989
rect 37715 172961 37749 172989
rect 37777 172961 37811 172989
rect 37839 172961 37887 172989
rect 37577 164175 37887 172961
rect 37577 164147 37625 164175
rect 37653 164147 37687 164175
rect 37715 164147 37749 164175
rect 37777 164147 37811 164175
rect 37839 164147 37887 164175
rect 37577 164113 37887 164147
rect 37577 164085 37625 164113
rect 37653 164085 37687 164113
rect 37715 164085 37749 164113
rect 37777 164085 37811 164113
rect 37839 164085 37887 164113
rect 37577 164051 37887 164085
rect 37577 164023 37625 164051
rect 37653 164023 37687 164051
rect 37715 164023 37749 164051
rect 37777 164023 37811 164051
rect 37839 164023 37887 164051
rect 37577 163989 37887 164023
rect 37577 163961 37625 163989
rect 37653 163961 37687 163989
rect 37715 163961 37749 163989
rect 37777 163961 37811 163989
rect 37839 163961 37887 163989
rect 37577 155175 37887 163961
rect 37577 155147 37625 155175
rect 37653 155147 37687 155175
rect 37715 155147 37749 155175
rect 37777 155147 37811 155175
rect 37839 155147 37887 155175
rect 37577 155113 37887 155147
rect 37577 155085 37625 155113
rect 37653 155085 37687 155113
rect 37715 155085 37749 155113
rect 37777 155085 37811 155113
rect 37839 155085 37887 155113
rect 37577 155051 37887 155085
rect 37577 155023 37625 155051
rect 37653 155023 37687 155051
rect 37715 155023 37749 155051
rect 37777 155023 37811 155051
rect 37839 155023 37887 155051
rect 37577 154989 37887 155023
rect 37577 154961 37625 154989
rect 37653 154961 37687 154989
rect 37715 154961 37749 154989
rect 37777 154961 37811 154989
rect 37839 154961 37887 154989
rect 37577 146175 37887 154961
rect 37577 146147 37625 146175
rect 37653 146147 37687 146175
rect 37715 146147 37749 146175
rect 37777 146147 37811 146175
rect 37839 146147 37887 146175
rect 37577 146113 37887 146147
rect 37577 146085 37625 146113
rect 37653 146085 37687 146113
rect 37715 146085 37749 146113
rect 37777 146085 37811 146113
rect 37839 146085 37887 146113
rect 37577 146051 37887 146085
rect 37577 146023 37625 146051
rect 37653 146023 37687 146051
rect 37715 146023 37749 146051
rect 37777 146023 37811 146051
rect 37839 146023 37887 146051
rect 37577 145989 37887 146023
rect 37577 145961 37625 145989
rect 37653 145961 37687 145989
rect 37715 145961 37749 145989
rect 37777 145961 37811 145989
rect 37839 145961 37887 145989
rect 37577 137175 37887 145961
rect 37577 137147 37625 137175
rect 37653 137147 37687 137175
rect 37715 137147 37749 137175
rect 37777 137147 37811 137175
rect 37839 137147 37887 137175
rect 37577 137113 37887 137147
rect 37577 137085 37625 137113
rect 37653 137085 37687 137113
rect 37715 137085 37749 137113
rect 37777 137085 37811 137113
rect 37839 137085 37887 137113
rect 37577 137051 37887 137085
rect 37577 137023 37625 137051
rect 37653 137023 37687 137051
rect 37715 137023 37749 137051
rect 37777 137023 37811 137051
rect 37839 137023 37887 137051
rect 37577 136989 37887 137023
rect 37577 136961 37625 136989
rect 37653 136961 37687 136989
rect 37715 136961 37749 136989
rect 37777 136961 37811 136989
rect 37839 136961 37887 136989
rect 37577 128175 37887 136961
rect 37577 128147 37625 128175
rect 37653 128147 37687 128175
rect 37715 128147 37749 128175
rect 37777 128147 37811 128175
rect 37839 128147 37887 128175
rect 37577 128113 37887 128147
rect 37577 128085 37625 128113
rect 37653 128085 37687 128113
rect 37715 128085 37749 128113
rect 37777 128085 37811 128113
rect 37839 128085 37887 128113
rect 37577 128051 37887 128085
rect 37577 128023 37625 128051
rect 37653 128023 37687 128051
rect 37715 128023 37749 128051
rect 37777 128023 37811 128051
rect 37839 128023 37887 128051
rect 37577 127989 37887 128023
rect 37577 127961 37625 127989
rect 37653 127961 37687 127989
rect 37715 127961 37749 127989
rect 37777 127961 37811 127989
rect 37839 127961 37887 127989
rect 37577 119175 37887 127961
rect 37577 119147 37625 119175
rect 37653 119147 37687 119175
rect 37715 119147 37749 119175
rect 37777 119147 37811 119175
rect 37839 119147 37887 119175
rect 37577 119113 37887 119147
rect 37577 119085 37625 119113
rect 37653 119085 37687 119113
rect 37715 119085 37749 119113
rect 37777 119085 37811 119113
rect 37839 119085 37887 119113
rect 37577 119051 37887 119085
rect 37577 119023 37625 119051
rect 37653 119023 37687 119051
rect 37715 119023 37749 119051
rect 37777 119023 37811 119051
rect 37839 119023 37887 119051
rect 37577 118989 37887 119023
rect 37577 118961 37625 118989
rect 37653 118961 37687 118989
rect 37715 118961 37749 118989
rect 37777 118961 37811 118989
rect 37839 118961 37887 118989
rect 37577 110175 37887 118961
rect 37577 110147 37625 110175
rect 37653 110147 37687 110175
rect 37715 110147 37749 110175
rect 37777 110147 37811 110175
rect 37839 110147 37887 110175
rect 37577 110113 37887 110147
rect 37577 110085 37625 110113
rect 37653 110085 37687 110113
rect 37715 110085 37749 110113
rect 37777 110085 37811 110113
rect 37839 110085 37887 110113
rect 37577 110051 37887 110085
rect 37577 110023 37625 110051
rect 37653 110023 37687 110051
rect 37715 110023 37749 110051
rect 37777 110023 37811 110051
rect 37839 110023 37887 110051
rect 37577 109989 37887 110023
rect 37577 109961 37625 109989
rect 37653 109961 37687 109989
rect 37715 109961 37749 109989
rect 37777 109961 37811 109989
rect 37839 109961 37887 109989
rect 37577 101175 37887 109961
rect 37577 101147 37625 101175
rect 37653 101147 37687 101175
rect 37715 101147 37749 101175
rect 37777 101147 37811 101175
rect 37839 101147 37887 101175
rect 37577 101113 37887 101147
rect 37577 101085 37625 101113
rect 37653 101085 37687 101113
rect 37715 101085 37749 101113
rect 37777 101085 37811 101113
rect 37839 101085 37887 101113
rect 37577 101051 37887 101085
rect 37577 101023 37625 101051
rect 37653 101023 37687 101051
rect 37715 101023 37749 101051
rect 37777 101023 37811 101051
rect 37839 101023 37887 101051
rect 37577 100989 37887 101023
rect 37577 100961 37625 100989
rect 37653 100961 37687 100989
rect 37715 100961 37749 100989
rect 37777 100961 37811 100989
rect 37839 100961 37887 100989
rect 37577 92175 37887 100961
rect 37577 92147 37625 92175
rect 37653 92147 37687 92175
rect 37715 92147 37749 92175
rect 37777 92147 37811 92175
rect 37839 92147 37887 92175
rect 37577 92113 37887 92147
rect 37577 92085 37625 92113
rect 37653 92085 37687 92113
rect 37715 92085 37749 92113
rect 37777 92085 37811 92113
rect 37839 92085 37887 92113
rect 37577 92051 37887 92085
rect 37577 92023 37625 92051
rect 37653 92023 37687 92051
rect 37715 92023 37749 92051
rect 37777 92023 37811 92051
rect 37839 92023 37887 92051
rect 37577 91989 37887 92023
rect 37577 91961 37625 91989
rect 37653 91961 37687 91989
rect 37715 91961 37749 91989
rect 37777 91961 37811 91989
rect 37839 91961 37887 91989
rect 37577 83175 37887 91961
rect 37577 83147 37625 83175
rect 37653 83147 37687 83175
rect 37715 83147 37749 83175
rect 37777 83147 37811 83175
rect 37839 83147 37887 83175
rect 37577 83113 37887 83147
rect 37577 83085 37625 83113
rect 37653 83085 37687 83113
rect 37715 83085 37749 83113
rect 37777 83085 37811 83113
rect 37839 83085 37887 83113
rect 37577 83051 37887 83085
rect 37577 83023 37625 83051
rect 37653 83023 37687 83051
rect 37715 83023 37749 83051
rect 37777 83023 37811 83051
rect 37839 83023 37887 83051
rect 37577 82989 37887 83023
rect 37577 82961 37625 82989
rect 37653 82961 37687 82989
rect 37715 82961 37749 82989
rect 37777 82961 37811 82989
rect 37839 82961 37887 82989
rect 37577 74175 37887 82961
rect 37577 74147 37625 74175
rect 37653 74147 37687 74175
rect 37715 74147 37749 74175
rect 37777 74147 37811 74175
rect 37839 74147 37887 74175
rect 37577 74113 37887 74147
rect 37577 74085 37625 74113
rect 37653 74085 37687 74113
rect 37715 74085 37749 74113
rect 37777 74085 37811 74113
rect 37839 74085 37887 74113
rect 37577 74051 37887 74085
rect 37577 74023 37625 74051
rect 37653 74023 37687 74051
rect 37715 74023 37749 74051
rect 37777 74023 37811 74051
rect 37839 74023 37887 74051
rect 37577 73989 37887 74023
rect 37577 73961 37625 73989
rect 37653 73961 37687 73989
rect 37715 73961 37749 73989
rect 37777 73961 37811 73989
rect 37839 73961 37887 73989
rect 37577 65175 37887 73961
rect 37577 65147 37625 65175
rect 37653 65147 37687 65175
rect 37715 65147 37749 65175
rect 37777 65147 37811 65175
rect 37839 65147 37887 65175
rect 37577 65113 37887 65147
rect 37577 65085 37625 65113
rect 37653 65085 37687 65113
rect 37715 65085 37749 65113
rect 37777 65085 37811 65113
rect 37839 65085 37887 65113
rect 37577 65051 37887 65085
rect 37577 65023 37625 65051
rect 37653 65023 37687 65051
rect 37715 65023 37749 65051
rect 37777 65023 37811 65051
rect 37839 65023 37887 65051
rect 37577 64989 37887 65023
rect 37577 64961 37625 64989
rect 37653 64961 37687 64989
rect 37715 64961 37749 64989
rect 37777 64961 37811 64989
rect 37839 64961 37887 64989
rect 37577 56175 37887 64961
rect 37577 56147 37625 56175
rect 37653 56147 37687 56175
rect 37715 56147 37749 56175
rect 37777 56147 37811 56175
rect 37839 56147 37887 56175
rect 37577 56113 37887 56147
rect 37577 56085 37625 56113
rect 37653 56085 37687 56113
rect 37715 56085 37749 56113
rect 37777 56085 37811 56113
rect 37839 56085 37887 56113
rect 37577 56051 37887 56085
rect 37577 56023 37625 56051
rect 37653 56023 37687 56051
rect 37715 56023 37749 56051
rect 37777 56023 37811 56051
rect 37839 56023 37887 56051
rect 37577 55989 37887 56023
rect 37577 55961 37625 55989
rect 37653 55961 37687 55989
rect 37715 55961 37749 55989
rect 37777 55961 37811 55989
rect 37839 55961 37887 55989
rect 37577 47175 37887 55961
rect 37577 47147 37625 47175
rect 37653 47147 37687 47175
rect 37715 47147 37749 47175
rect 37777 47147 37811 47175
rect 37839 47147 37887 47175
rect 37577 47113 37887 47147
rect 37577 47085 37625 47113
rect 37653 47085 37687 47113
rect 37715 47085 37749 47113
rect 37777 47085 37811 47113
rect 37839 47085 37887 47113
rect 37577 47051 37887 47085
rect 37577 47023 37625 47051
rect 37653 47023 37687 47051
rect 37715 47023 37749 47051
rect 37777 47023 37811 47051
rect 37839 47023 37887 47051
rect 37577 46989 37887 47023
rect 37577 46961 37625 46989
rect 37653 46961 37687 46989
rect 37715 46961 37749 46989
rect 37777 46961 37811 46989
rect 37839 46961 37887 46989
rect 37577 38175 37887 46961
rect 37577 38147 37625 38175
rect 37653 38147 37687 38175
rect 37715 38147 37749 38175
rect 37777 38147 37811 38175
rect 37839 38147 37887 38175
rect 37577 38113 37887 38147
rect 37577 38085 37625 38113
rect 37653 38085 37687 38113
rect 37715 38085 37749 38113
rect 37777 38085 37811 38113
rect 37839 38085 37887 38113
rect 37577 38051 37887 38085
rect 37577 38023 37625 38051
rect 37653 38023 37687 38051
rect 37715 38023 37749 38051
rect 37777 38023 37811 38051
rect 37839 38023 37887 38051
rect 37577 37989 37887 38023
rect 37577 37961 37625 37989
rect 37653 37961 37687 37989
rect 37715 37961 37749 37989
rect 37777 37961 37811 37989
rect 37839 37961 37887 37989
rect 37577 29175 37887 37961
rect 37577 29147 37625 29175
rect 37653 29147 37687 29175
rect 37715 29147 37749 29175
rect 37777 29147 37811 29175
rect 37839 29147 37887 29175
rect 37577 29113 37887 29147
rect 37577 29085 37625 29113
rect 37653 29085 37687 29113
rect 37715 29085 37749 29113
rect 37777 29085 37811 29113
rect 37839 29085 37887 29113
rect 37577 29051 37887 29085
rect 37577 29023 37625 29051
rect 37653 29023 37687 29051
rect 37715 29023 37749 29051
rect 37777 29023 37811 29051
rect 37839 29023 37887 29051
rect 37577 28989 37887 29023
rect 37577 28961 37625 28989
rect 37653 28961 37687 28989
rect 37715 28961 37749 28989
rect 37777 28961 37811 28989
rect 37839 28961 37887 28989
rect 37577 20175 37887 28961
rect 37577 20147 37625 20175
rect 37653 20147 37687 20175
rect 37715 20147 37749 20175
rect 37777 20147 37811 20175
rect 37839 20147 37887 20175
rect 37577 20113 37887 20147
rect 37577 20085 37625 20113
rect 37653 20085 37687 20113
rect 37715 20085 37749 20113
rect 37777 20085 37811 20113
rect 37839 20085 37887 20113
rect 37577 20051 37887 20085
rect 37577 20023 37625 20051
rect 37653 20023 37687 20051
rect 37715 20023 37749 20051
rect 37777 20023 37811 20051
rect 37839 20023 37887 20051
rect 37577 19989 37887 20023
rect 37577 19961 37625 19989
rect 37653 19961 37687 19989
rect 37715 19961 37749 19989
rect 37777 19961 37811 19989
rect 37839 19961 37887 19989
rect 37577 11175 37887 19961
rect 37577 11147 37625 11175
rect 37653 11147 37687 11175
rect 37715 11147 37749 11175
rect 37777 11147 37811 11175
rect 37839 11147 37887 11175
rect 37577 11113 37887 11147
rect 37577 11085 37625 11113
rect 37653 11085 37687 11113
rect 37715 11085 37749 11113
rect 37777 11085 37811 11113
rect 37839 11085 37887 11113
rect 37577 11051 37887 11085
rect 37577 11023 37625 11051
rect 37653 11023 37687 11051
rect 37715 11023 37749 11051
rect 37777 11023 37811 11051
rect 37839 11023 37887 11051
rect 37577 10989 37887 11023
rect 37577 10961 37625 10989
rect 37653 10961 37687 10989
rect 37715 10961 37749 10989
rect 37777 10961 37811 10989
rect 37839 10961 37887 10989
rect 37577 2175 37887 10961
rect 37577 2147 37625 2175
rect 37653 2147 37687 2175
rect 37715 2147 37749 2175
rect 37777 2147 37811 2175
rect 37839 2147 37887 2175
rect 37577 2113 37887 2147
rect 37577 2085 37625 2113
rect 37653 2085 37687 2113
rect 37715 2085 37749 2113
rect 37777 2085 37811 2113
rect 37839 2085 37887 2113
rect 37577 2051 37887 2085
rect 37577 2023 37625 2051
rect 37653 2023 37687 2051
rect 37715 2023 37749 2051
rect 37777 2023 37811 2051
rect 37839 2023 37887 2051
rect 37577 1989 37887 2023
rect 37577 1961 37625 1989
rect 37653 1961 37687 1989
rect 37715 1961 37749 1989
rect 37777 1961 37811 1989
rect 37839 1961 37887 1989
rect 37577 -80 37887 1961
rect 37577 -108 37625 -80
rect 37653 -108 37687 -80
rect 37715 -108 37749 -80
rect 37777 -108 37811 -80
rect 37839 -108 37887 -80
rect 37577 -142 37887 -108
rect 37577 -170 37625 -142
rect 37653 -170 37687 -142
rect 37715 -170 37749 -142
rect 37777 -170 37811 -142
rect 37839 -170 37887 -142
rect 37577 -204 37887 -170
rect 37577 -232 37625 -204
rect 37653 -232 37687 -204
rect 37715 -232 37749 -204
rect 37777 -232 37811 -204
rect 37839 -232 37887 -204
rect 37577 -266 37887 -232
rect 37577 -294 37625 -266
rect 37653 -294 37687 -266
rect 37715 -294 37749 -266
rect 37777 -294 37811 -266
rect 37839 -294 37887 -266
rect 37577 -822 37887 -294
rect 39437 299086 39747 299134
rect 39437 299058 39485 299086
rect 39513 299058 39547 299086
rect 39575 299058 39609 299086
rect 39637 299058 39671 299086
rect 39699 299058 39747 299086
rect 39437 299024 39747 299058
rect 39437 298996 39485 299024
rect 39513 298996 39547 299024
rect 39575 298996 39609 299024
rect 39637 298996 39671 299024
rect 39699 298996 39747 299024
rect 39437 298962 39747 298996
rect 39437 298934 39485 298962
rect 39513 298934 39547 298962
rect 39575 298934 39609 298962
rect 39637 298934 39671 298962
rect 39699 298934 39747 298962
rect 39437 298900 39747 298934
rect 39437 298872 39485 298900
rect 39513 298872 39547 298900
rect 39575 298872 39609 298900
rect 39637 298872 39671 298900
rect 39699 298872 39747 298900
rect 39437 293175 39747 298872
rect 39437 293147 39485 293175
rect 39513 293147 39547 293175
rect 39575 293147 39609 293175
rect 39637 293147 39671 293175
rect 39699 293147 39747 293175
rect 39437 293113 39747 293147
rect 39437 293085 39485 293113
rect 39513 293085 39547 293113
rect 39575 293085 39609 293113
rect 39637 293085 39671 293113
rect 39699 293085 39747 293113
rect 39437 293051 39747 293085
rect 39437 293023 39485 293051
rect 39513 293023 39547 293051
rect 39575 293023 39609 293051
rect 39637 293023 39671 293051
rect 39699 293023 39747 293051
rect 39437 292989 39747 293023
rect 39437 292961 39485 292989
rect 39513 292961 39547 292989
rect 39575 292961 39609 292989
rect 39637 292961 39671 292989
rect 39699 292961 39747 292989
rect 39437 284175 39747 292961
rect 39437 284147 39485 284175
rect 39513 284147 39547 284175
rect 39575 284147 39609 284175
rect 39637 284147 39671 284175
rect 39699 284147 39747 284175
rect 39437 284113 39747 284147
rect 39437 284085 39485 284113
rect 39513 284085 39547 284113
rect 39575 284085 39609 284113
rect 39637 284085 39671 284113
rect 39699 284085 39747 284113
rect 39437 284051 39747 284085
rect 39437 284023 39485 284051
rect 39513 284023 39547 284051
rect 39575 284023 39609 284051
rect 39637 284023 39671 284051
rect 39699 284023 39747 284051
rect 39437 283989 39747 284023
rect 39437 283961 39485 283989
rect 39513 283961 39547 283989
rect 39575 283961 39609 283989
rect 39637 283961 39671 283989
rect 39699 283961 39747 283989
rect 39437 275175 39747 283961
rect 39437 275147 39485 275175
rect 39513 275147 39547 275175
rect 39575 275147 39609 275175
rect 39637 275147 39671 275175
rect 39699 275147 39747 275175
rect 39437 275113 39747 275147
rect 39437 275085 39485 275113
rect 39513 275085 39547 275113
rect 39575 275085 39609 275113
rect 39637 275085 39671 275113
rect 39699 275085 39747 275113
rect 39437 275051 39747 275085
rect 39437 275023 39485 275051
rect 39513 275023 39547 275051
rect 39575 275023 39609 275051
rect 39637 275023 39671 275051
rect 39699 275023 39747 275051
rect 39437 274989 39747 275023
rect 39437 274961 39485 274989
rect 39513 274961 39547 274989
rect 39575 274961 39609 274989
rect 39637 274961 39671 274989
rect 39699 274961 39747 274989
rect 39437 266175 39747 274961
rect 39437 266147 39485 266175
rect 39513 266147 39547 266175
rect 39575 266147 39609 266175
rect 39637 266147 39671 266175
rect 39699 266147 39747 266175
rect 39437 266113 39747 266147
rect 39437 266085 39485 266113
rect 39513 266085 39547 266113
rect 39575 266085 39609 266113
rect 39637 266085 39671 266113
rect 39699 266085 39747 266113
rect 39437 266051 39747 266085
rect 39437 266023 39485 266051
rect 39513 266023 39547 266051
rect 39575 266023 39609 266051
rect 39637 266023 39671 266051
rect 39699 266023 39747 266051
rect 39437 265989 39747 266023
rect 39437 265961 39485 265989
rect 39513 265961 39547 265989
rect 39575 265961 39609 265989
rect 39637 265961 39671 265989
rect 39699 265961 39747 265989
rect 39437 257175 39747 265961
rect 39437 257147 39485 257175
rect 39513 257147 39547 257175
rect 39575 257147 39609 257175
rect 39637 257147 39671 257175
rect 39699 257147 39747 257175
rect 39437 257113 39747 257147
rect 39437 257085 39485 257113
rect 39513 257085 39547 257113
rect 39575 257085 39609 257113
rect 39637 257085 39671 257113
rect 39699 257085 39747 257113
rect 39437 257051 39747 257085
rect 39437 257023 39485 257051
rect 39513 257023 39547 257051
rect 39575 257023 39609 257051
rect 39637 257023 39671 257051
rect 39699 257023 39747 257051
rect 39437 256989 39747 257023
rect 39437 256961 39485 256989
rect 39513 256961 39547 256989
rect 39575 256961 39609 256989
rect 39637 256961 39671 256989
rect 39699 256961 39747 256989
rect 39437 248175 39747 256961
rect 39437 248147 39485 248175
rect 39513 248147 39547 248175
rect 39575 248147 39609 248175
rect 39637 248147 39671 248175
rect 39699 248147 39747 248175
rect 39437 248113 39747 248147
rect 39437 248085 39485 248113
rect 39513 248085 39547 248113
rect 39575 248085 39609 248113
rect 39637 248085 39671 248113
rect 39699 248085 39747 248113
rect 39437 248051 39747 248085
rect 39437 248023 39485 248051
rect 39513 248023 39547 248051
rect 39575 248023 39609 248051
rect 39637 248023 39671 248051
rect 39699 248023 39747 248051
rect 39437 247989 39747 248023
rect 39437 247961 39485 247989
rect 39513 247961 39547 247989
rect 39575 247961 39609 247989
rect 39637 247961 39671 247989
rect 39699 247961 39747 247989
rect 39437 239175 39747 247961
rect 39437 239147 39485 239175
rect 39513 239147 39547 239175
rect 39575 239147 39609 239175
rect 39637 239147 39671 239175
rect 39699 239147 39747 239175
rect 39437 239113 39747 239147
rect 39437 239085 39485 239113
rect 39513 239085 39547 239113
rect 39575 239085 39609 239113
rect 39637 239085 39671 239113
rect 39699 239085 39747 239113
rect 39437 239051 39747 239085
rect 39437 239023 39485 239051
rect 39513 239023 39547 239051
rect 39575 239023 39609 239051
rect 39637 239023 39671 239051
rect 39699 239023 39747 239051
rect 39437 238989 39747 239023
rect 39437 238961 39485 238989
rect 39513 238961 39547 238989
rect 39575 238961 39609 238989
rect 39637 238961 39671 238989
rect 39699 238961 39747 238989
rect 39437 230175 39747 238961
rect 39437 230147 39485 230175
rect 39513 230147 39547 230175
rect 39575 230147 39609 230175
rect 39637 230147 39671 230175
rect 39699 230147 39747 230175
rect 39437 230113 39747 230147
rect 39437 230085 39485 230113
rect 39513 230085 39547 230113
rect 39575 230085 39609 230113
rect 39637 230085 39671 230113
rect 39699 230085 39747 230113
rect 39437 230051 39747 230085
rect 39437 230023 39485 230051
rect 39513 230023 39547 230051
rect 39575 230023 39609 230051
rect 39637 230023 39671 230051
rect 39699 230023 39747 230051
rect 39437 229989 39747 230023
rect 39437 229961 39485 229989
rect 39513 229961 39547 229989
rect 39575 229961 39609 229989
rect 39637 229961 39671 229989
rect 39699 229961 39747 229989
rect 39437 221175 39747 229961
rect 39437 221147 39485 221175
rect 39513 221147 39547 221175
rect 39575 221147 39609 221175
rect 39637 221147 39671 221175
rect 39699 221147 39747 221175
rect 39437 221113 39747 221147
rect 39437 221085 39485 221113
rect 39513 221085 39547 221113
rect 39575 221085 39609 221113
rect 39637 221085 39671 221113
rect 39699 221085 39747 221113
rect 39437 221051 39747 221085
rect 39437 221023 39485 221051
rect 39513 221023 39547 221051
rect 39575 221023 39609 221051
rect 39637 221023 39671 221051
rect 39699 221023 39747 221051
rect 39437 220989 39747 221023
rect 39437 220961 39485 220989
rect 39513 220961 39547 220989
rect 39575 220961 39609 220989
rect 39637 220961 39671 220989
rect 39699 220961 39747 220989
rect 39437 212175 39747 220961
rect 39437 212147 39485 212175
rect 39513 212147 39547 212175
rect 39575 212147 39609 212175
rect 39637 212147 39671 212175
rect 39699 212147 39747 212175
rect 39437 212113 39747 212147
rect 39437 212085 39485 212113
rect 39513 212085 39547 212113
rect 39575 212085 39609 212113
rect 39637 212085 39671 212113
rect 39699 212085 39747 212113
rect 39437 212051 39747 212085
rect 39437 212023 39485 212051
rect 39513 212023 39547 212051
rect 39575 212023 39609 212051
rect 39637 212023 39671 212051
rect 39699 212023 39747 212051
rect 39437 211989 39747 212023
rect 39437 211961 39485 211989
rect 39513 211961 39547 211989
rect 39575 211961 39609 211989
rect 39637 211961 39671 211989
rect 39699 211961 39747 211989
rect 39437 203175 39747 211961
rect 39437 203147 39485 203175
rect 39513 203147 39547 203175
rect 39575 203147 39609 203175
rect 39637 203147 39671 203175
rect 39699 203147 39747 203175
rect 39437 203113 39747 203147
rect 39437 203085 39485 203113
rect 39513 203085 39547 203113
rect 39575 203085 39609 203113
rect 39637 203085 39671 203113
rect 39699 203085 39747 203113
rect 39437 203051 39747 203085
rect 39437 203023 39485 203051
rect 39513 203023 39547 203051
rect 39575 203023 39609 203051
rect 39637 203023 39671 203051
rect 39699 203023 39747 203051
rect 39437 202989 39747 203023
rect 39437 202961 39485 202989
rect 39513 202961 39547 202989
rect 39575 202961 39609 202989
rect 39637 202961 39671 202989
rect 39699 202961 39747 202989
rect 39437 194175 39747 202961
rect 39437 194147 39485 194175
rect 39513 194147 39547 194175
rect 39575 194147 39609 194175
rect 39637 194147 39671 194175
rect 39699 194147 39747 194175
rect 39437 194113 39747 194147
rect 39437 194085 39485 194113
rect 39513 194085 39547 194113
rect 39575 194085 39609 194113
rect 39637 194085 39671 194113
rect 39699 194085 39747 194113
rect 39437 194051 39747 194085
rect 39437 194023 39485 194051
rect 39513 194023 39547 194051
rect 39575 194023 39609 194051
rect 39637 194023 39671 194051
rect 39699 194023 39747 194051
rect 39437 193989 39747 194023
rect 39437 193961 39485 193989
rect 39513 193961 39547 193989
rect 39575 193961 39609 193989
rect 39637 193961 39671 193989
rect 39699 193961 39747 193989
rect 39437 185175 39747 193961
rect 39437 185147 39485 185175
rect 39513 185147 39547 185175
rect 39575 185147 39609 185175
rect 39637 185147 39671 185175
rect 39699 185147 39747 185175
rect 39437 185113 39747 185147
rect 39437 185085 39485 185113
rect 39513 185085 39547 185113
rect 39575 185085 39609 185113
rect 39637 185085 39671 185113
rect 39699 185085 39747 185113
rect 39437 185051 39747 185085
rect 39437 185023 39485 185051
rect 39513 185023 39547 185051
rect 39575 185023 39609 185051
rect 39637 185023 39671 185051
rect 39699 185023 39747 185051
rect 39437 184989 39747 185023
rect 39437 184961 39485 184989
rect 39513 184961 39547 184989
rect 39575 184961 39609 184989
rect 39637 184961 39671 184989
rect 39699 184961 39747 184989
rect 39437 176175 39747 184961
rect 39437 176147 39485 176175
rect 39513 176147 39547 176175
rect 39575 176147 39609 176175
rect 39637 176147 39671 176175
rect 39699 176147 39747 176175
rect 39437 176113 39747 176147
rect 39437 176085 39485 176113
rect 39513 176085 39547 176113
rect 39575 176085 39609 176113
rect 39637 176085 39671 176113
rect 39699 176085 39747 176113
rect 39437 176051 39747 176085
rect 39437 176023 39485 176051
rect 39513 176023 39547 176051
rect 39575 176023 39609 176051
rect 39637 176023 39671 176051
rect 39699 176023 39747 176051
rect 39437 175989 39747 176023
rect 39437 175961 39485 175989
rect 39513 175961 39547 175989
rect 39575 175961 39609 175989
rect 39637 175961 39671 175989
rect 39699 175961 39747 175989
rect 39437 167175 39747 175961
rect 39437 167147 39485 167175
rect 39513 167147 39547 167175
rect 39575 167147 39609 167175
rect 39637 167147 39671 167175
rect 39699 167147 39747 167175
rect 39437 167113 39747 167147
rect 39437 167085 39485 167113
rect 39513 167085 39547 167113
rect 39575 167085 39609 167113
rect 39637 167085 39671 167113
rect 39699 167085 39747 167113
rect 39437 167051 39747 167085
rect 39437 167023 39485 167051
rect 39513 167023 39547 167051
rect 39575 167023 39609 167051
rect 39637 167023 39671 167051
rect 39699 167023 39747 167051
rect 39437 166989 39747 167023
rect 39437 166961 39485 166989
rect 39513 166961 39547 166989
rect 39575 166961 39609 166989
rect 39637 166961 39671 166989
rect 39699 166961 39747 166989
rect 39437 158175 39747 166961
rect 39437 158147 39485 158175
rect 39513 158147 39547 158175
rect 39575 158147 39609 158175
rect 39637 158147 39671 158175
rect 39699 158147 39747 158175
rect 39437 158113 39747 158147
rect 39437 158085 39485 158113
rect 39513 158085 39547 158113
rect 39575 158085 39609 158113
rect 39637 158085 39671 158113
rect 39699 158085 39747 158113
rect 39437 158051 39747 158085
rect 39437 158023 39485 158051
rect 39513 158023 39547 158051
rect 39575 158023 39609 158051
rect 39637 158023 39671 158051
rect 39699 158023 39747 158051
rect 39437 157989 39747 158023
rect 39437 157961 39485 157989
rect 39513 157961 39547 157989
rect 39575 157961 39609 157989
rect 39637 157961 39671 157989
rect 39699 157961 39747 157989
rect 39437 149175 39747 157961
rect 39437 149147 39485 149175
rect 39513 149147 39547 149175
rect 39575 149147 39609 149175
rect 39637 149147 39671 149175
rect 39699 149147 39747 149175
rect 39437 149113 39747 149147
rect 39437 149085 39485 149113
rect 39513 149085 39547 149113
rect 39575 149085 39609 149113
rect 39637 149085 39671 149113
rect 39699 149085 39747 149113
rect 39437 149051 39747 149085
rect 39437 149023 39485 149051
rect 39513 149023 39547 149051
rect 39575 149023 39609 149051
rect 39637 149023 39671 149051
rect 39699 149023 39747 149051
rect 39437 148989 39747 149023
rect 39437 148961 39485 148989
rect 39513 148961 39547 148989
rect 39575 148961 39609 148989
rect 39637 148961 39671 148989
rect 39699 148961 39747 148989
rect 39437 140175 39747 148961
rect 39437 140147 39485 140175
rect 39513 140147 39547 140175
rect 39575 140147 39609 140175
rect 39637 140147 39671 140175
rect 39699 140147 39747 140175
rect 39437 140113 39747 140147
rect 39437 140085 39485 140113
rect 39513 140085 39547 140113
rect 39575 140085 39609 140113
rect 39637 140085 39671 140113
rect 39699 140085 39747 140113
rect 39437 140051 39747 140085
rect 39437 140023 39485 140051
rect 39513 140023 39547 140051
rect 39575 140023 39609 140051
rect 39637 140023 39671 140051
rect 39699 140023 39747 140051
rect 39437 139989 39747 140023
rect 39437 139961 39485 139989
rect 39513 139961 39547 139989
rect 39575 139961 39609 139989
rect 39637 139961 39671 139989
rect 39699 139961 39747 139989
rect 39437 131175 39747 139961
rect 39437 131147 39485 131175
rect 39513 131147 39547 131175
rect 39575 131147 39609 131175
rect 39637 131147 39671 131175
rect 39699 131147 39747 131175
rect 39437 131113 39747 131147
rect 39437 131085 39485 131113
rect 39513 131085 39547 131113
rect 39575 131085 39609 131113
rect 39637 131085 39671 131113
rect 39699 131085 39747 131113
rect 39437 131051 39747 131085
rect 39437 131023 39485 131051
rect 39513 131023 39547 131051
rect 39575 131023 39609 131051
rect 39637 131023 39671 131051
rect 39699 131023 39747 131051
rect 39437 130989 39747 131023
rect 39437 130961 39485 130989
rect 39513 130961 39547 130989
rect 39575 130961 39609 130989
rect 39637 130961 39671 130989
rect 39699 130961 39747 130989
rect 39437 122175 39747 130961
rect 39437 122147 39485 122175
rect 39513 122147 39547 122175
rect 39575 122147 39609 122175
rect 39637 122147 39671 122175
rect 39699 122147 39747 122175
rect 39437 122113 39747 122147
rect 39437 122085 39485 122113
rect 39513 122085 39547 122113
rect 39575 122085 39609 122113
rect 39637 122085 39671 122113
rect 39699 122085 39747 122113
rect 39437 122051 39747 122085
rect 39437 122023 39485 122051
rect 39513 122023 39547 122051
rect 39575 122023 39609 122051
rect 39637 122023 39671 122051
rect 39699 122023 39747 122051
rect 39437 121989 39747 122023
rect 39437 121961 39485 121989
rect 39513 121961 39547 121989
rect 39575 121961 39609 121989
rect 39637 121961 39671 121989
rect 39699 121961 39747 121989
rect 39437 113175 39747 121961
rect 39437 113147 39485 113175
rect 39513 113147 39547 113175
rect 39575 113147 39609 113175
rect 39637 113147 39671 113175
rect 39699 113147 39747 113175
rect 39437 113113 39747 113147
rect 39437 113085 39485 113113
rect 39513 113085 39547 113113
rect 39575 113085 39609 113113
rect 39637 113085 39671 113113
rect 39699 113085 39747 113113
rect 39437 113051 39747 113085
rect 39437 113023 39485 113051
rect 39513 113023 39547 113051
rect 39575 113023 39609 113051
rect 39637 113023 39671 113051
rect 39699 113023 39747 113051
rect 39437 112989 39747 113023
rect 39437 112961 39485 112989
rect 39513 112961 39547 112989
rect 39575 112961 39609 112989
rect 39637 112961 39671 112989
rect 39699 112961 39747 112989
rect 39437 104175 39747 112961
rect 39437 104147 39485 104175
rect 39513 104147 39547 104175
rect 39575 104147 39609 104175
rect 39637 104147 39671 104175
rect 39699 104147 39747 104175
rect 39437 104113 39747 104147
rect 39437 104085 39485 104113
rect 39513 104085 39547 104113
rect 39575 104085 39609 104113
rect 39637 104085 39671 104113
rect 39699 104085 39747 104113
rect 39437 104051 39747 104085
rect 39437 104023 39485 104051
rect 39513 104023 39547 104051
rect 39575 104023 39609 104051
rect 39637 104023 39671 104051
rect 39699 104023 39747 104051
rect 39437 103989 39747 104023
rect 39437 103961 39485 103989
rect 39513 103961 39547 103989
rect 39575 103961 39609 103989
rect 39637 103961 39671 103989
rect 39699 103961 39747 103989
rect 39437 95175 39747 103961
rect 39437 95147 39485 95175
rect 39513 95147 39547 95175
rect 39575 95147 39609 95175
rect 39637 95147 39671 95175
rect 39699 95147 39747 95175
rect 39437 95113 39747 95147
rect 39437 95085 39485 95113
rect 39513 95085 39547 95113
rect 39575 95085 39609 95113
rect 39637 95085 39671 95113
rect 39699 95085 39747 95113
rect 39437 95051 39747 95085
rect 39437 95023 39485 95051
rect 39513 95023 39547 95051
rect 39575 95023 39609 95051
rect 39637 95023 39671 95051
rect 39699 95023 39747 95051
rect 39437 94989 39747 95023
rect 39437 94961 39485 94989
rect 39513 94961 39547 94989
rect 39575 94961 39609 94989
rect 39637 94961 39671 94989
rect 39699 94961 39747 94989
rect 39437 86175 39747 94961
rect 39437 86147 39485 86175
rect 39513 86147 39547 86175
rect 39575 86147 39609 86175
rect 39637 86147 39671 86175
rect 39699 86147 39747 86175
rect 39437 86113 39747 86147
rect 39437 86085 39485 86113
rect 39513 86085 39547 86113
rect 39575 86085 39609 86113
rect 39637 86085 39671 86113
rect 39699 86085 39747 86113
rect 39437 86051 39747 86085
rect 39437 86023 39485 86051
rect 39513 86023 39547 86051
rect 39575 86023 39609 86051
rect 39637 86023 39671 86051
rect 39699 86023 39747 86051
rect 39437 85989 39747 86023
rect 39437 85961 39485 85989
rect 39513 85961 39547 85989
rect 39575 85961 39609 85989
rect 39637 85961 39671 85989
rect 39699 85961 39747 85989
rect 39437 77175 39747 85961
rect 39437 77147 39485 77175
rect 39513 77147 39547 77175
rect 39575 77147 39609 77175
rect 39637 77147 39671 77175
rect 39699 77147 39747 77175
rect 39437 77113 39747 77147
rect 39437 77085 39485 77113
rect 39513 77085 39547 77113
rect 39575 77085 39609 77113
rect 39637 77085 39671 77113
rect 39699 77085 39747 77113
rect 39437 77051 39747 77085
rect 39437 77023 39485 77051
rect 39513 77023 39547 77051
rect 39575 77023 39609 77051
rect 39637 77023 39671 77051
rect 39699 77023 39747 77051
rect 39437 76989 39747 77023
rect 39437 76961 39485 76989
rect 39513 76961 39547 76989
rect 39575 76961 39609 76989
rect 39637 76961 39671 76989
rect 39699 76961 39747 76989
rect 39437 68175 39747 76961
rect 39437 68147 39485 68175
rect 39513 68147 39547 68175
rect 39575 68147 39609 68175
rect 39637 68147 39671 68175
rect 39699 68147 39747 68175
rect 39437 68113 39747 68147
rect 39437 68085 39485 68113
rect 39513 68085 39547 68113
rect 39575 68085 39609 68113
rect 39637 68085 39671 68113
rect 39699 68085 39747 68113
rect 39437 68051 39747 68085
rect 39437 68023 39485 68051
rect 39513 68023 39547 68051
rect 39575 68023 39609 68051
rect 39637 68023 39671 68051
rect 39699 68023 39747 68051
rect 39437 67989 39747 68023
rect 39437 67961 39485 67989
rect 39513 67961 39547 67989
rect 39575 67961 39609 67989
rect 39637 67961 39671 67989
rect 39699 67961 39747 67989
rect 39437 59175 39747 67961
rect 39437 59147 39485 59175
rect 39513 59147 39547 59175
rect 39575 59147 39609 59175
rect 39637 59147 39671 59175
rect 39699 59147 39747 59175
rect 39437 59113 39747 59147
rect 39437 59085 39485 59113
rect 39513 59085 39547 59113
rect 39575 59085 39609 59113
rect 39637 59085 39671 59113
rect 39699 59085 39747 59113
rect 39437 59051 39747 59085
rect 39437 59023 39485 59051
rect 39513 59023 39547 59051
rect 39575 59023 39609 59051
rect 39637 59023 39671 59051
rect 39699 59023 39747 59051
rect 39437 58989 39747 59023
rect 39437 58961 39485 58989
rect 39513 58961 39547 58989
rect 39575 58961 39609 58989
rect 39637 58961 39671 58989
rect 39699 58961 39747 58989
rect 39437 50175 39747 58961
rect 39437 50147 39485 50175
rect 39513 50147 39547 50175
rect 39575 50147 39609 50175
rect 39637 50147 39671 50175
rect 39699 50147 39747 50175
rect 39437 50113 39747 50147
rect 39437 50085 39485 50113
rect 39513 50085 39547 50113
rect 39575 50085 39609 50113
rect 39637 50085 39671 50113
rect 39699 50085 39747 50113
rect 39437 50051 39747 50085
rect 39437 50023 39485 50051
rect 39513 50023 39547 50051
rect 39575 50023 39609 50051
rect 39637 50023 39671 50051
rect 39699 50023 39747 50051
rect 39437 49989 39747 50023
rect 39437 49961 39485 49989
rect 39513 49961 39547 49989
rect 39575 49961 39609 49989
rect 39637 49961 39671 49989
rect 39699 49961 39747 49989
rect 39437 41175 39747 49961
rect 39437 41147 39485 41175
rect 39513 41147 39547 41175
rect 39575 41147 39609 41175
rect 39637 41147 39671 41175
rect 39699 41147 39747 41175
rect 39437 41113 39747 41147
rect 39437 41085 39485 41113
rect 39513 41085 39547 41113
rect 39575 41085 39609 41113
rect 39637 41085 39671 41113
rect 39699 41085 39747 41113
rect 39437 41051 39747 41085
rect 39437 41023 39485 41051
rect 39513 41023 39547 41051
rect 39575 41023 39609 41051
rect 39637 41023 39671 41051
rect 39699 41023 39747 41051
rect 39437 40989 39747 41023
rect 39437 40961 39485 40989
rect 39513 40961 39547 40989
rect 39575 40961 39609 40989
rect 39637 40961 39671 40989
rect 39699 40961 39747 40989
rect 39437 32175 39747 40961
rect 39437 32147 39485 32175
rect 39513 32147 39547 32175
rect 39575 32147 39609 32175
rect 39637 32147 39671 32175
rect 39699 32147 39747 32175
rect 39437 32113 39747 32147
rect 39437 32085 39485 32113
rect 39513 32085 39547 32113
rect 39575 32085 39609 32113
rect 39637 32085 39671 32113
rect 39699 32085 39747 32113
rect 39437 32051 39747 32085
rect 39437 32023 39485 32051
rect 39513 32023 39547 32051
rect 39575 32023 39609 32051
rect 39637 32023 39671 32051
rect 39699 32023 39747 32051
rect 39437 31989 39747 32023
rect 39437 31961 39485 31989
rect 39513 31961 39547 31989
rect 39575 31961 39609 31989
rect 39637 31961 39671 31989
rect 39699 31961 39747 31989
rect 39437 23175 39747 31961
rect 39437 23147 39485 23175
rect 39513 23147 39547 23175
rect 39575 23147 39609 23175
rect 39637 23147 39671 23175
rect 39699 23147 39747 23175
rect 39437 23113 39747 23147
rect 39437 23085 39485 23113
rect 39513 23085 39547 23113
rect 39575 23085 39609 23113
rect 39637 23085 39671 23113
rect 39699 23085 39747 23113
rect 39437 23051 39747 23085
rect 39437 23023 39485 23051
rect 39513 23023 39547 23051
rect 39575 23023 39609 23051
rect 39637 23023 39671 23051
rect 39699 23023 39747 23051
rect 39437 22989 39747 23023
rect 39437 22961 39485 22989
rect 39513 22961 39547 22989
rect 39575 22961 39609 22989
rect 39637 22961 39671 22989
rect 39699 22961 39747 22989
rect 39437 14175 39747 22961
rect 39437 14147 39485 14175
rect 39513 14147 39547 14175
rect 39575 14147 39609 14175
rect 39637 14147 39671 14175
rect 39699 14147 39747 14175
rect 39437 14113 39747 14147
rect 39437 14085 39485 14113
rect 39513 14085 39547 14113
rect 39575 14085 39609 14113
rect 39637 14085 39671 14113
rect 39699 14085 39747 14113
rect 39437 14051 39747 14085
rect 39437 14023 39485 14051
rect 39513 14023 39547 14051
rect 39575 14023 39609 14051
rect 39637 14023 39671 14051
rect 39699 14023 39747 14051
rect 39437 13989 39747 14023
rect 39437 13961 39485 13989
rect 39513 13961 39547 13989
rect 39575 13961 39609 13989
rect 39637 13961 39671 13989
rect 39699 13961 39747 13989
rect 39437 5175 39747 13961
rect 39437 5147 39485 5175
rect 39513 5147 39547 5175
rect 39575 5147 39609 5175
rect 39637 5147 39671 5175
rect 39699 5147 39747 5175
rect 39437 5113 39747 5147
rect 39437 5085 39485 5113
rect 39513 5085 39547 5113
rect 39575 5085 39609 5113
rect 39637 5085 39671 5113
rect 39699 5085 39747 5113
rect 39437 5051 39747 5085
rect 39437 5023 39485 5051
rect 39513 5023 39547 5051
rect 39575 5023 39609 5051
rect 39637 5023 39671 5051
rect 39699 5023 39747 5051
rect 39437 4989 39747 5023
rect 39437 4961 39485 4989
rect 39513 4961 39547 4989
rect 39575 4961 39609 4989
rect 39637 4961 39671 4989
rect 39699 4961 39747 4989
rect 39437 -560 39747 4961
rect 39437 -588 39485 -560
rect 39513 -588 39547 -560
rect 39575 -588 39609 -560
rect 39637 -588 39671 -560
rect 39699 -588 39747 -560
rect 39437 -622 39747 -588
rect 39437 -650 39485 -622
rect 39513 -650 39547 -622
rect 39575 -650 39609 -622
rect 39637 -650 39671 -622
rect 39699 -650 39747 -622
rect 39437 -684 39747 -650
rect 39437 -712 39485 -684
rect 39513 -712 39547 -684
rect 39575 -712 39609 -684
rect 39637 -712 39671 -684
rect 39699 -712 39747 -684
rect 39437 -746 39747 -712
rect 39437 -774 39485 -746
rect 39513 -774 39547 -746
rect 39575 -774 39609 -746
rect 39637 -774 39671 -746
rect 39699 -774 39747 -746
rect 39437 -822 39747 -774
rect 46577 298606 46887 299134
rect 46577 298578 46625 298606
rect 46653 298578 46687 298606
rect 46715 298578 46749 298606
rect 46777 298578 46811 298606
rect 46839 298578 46887 298606
rect 46577 298544 46887 298578
rect 46577 298516 46625 298544
rect 46653 298516 46687 298544
rect 46715 298516 46749 298544
rect 46777 298516 46811 298544
rect 46839 298516 46887 298544
rect 46577 298482 46887 298516
rect 46577 298454 46625 298482
rect 46653 298454 46687 298482
rect 46715 298454 46749 298482
rect 46777 298454 46811 298482
rect 46839 298454 46887 298482
rect 46577 298420 46887 298454
rect 46577 298392 46625 298420
rect 46653 298392 46687 298420
rect 46715 298392 46749 298420
rect 46777 298392 46811 298420
rect 46839 298392 46887 298420
rect 46577 290175 46887 298392
rect 46577 290147 46625 290175
rect 46653 290147 46687 290175
rect 46715 290147 46749 290175
rect 46777 290147 46811 290175
rect 46839 290147 46887 290175
rect 46577 290113 46887 290147
rect 46577 290085 46625 290113
rect 46653 290085 46687 290113
rect 46715 290085 46749 290113
rect 46777 290085 46811 290113
rect 46839 290085 46887 290113
rect 46577 290051 46887 290085
rect 46577 290023 46625 290051
rect 46653 290023 46687 290051
rect 46715 290023 46749 290051
rect 46777 290023 46811 290051
rect 46839 290023 46887 290051
rect 46577 289989 46887 290023
rect 46577 289961 46625 289989
rect 46653 289961 46687 289989
rect 46715 289961 46749 289989
rect 46777 289961 46811 289989
rect 46839 289961 46887 289989
rect 46577 281175 46887 289961
rect 46577 281147 46625 281175
rect 46653 281147 46687 281175
rect 46715 281147 46749 281175
rect 46777 281147 46811 281175
rect 46839 281147 46887 281175
rect 46577 281113 46887 281147
rect 46577 281085 46625 281113
rect 46653 281085 46687 281113
rect 46715 281085 46749 281113
rect 46777 281085 46811 281113
rect 46839 281085 46887 281113
rect 46577 281051 46887 281085
rect 46577 281023 46625 281051
rect 46653 281023 46687 281051
rect 46715 281023 46749 281051
rect 46777 281023 46811 281051
rect 46839 281023 46887 281051
rect 46577 280989 46887 281023
rect 46577 280961 46625 280989
rect 46653 280961 46687 280989
rect 46715 280961 46749 280989
rect 46777 280961 46811 280989
rect 46839 280961 46887 280989
rect 46577 272175 46887 280961
rect 46577 272147 46625 272175
rect 46653 272147 46687 272175
rect 46715 272147 46749 272175
rect 46777 272147 46811 272175
rect 46839 272147 46887 272175
rect 46577 272113 46887 272147
rect 46577 272085 46625 272113
rect 46653 272085 46687 272113
rect 46715 272085 46749 272113
rect 46777 272085 46811 272113
rect 46839 272085 46887 272113
rect 46577 272051 46887 272085
rect 46577 272023 46625 272051
rect 46653 272023 46687 272051
rect 46715 272023 46749 272051
rect 46777 272023 46811 272051
rect 46839 272023 46887 272051
rect 46577 271989 46887 272023
rect 46577 271961 46625 271989
rect 46653 271961 46687 271989
rect 46715 271961 46749 271989
rect 46777 271961 46811 271989
rect 46839 271961 46887 271989
rect 46577 263175 46887 271961
rect 46577 263147 46625 263175
rect 46653 263147 46687 263175
rect 46715 263147 46749 263175
rect 46777 263147 46811 263175
rect 46839 263147 46887 263175
rect 46577 263113 46887 263147
rect 46577 263085 46625 263113
rect 46653 263085 46687 263113
rect 46715 263085 46749 263113
rect 46777 263085 46811 263113
rect 46839 263085 46887 263113
rect 46577 263051 46887 263085
rect 46577 263023 46625 263051
rect 46653 263023 46687 263051
rect 46715 263023 46749 263051
rect 46777 263023 46811 263051
rect 46839 263023 46887 263051
rect 46577 262989 46887 263023
rect 46577 262961 46625 262989
rect 46653 262961 46687 262989
rect 46715 262961 46749 262989
rect 46777 262961 46811 262989
rect 46839 262961 46887 262989
rect 46577 254175 46887 262961
rect 46577 254147 46625 254175
rect 46653 254147 46687 254175
rect 46715 254147 46749 254175
rect 46777 254147 46811 254175
rect 46839 254147 46887 254175
rect 46577 254113 46887 254147
rect 46577 254085 46625 254113
rect 46653 254085 46687 254113
rect 46715 254085 46749 254113
rect 46777 254085 46811 254113
rect 46839 254085 46887 254113
rect 46577 254051 46887 254085
rect 46577 254023 46625 254051
rect 46653 254023 46687 254051
rect 46715 254023 46749 254051
rect 46777 254023 46811 254051
rect 46839 254023 46887 254051
rect 46577 253989 46887 254023
rect 46577 253961 46625 253989
rect 46653 253961 46687 253989
rect 46715 253961 46749 253989
rect 46777 253961 46811 253989
rect 46839 253961 46887 253989
rect 46577 245175 46887 253961
rect 46577 245147 46625 245175
rect 46653 245147 46687 245175
rect 46715 245147 46749 245175
rect 46777 245147 46811 245175
rect 46839 245147 46887 245175
rect 46577 245113 46887 245147
rect 46577 245085 46625 245113
rect 46653 245085 46687 245113
rect 46715 245085 46749 245113
rect 46777 245085 46811 245113
rect 46839 245085 46887 245113
rect 46577 245051 46887 245085
rect 46577 245023 46625 245051
rect 46653 245023 46687 245051
rect 46715 245023 46749 245051
rect 46777 245023 46811 245051
rect 46839 245023 46887 245051
rect 46577 244989 46887 245023
rect 46577 244961 46625 244989
rect 46653 244961 46687 244989
rect 46715 244961 46749 244989
rect 46777 244961 46811 244989
rect 46839 244961 46887 244989
rect 46577 236175 46887 244961
rect 46577 236147 46625 236175
rect 46653 236147 46687 236175
rect 46715 236147 46749 236175
rect 46777 236147 46811 236175
rect 46839 236147 46887 236175
rect 46577 236113 46887 236147
rect 46577 236085 46625 236113
rect 46653 236085 46687 236113
rect 46715 236085 46749 236113
rect 46777 236085 46811 236113
rect 46839 236085 46887 236113
rect 46577 236051 46887 236085
rect 46577 236023 46625 236051
rect 46653 236023 46687 236051
rect 46715 236023 46749 236051
rect 46777 236023 46811 236051
rect 46839 236023 46887 236051
rect 46577 235989 46887 236023
rect 46577 235961 46625 235989
rect 46653 235961 46687 235989
rect 46715 235961 46749 235989
rect 46777 235961 46811 235989
rect 46839 235961 46887 235989
rect 46577 227175 46887 235961
rect 46577 227147 46625 227175
rect 46653 227147 46687 227175
rect 46715 227147 46749 227175
rect 46777 227147 46811 227175
rect 46839 227147 46887 227175
rect 46577 227113 46887 227147
rect 46577 227085 46625 227113
rect 46653 227085 46687 227113
rect 46715 227085 46749 227113
rect 46777 227085 46811 227113
rect 46839 227085 46887 227113
rect 46577 227051 46887 227085
rect 46577 227023 46625 227051
rect 46653 227023 46687 227051
rect 46715 227023 46749 227051
rect 46777 227023 46811 227051
rect 46839 227023 46887 227051
rect 46577 226989 46887 227023
rect 46577 226961 46625 226989
rect 46653 226961 46687 226989
rect 46715 226961 46749 226989
rect 46777 226961 46811 226989
rect 46839 226961 46887 226989
rect 46577 218175 46887 226961
rect 46577 218147 46625 218175
rect 46653 218147 46687 218175
rect 46715 218147 46749 218175
rect 46777 218147 46811 218175
rect 46839 218147 46887 218175
rect 46577 218113 46887 218147
rect 46577 218085 46625 218113
rect 46653 218085 46687 218113
rect 46715 218085 46749 218113
rect 46777 218085 46811 218113
rect 46839 218085 46887 218113
rect 46577 218051 46887 218085
rect 46577 218023 46625 218051
rect 46653 218023 46687 218051
rect 46715 218023 46749 218051
rect 46777 218023 46811 218051
rect 46839 218023 46887 218051
rect 46577 217989 46887 218023
rect 46577 217961 46625 217989
rect 46653 217961 46687 217989
rect 46715 217961 46749 217989
rect 46777 217961 46811 217989
rect 46839 217961 46887 217989
rect 46577 209175 46887 217961
rect 46577 209147 46625 209175
rect 46653 209147 46687 209175
rect 46715 209147 46749 209175
rect 46777 209147 46811 209175
rect 46839 209147 46887 209175
rect 46577 209113 46887 209147
rect 46577 209085 46625 209113
rect 46653 209085 46687 209113
rect 46715 209085 46749 209113
rect 46777 209085 46811 209113
rect 46839 209085 46887 209113
rect 46577 209051 46887 209085
rect 46577 209023 46625 209051
rect 46653 209023 46687 209051
rect 46715 209023 46749 209051
rect 46777 209023 46811 209051
rect 46839 209023 46887 209051
rect 46577 208989 46887 209023
rect 46577 208961 46625 208989
rect 46653 208961 46687 208989
rect 46715 208961 46749 208989
rect 46777 208961 46811 208989
rect 46839 208961 46887 208989
rect 46577 200175 46887 208961
rect 46577 200147 46625 200175
rect 46653 200147 46687 200175
rect 46715 200147 46749 200175
rect 46777 200147 46811 200175
rect 46839 200147 46887 200175
rect 46577 200113 46887 200147
rect 46577 200085 46625 200113
rect 46653 200085 46687 200113
rect 46715 200085 46749 200113
rect 46777 200085 46811 200113
rect 46839 200085 46887 200113
rect 46577 200051 46887 200085
rect 46577 200023 46625 200051
rect 46653 200023 46687 200051
rect 46715 200023 46749 200051
rect 46777 200023 46811 200051
rect 46839 200023 46887 200051
rect 46577 199989 46887 200023
rect 46577 199961 46625 199989
rect 46653 199961 46687 199989
rect 46715 199961 46749 199989
rect 46777 199961 46811 199989
rect 46839 199961 46887 199989
rect 46577 191175 46887 199961
rect 46577 191147 46625 191175
rect 46653 191147 46687 191175
rect 46715 191147 46749 191175
rect 46777 191147 46811 191175
rect 46839 191147 46887 191175
rect 46577 191113 46887 191147
rect 46577 191085 46625 191113
rect 46653 191085 46687 191113
rect 46715 191085 46749 191113
rect 46777 191085 46811 191113
rect 46839 191085 46887 191113
rect 46577 191051 46887 191085
rect 46577 191023 46625 191051
rect 46653 191023 46687 191051
rect 46715 191023 46749 191051
rect 46777 191023 46811 191051
rect 46839 191023 46887 191051
rect 46577 190989 46887 191023
rect 46577 190961 46625 190989
rect 46653 190961 46687 190989
rect 46715 190961 46749 190989
rect 46777 190961 46811 190989
rect 46839 190961 46887 190989
rect 46577 182175 46887 190961
rect 46577 182147 46625 182175
rect 46653 182147 46687 182175
rect 46715 182147 46749 182175
rect 46777 182147 46811 182175
rect 46839 182147 46887 182175
rect 46577 182113 46887 182147
rect 46577 182085 46625 182113
rect 46653 182085 46687 182113
rect 46715 182085 46749 182113
rect 46777 182085 46811 182113
rect 46839 182085 46887 182113
rect 46577 182051 46887 182085
rect 46577 182023 46625 182051
rect 46653 182023 46687 182051
rect 46715 182023 46749 182051
rect 46777 182023 46811 182051
rect 46839 182023 46887 182051
rect 46577 181989 46887 182023
rect 46577 181961 46625 181989
rect 46653 181961 46687 181989
rect 46715 181961 46749 181989
rect 46777 181961 46811 181989
rect 46839 181961 46887 181989
rect 46577 173175 46887 181961
rect 46577 173147 46625 173175
rect 46653 173147 46687 173175
rect 46715 173147 46749 173175
rect 46777 173147 46811 173175
rect 46839 173147 46887 173175
rect 46577 173113 46887 173147
rect 46577 173085 46625 173113
rect 46653 173085 46687 173113
rect 46715 173085 46749 173113
rect 46777 173085 46811 173113
rect 46839 173085 46887 173113
rect 46577 173051 46887 173085
rect 46577 173023 46625 173051
rect 46653 173023 46687 173051
rect 46715 173023 46749 173051
rect 46777 173023 46811 173051
rect 46839 173023 46887 173051
rect 46577 172989 46887 173023
rect 46577 172961 46625 172989
rect 46653 172961 46687 172989
rect 46715 172961 46749 172989
rect 46777 172961 46811 172989
rect 46839 172961 46887 172989
rect 46577 164175 46887 172961
rect 46577 164147 46625 164175
rect 46653 164147 46687 164175
rect 46715 164147 46749 164175
rect 46777 164147 46811 164175
rect 46839 164147 46887 164175
rect 46577 164113 46887 164147
rect 46577 164085 46625 164113
rect 46653 164085 46687 164113
rect 46715 164085 46749 164113
rect 46777 164085 46811 164113
rect 46839 164085 46887 164113
rect 46577 164051 46887 164085
rect 46577 164023 46625 164051
rect 46653 164023 46687 164051
rect 46715 164023 46749 164051
rect 46777 164023 46811 164051
rect 46839 164023 46887 164051
rect 46577 163989 46887 164023
rect 46577 163961 46625 163989
rect 46653 163961 46687 163989
rect 46715 163961 46749 163989
rect 46777 163961 46811 163989
rect 46839 163961 46887 163989
rect 46577 155175 46887 163961
rect 46577 155147 46625 155175
rect 46653 155147 46687 155175
rect 46715 155147 46749 155175
rect 46777 155147 46811 155175
rect 46839 155147 46887 155175
rect 46577 155113 46887 155147
rect 46577 155085 46625 155113
rect 46653 155085 46687 155113
rect 46715 155085 46749 155113
rect 46777 155085 46811 155113
rect 46839 155085 46887 155113
rect 46577 155051 46887 155085
rect 46577 155023 46625 155051
rect 46653 155023 46687 155051
rect 46715 155023 46749 155051
rect 46777 155023 46811 155051
rect 46839 155023 46887 155051
rect 46577 154989 46887 155023
rect 46577 154961 46625 154989
rect 46653 154961 46687 154989
rect 46715 154961 46749 154989
rect 46777 154961 46811 154989
rect 46839 154961 46887 154989
rect 46577 146175 46887 154961
rect 46577 146147 46625 146175
rect 46653 146147 46687 146175
rect 46715 146147 46749 146175
rect 46777 146147 46811 146175
rect 46839 146147 46887 146175
rect 46577 146113 46887 146147
rect 46577 146085 46625 146113
rect 46653 146085 46687 146113
rect 46715 146085 46749 146113
rect 46777 146085 46811 146113
rect 46839 146085 46887 146113
rect 46577 146051 46887 146085
rect 46577 146023 46625 146051
rect 46653 146023 46687 146051
rect 46715 146023 46749 146051
rect 46777 146023 46811 146051
rect 46839 146023 46887 146051
rect 46577 145989 46887 146023
rect 46577 145961 46625 145989
rect 46653 145961 46687 145989
rect 46715 145961 46749 145989
rect 46777 145961 46811 145989
rect 46839 145961 46887 145989
rect 46577 137175 46887 145961
rect 46577 137147 46625 137175
rect 46653 137147 46687 137175
rect 46715 137147 46749 137175
rect 46777 137147 46811 137175
rect 46839 137147 46887 137175
rect 46577 137113 46887 137147
rect 46577 137085 46625 137113
rect 46653 137085 46687 137113
rect 46715 137085 46749 137113
rect 46777 137085 46811 137113
rect 46839 137085 46887 137113
rect 46577 137051 46887 137085
rect 46577 137023 46625 137051
rect 46653 137023 46687 137051
rect 46715 137023 46749 137051
rect 46777 137023 46811 137051
rect 46839 137023 46887 137051
rect 46577 136989 46887 137023
rect 46577 136961 46625 136989
rect 46653 136961 46687 136989
rect 46715 136961 46749 136989
rect 46777 136961 46811 136989
rect 46839 136961 46887 136989
rect 46577 128175 46887 136961
rect 46577 128147 46625 128175
rect 46653 128147 46687 128175
rect 46715 128147 46749 128175
rect 46777 128147 46811 128175
rect 46839 128147 46887 128175
rect 46577 128113 46887 128147
rect 46577 128085 46625 128113
rect 46653 128085 46687 128113
rect 46715 128085 46749 128113
rect 46777 128085 46811 128113
rect 46839 128085 46887 128113
rect 46577 128051 46887 128085
rect 46577 128023 46625 128051
rect 46653 128023 46687 128051
rect 46715 128023 46749 128051
rect 46777 128023 46811 128051
rect 46839 128023 46887 128051
rect 46577 127989 46887 128023
rect 46577 127961 46625 127989
rect 46653 127961 46687 127989
rect 46715 127961 46749 127989
rect 46777 127961 46811 127989
rect 46839 127961 46887 127989
rect 46577 119175 46887 127961
rect 46577 119147 46625 119175
rect 46653 119147 46687 119175
rect 46715 119147 46749 119175
rect 46777 119147 46811 119175
rect 46839 119147 46887 119175
rect 46577 119113 46887 119147
rect 46577 119085 46625 119113
rect 46653 119085 46687 119113
rect 46715 119085 46749 119113
rect 46777 119085 46811 119113
rect 46839 119085 46887 119113
rect 46577 119051 46887 119085
rect 46577 119023 46625 119051
rect 46653 119023 46687 119051
rect 46715 119023 46749 119051
rect 46777 119023 46811 119051
rect 46839 119023 46887 119051
rect 46577 118989 46887 119023
rect 46577 118961 46625 118989
rect 46653 118961 46687 118989
rect 46715 118961 46749 118989
rect 46777 118961 46811 118989
rect 46839 118961 46887 118989
rect 46577 110175 46887 118961
rect 46577 110147 46625 110175
rect 46653 110147 46687 110175
rect 46715 110147 46749 110175
rect 46777 110147 46811 110175
rect 46839 110147 46887 110175
rect 46577 110113 46887 110147
rect 46577 110085 46625 110113
rect 46653 110085 46687 110113
rect 46715 110085 46749 110113
rect 46777 110085 46811 110113
rect 46839 110085 46887 110113
rect 46577 110051 46887 110085
rect 46577 110023 46625 110051
rect 46653 110023 46687 110051
rect 46715 110023 46749 110051
rect 46777 110023 46811 110051
rect 46839 110023 46887 110051
rect 46577 109989 46887 110023
rect 46577 109961 46625 109989
rect 46653 109961 46687 109989
rect 46715 109961 46749 109989
rect 46777 109961 46811 109989
rect 46839 109961 46887 109989
rect 46577 101175 46887 109961
rect 46577 101147 46625 101175
rect 46653 101147 46687 101175
rect 46715 101147 46749 101175
rect 46777 101147 46811 101175
rect 46839 101147 46887 101175
rect 46577 101113 46887 101147
rect 46577 101085 46625 101113
rect 46653 101085 46687 101113
rect 46715 101085 46749 101113
rect 46777 101085 46811 101113
rect 46839 101085 46887 101113
rect 46577 101051 46887 101085
rect 46577 101023 46625 101051
rect 46653 101023 46687 101051
rect 46715 101023 46749 101051
rect 46777 101023 46811 101051
rect 46839 101023 46887 101051
rect 46577 100989 46887 101023
rect 46577 100961 46625 100989
rect 46653 100961 46687 100989
rect 46715 100961 46749 100989
rect 46777 100961 46811 100989
rect 46839 100961 46887 100989
rect 46577 92175 46887 100961
rect 46577 92147 46625 92175
rect 46653 92147 46687 92175
rect 46715 92147 46749 92175
rect 46777 92147 46811 92175
rect 46839 92147 46887 92175
rect 46577 92113 46887 92147
rect 46577 92085 46625 92113
rect 46653 92085 46687 92113
rect 46715 92085 46749 92113
rect 46777 92085 46811 92113
rect 46839 92085 46887 92113
rect 46577 92051 46887 92085
rect 46577 92023 46625 92051
rect 46653 92023 46687 92051
rect 46715 92023 46749 92051
rect 46777 92023 46811 92051
rect 46839 92023 46887 92051
rect 46577 91989 46887 92023
rect 46577 91961 46625 91989
rect 46653 91961 46687 91989
rect 46715 91961 46749 91989
rect 46777 91961 46811 91989
rect 46839 91961 46887 91989
rect 46577 83175 46887 91961
rect 46577 83147 46625 83175
rect 46653 83147 46687 83175
rect 46715 83147 46749 83175
rect 46777 83147 46811 83175
rect 46839 83147 46887 83175
rect 46577 83113 46887 83147
rect 46577 83085 46625 83113
rect 46653 83085 46687 83113
rect 46715 83085 46749 83113
rect 46777 83085 46811 83113
rect 46839 83085 46887 83113
rect 46577 83051 46887 83085
rect 46577 83023 46625 83051
rect 46653 83023 46687 83051
rect 46715 83023 46749 83051
rect 46777 83023 46811 83051
rect 46839 83023 46887 83051
rect 46577 82989 46887 83023
rect 46577 82961 46625 82989
rect 46653 82961 46687 82989
rect 46715 82961 46749 82989
rect 46777 82961 46811 82989
rect 46839 82961 46887 82989
rect 46577 74175 46887 82961
rect 46577 74147 46625 74175
rect 46653 74147 46687 74175
rect 46715 74147 46749 74175
rect 46777 74147 46811 74175
rect 46839 74147 46887 74175
rect 46577 74113 46887 74147
rect 46577 74085 46625 74113
rect 46653 74085 46687 74113
rect 46715 74085 46749 74113
rect 46777 74085 46811 74113
rect 46839 74085 46887 74113
rect 46577 74051 46887 74085
rect 46577 74023 46625 74051
rect 46653 74023 46687 74051
rect 46715 74023 46749 74051
rect 46777 74023 46811 74051
rect 46839 74023 46887 74051
rect 46577 73989 46887 74023
rect 46577 73961 46625 73989
rect 46653 73961 46687 73989
rect 46715 73961 46749 73989
rect 46777 73961 46811 73989
rect 46839 73961 46887 73989
rect 46577 65175 46887 73961
rect 46577 65147 46625 65175
rect 46653 65147 46687 65175
rect 46715 65147 46749 65175
rect 46777 65147 46811 65175
rect 46839 65147 46887 65175
rect 46577 65113 46887 65147
rect 46577 65085 46625 65113
rect 46653 65085 46687 65113
rect 46715 65085 46749 65113
rect 46777 65085 46811 65113
rect 46839 65085 46887 65113
rect 46577 65051 46887 65085
rect 46577 65023 46625 65051
rect 46653 65023 46687 65051
rect 46715 65023 46749 65051
rect 46777 65023 46811 65051
rect 46839 65023 46887 65051
rect 46577 64989 46887 65023
rect 46577 64961 46625 64989
rect 46653 64961 46687 64989
rect 46715 64961 46749 64989
rect 46777 64961 46811 64989
rect 46839 64961 46887 64989
rect 46577 56175 46887 64961
rect 46577 56147 46625 56175
rect 46653 56147 46687 56175
rect 46715 56147 46749 56175
rect 46777 56147 46811 56175
rect 46839 56147 46887 56175
rect 46577 56113 46887 56147
rect 46577 56085 46625 56113
rect 46653 56085 46687 56113
rect 46715 56085 46749 56113
rect 46777 56085 46811 56113
rect 46839 56085 46887 56113
rect 46577 56051 46887 56085
rect 46577 56023 46625 56051
rect 46653 56023 46687 56051
rect 46715 56023 46749 56051
rect 46777 56023 46811 56051
rect 46839 56023 46887 56051
rect 46577 55989 46887 56023
rect 46577 55961 46625 55989
rect 46653 55961 46687 55989
rect 46715 55961 46749 55989
rect 46777 55961 46811 55989
rect 46839 55961 46887 55989
rect 46577 47175 46887 55961
rect 46577 47147 46625 47175
rect 46653 47147 46687 47175
rect 46715 47147 46749 47175
rect 46777 47147 46811 47175
rect 46839 47147 46887 47175
rect 46577 47113 46887 47147
rect 46577 47085 46625 47113
rect 46653 47085 46687 47113
rect 46715 47085 46749 47113
rect 46777 47085 46811 47113
rect 46839 47085 46887 47113
rect 46577 47051 46887 47085
rect 46577 47023 46625 47051
rect 46653 47023 46687 47051
rect 46715 47023 46749 47051
rect 46777 47023 46811 47051
rect 46839 47023 46887 47051
rect 46577 46989 46887 47023
rect 46577 46961 46625 46989
rect 46653 46961 46687 46989
rect 46715 46961 46749 46989
rect 46777 46961 46811 46989
rect 46839 46961 46887 46989
rect 46577 38175 46887 46961
rect 46577 38147 46625 38175
rect 46653 38147 46687 38175
rect 46715 38147 46749 38175
rect 46777 38147 46811 38175
rect 46839 38147 46887 38175
rect 46577 38113 46887 38147
rect 46577 38085 46625 38113
rect 46653 38085 46687 38113
rect 46715 38085 46749 38113
rect 46777 38085 46811 38113
rect 46839 38085 46887 38113
rect 46577 38051 46887 38085
rect 46577 38023 46625 38051
rect 46653 38023 46687 38051
rect 46715 38023 46749 38051
rect 46777 38023 46811 38051
rect 46839 38023 46887 38051
rect 46577 37989 46887 38023
rect 46577 37961 46625 37989
rect 46653 37961 46687 37989
rect 46715 37961 46749 37989
rect 46777 37961 46811 37989
rect 46839 37961 46887 37989
rect 46577 29175 46887 37961
rect 46577 29147 46625 29175
rect 46653 29147 46687 29175
rect 46715 29147 46749 29175
rect 46777 29147 46811 29175
rect 46839 29147 46887 29175
rect 46577 29113 46887 29147
rect 46577 29085 46625 29113
rect 46653 29085 46687 29113
rect 46715 29085 46749 29113
rect 46777 29085 46811 29113
rect 46839 29085 46887 29113
rect 46577 29051 46887 29085
rect 46577 29023 46625 29051
rect 46653 29023 46687 29051
rect 46715 29023 46749 29051
rect 46777 29023 46811 29051
rect 46839 29023 46887 29051
rect 46577 28989 46887 29023
rect 46577 28961 46625 28989
rect 46653 28961 46687 28989
rect 46715 28961 46749 28989
rect 46777 28961 46811 28989
rect 46839 28961 46887 28989
rect 46577 20175 46887 28961
rect 46577 20147 46625 20175
rect 46653 20147 46687 20175
rect 46715 20147 46749 20175
rect 46777 20147 46811 20175
rect 46839 20147 46887 20175
rect 46577 20113 46887 20147
rect 46577 20085 46625 20113
rect 46653 20085 46687 20113
rect 46715 20085 46749 20113
rect 46777 20085 46811 20113
rect 46839 20085 46887 20113
rect 46577 20051 46887 20085
rect 46577 20023 46625 20051
rect 46653 20023 46687 20051
rect 46715 20023 46749 20051
rect 46777 20023 46811 20051
rect 46839 20023 46887 20051
rect 46577 19989 46887 20023
rect 46577 19961 46625 19989
rect 46653 19961 46687 19989
rect 46715 19961 46749 19989
rect 46777 19961 46811 19989
rect 46839 19961 46887 19989
rect 46577 11175 46887 19961
rect 46577 11147 46625 11175
rect 46653 11147 46687 11175
rect 46715 11147 46749 11175
rect 46777 11147 46811 11175
rect 46839 11147 46887 11175
rect 46577 11113 46887 11147
rect 46577 11085 46625 11113
rect 46653 11085 46687 11113
rect 46715 11085 46749 11113
rect 46777 11085 46811 11113
rect 46839 11085 46887 11113
rect 46577 11051 46887 11085
rect 46577 11023 46625 11051
rect 46653 11023 46687 11051
rect 46715 11023 46749 11051
rect 46777 11023 46811 11051
rect 46839 11023 46887 11051
rect 46577 10989 46887 11023
rect 46577 10961 46625 10989
rect 46653 10961 46687 10989
rect 46715 10961 46749 10989
rect 46777 10961 46811 10989
rect 46839 10961 46887 10989
rect 46577 2175 46887 10961
rect 46577 2147 46625 2175
rect 46653 2147 46687 2175
rect 46715 2147 46749 2175
rect 46777 2147 46811 2175
rect 46839 2147 46887 2175
rect 46577 2113 46887 2147
rect 46577 2085 46625 2113
rect 46653 2085 46687 2113
rect 46715 2085 46749 2113
rect 46777 2085 46811 2113
rect 46839 2085 46887 2113
rect 46577 2051 46887 2085
rect 46577 2023 46625 2051
rect 46653 2023 46687 2051
rect 46715 2023 46749 2051
rect 46777 2023 46811 2051
rect 46839 2023 46887 2051
rect 46577 1989 46887 2023
rect 46577 1961 46625 1989
rect 46653 1961 46687 1989
rect 46715 1961 46749 1989
rect 46777 1961 46811 1989
rect 46839 1961 46887 1989
rect 46577 -80 46887 1961
rect 46577 -108 46625 -80
rect 46653 -108 46687 -80
rect 46715 -108 46749 -80
rect 46777 -108 46811 -80
rect 46839 -108 46887 -80
rect 46577 -142 46887 -108
rect 46577 -170 46625 -142
rect 46653 -170 46687 -142
rect 46715 -170 46749 -142
rect 46777 -170 46811 -142
rect 46839 -170 46887 -142
rect 46577 -204 46887 -170
rect 46577 -232 46625 -204
rect 46653 -232 46687 -204
rect 46715 -232 46749 -204
rect 46777 -232 46811 -204
rect 46839 -232 46887 -204
rect 46577 -266 46887 -232
rect 46577 -294 46625 -266
rect 46653 -294 46687 -266
rect 46715 -294 46749 -266
rect 46777 -294 46811 -266
rect 46839 -294 46887 -266
rect 46577 -822 46887 -294
rect 48437 299086 48747 299134
rect 48437 299058 48485 299086
rect 48513 299058 48547 299086
rect 48575 299058 48609 299086
rect 48637 299058 48671 299086
rect 48699 299058 48747 299086
rect 48437 299024 48747 299058
rect 48437 298996 48485 299024
rect 48513 298996 48547 299024
rect 48575 298996 48609 299024
rect 48637 298996 48671 299024
rect 48699 298996 48747 299024
rect 48437 298962 48747 298996
rect 48437 298934 48485 298962
rect 48513 298934 48547 298962
rect 48575 298934 48609 298962
rect 48637 298934 48671 298962
rect 48699 298934 48747 298962
rect 48437 298900 48747 298934
rect 48437 298872 48485 298900
rect 48513 298872 48547 298900
rect 48575 298872 48609 298900
rect 48637 298872 48671 298900
rect 48699 298872 48747 298900
rect 48437 293175 48747 298872
rect 48437 293147 48485 293175
rect 48513 293147 48547 293175
rect 48575 293147 48609 293175
rect 48637 293147 48671 293175
rect 48699 293147 48747 293175
rect 48437 293113 48747 293147
rect 48437 293085 48485 293113
rect 48513 293085 48547 293113
rect 48575 293085 48609 293113
rect 48637 293085 48671 293113
rect 48699 293085 48747 293113
rect 48437 293051 48747 293085
rect 48437 293023 48485 293051
rect 48513 293023 48547 293051
rect 48575 293023 48609 293051
rect 48637 293023 48671 293051
rect 48699 293023 48747 293051
rect 48437 292989 48747 293023
rect 48437 292961 48485 292989
rect 48513 292961 48547 292989
rect 48575 292961 48609 292989
rect 48637 292961 48671 292989
rect 48699 292961 48747 292989
rect 48437 284175 48747 292961
rect 48437 284147 48485 284175
rect 48513 284147 48547 284175
rect 48575 284147 48609 284175
rect 48637 284147 48671 284175
rect 48699 284147 48747 284175
rect 48437 284113 48747 284147
rect 48437 284085 48485 284113
rect 48513 284085 48547 284113
rect 48575 284085 48609 284113
rect 48637 284085 48671 284113
rect 48699 284085 48747 284113
rect 48437 284051 48747 284085
rect 48437 284023 48485 284051
rect 48513 284023 48547 284051
rect 48575 284023 48609 284051
rect 48637 284023 48671 284051
rect 48699 284023 48747 284051
rect 48437 283989 48747 284023
rect 48437 283961 48485 283989
rect 48513 283961 48547 283989
rect 48575 283961 48609 283989
rect 48637 283961 48671 283989
rect 48699 283961 48747 283989
rect 48437 275175 48747 283961
rect 48437 275147 48485 275175
rect 48513 275147 48547 275175
rect 48575 275147 48609 275175
rect 48637 275147 48671 275175
rect 48699 275147 48747 275175
rect 48437 275113 48747 275147
rect 48437 275085 48485 275113
rect 48513 275085 48547 275113
rect 48575 275085 48609 275113
rect 48637 275085 48671 275113
rect 48699 275085 48747 275113
rect 48437 275051 48747 275085
rect 48437 275023 48485 275051
rect 48513 275023 48547 275051
rect 48575 275023 48609 275051
rect 48637 275023 48671 275051
rect 48699 275023 48747 275051
rect 48437 274989 48747 275023
rect 48437 274961 48485 274989
rect 48513 274961 48547 274989
rect 48575 274961 48609 274989
rect 48637 274961 48671 274989
rect 48699 274961 48747 274989
rect 48437 266175 48747 274961
rect 48437 266147 48485 266175
rect 48513 266147 48547 266175
rect 48575 266147 48609 266175
rect 48637 266147 48671 266175
rect 48699 266147 48747 266175
rect 48437 266113 48747 266147
rect 48437 266085 48485 266113
rect 48513 266085 48547 266113
rect 48575 266085 48609 266113
rect 48637 266085 48671 266113
rect 48699 266085 48747 266113
rect 48437 266051 48747 266085
rect 48437 266023 48485 266051
rect 48513 266023 48547 266051
rect 48575 266023 48609 266051
rect 48637 266023 48671 266051
rect 48699 266023 48747 266051
rect 48437 265989 48747 266023
rect 48437 265961 48485 265989
rect 48513 265961 48547 265989
rect 48575 265961 48609 265989
rect 48637 265961 48671 265989
rect 48699 265961 48747 265989
rect 48437 257175 48747 265961
rect 55577 298606 55887 299134
rect 55577 298578 55625 298606
rect 55653 298578 55687 298606
rect 55715 298578 55749 298606
rect 55777 298578 55811 298606
rect 55839 298578 55887 298606
rect 55577 298544 55887 298578
rect 55577 298516 55625 298544
rect 55653 298516 55687 298544
rect 55715 298516 55749 298544
rect 55777 298516 55811 298544
rect 55839 298516 55887 298544
rect 55577 298482 55887 298516
rect 55577 298454 55625 298482
rect 55653 298454 55687 298482
rect 55715 298454 55749 298482
rect 55777 298454 55811 298482
rect 55839 298454 55887 298482
rect 55577 298420 55887 298454
rect 55577 298392 55625 298420
rect 55653 298392 55687 298420
rect 55715 298392 55749 298420
rect 55777 298392 55811 298420
rect 55839 298392 55887 298420
rect 55577 290175 55887 298392
rect 55577 290147 55625 290175
rect 55653 290147 55687 290175
rect 55715 290147 55749 290175
rect 55777 290147 55811 290175
rect 55839 290147 55887 290175
rect 55577 290113 55887 290147
rect 55577 290085 55625 290113
rect 55653 290085 55687 290113
rect 55715 290085 55749 290113
rect 55777 290085 55811 290113
rect 55839 290085 55887 290113
rect 55577 290051 55887 290085
rect 55577 290023 55625 290051
rect 55653 290023 55687 290051
rect 55715 290023 55749 290051
rect 55777 290023 55811 290051
rect 55839 290023 55887 290051
rect 55577 289989 55887 290023
rect 55577 289961 55625 289989
rect 55653 289961 55687 289989
rect 55715 289961 55749 289989
rect 55777 289961 55811 289989
rect 55839 289961 55887 289989
rect 55577 281175 55887 289961
rect 55577 281147 55625 281175
rect 55653 281147 55687 281175
rect 55715 281147 55749 281175
rect 55777 281147 55811 281175
rect 55839 281147 55887 281175
rect 55577 281113 55887 281147
rect 55577 281085 55625 281113
rect 55653 281085 55687 281113
rect 55715 281085 55749 281113
rect 55777 281085 55811 281113
rect 55839 281085 55887 281113
rect 55577 281051 55887 281085
rect 55577 281023 55625 281051
rect 55653 281023 55687 281051
rect 55715 281023 55749 281051
rect 55777 281023 55811 281051
rect 55839 281023 55887 281051
rect 55577 280989 55887 281023
rect 55577 280961 55625 280989
rect 55653 280961 55687 280989
rect 55715 280961 55749 280989
rect 55777 280961 55811 280989
rect 55839 280961 55887 280989
rect 55577 272175 55887 280961
rect 55577 272147 55625 272175
rect 55653 272147 55687 272175
rect 55715 272147 55749 272175
rect 55777 272147 55811 272175
rect 55839 272147 55887 272175
rect 55577 272113 55887 272147
rect 55577 272085 55625 272113
rect 55653 272085 55687 272113
rect 55715 272085 55749 272113
rect 55777 272085 55811 272113
rect 55839 272085 55887 272113
rect 55577 272051 55887 272085
rect 55577 272023 55625 272051
rect 55653 272023 55687 272051
rect 55715 272023 55749 272051
rect 55777 272023 55811 272051
rect 55839 272023 55887 272051
rect 55577 271989 55887 272023
rect 55577 271961 55625 271989
rect 55653 271961 55687 271989
rect 55715 271961 55749 271989
rect 55777 271961 55811 271989
rect 55839 271961 55887 271989
rect 55577 263175 55887 271961
rect 55577 263147 55625 263175
rect 55653 263147 55687 263175
rect 55715 263147 55749 263175
rect 55777 263147 55811 263175
rect 55839 263147 55887 263175
rect 55577 263113 55887 263147
rect 55577 263085 55625 263113
rect 55653 263085 55687 263113
rect 55715 263085 55749 263113
rect 55777 263085 55811 263113
rect 55839 263085 55887 263113
rect 55577 263051 55887 263085
rect 55577 263023 55625 263051
rect 55653 263023 55687 263051
rect 55715 263023 55749 263051
rect 55777 263023 55811 263051
rect 55839 263023 55887 263051
rect 55577 262989 55887 263023
rect 55577 262961 55625 262989
rect 55653 262961 55687 262989
rect 55715 262961 55749 262989
rect 55777 262961 55811 262989
rect 55839 262961 55887 262989
rect 55577 260603 55887 262961
rect 57437 299086 57747 299134
rect 57437 299058 57485 299086
rect 57513 299058 57547 299086
rect 57575 299058 57609 299086
rect 57637 299058 57671 299086
rect 57699 299058 57747 299086
rect 57437 299024 57747 299058
rect 57437 298996 57485 299024
rect 57513 298996 57547 299024
rect 57575 298996 57609 299024
rect 57637 298996 57671 299024
rect 57699 298996 57747 299024
rect 57437 298962 57747 298996
rect 57437 298934 57485 298962
rect 57513 298934 57547 298962
rect 57575 298934 57609 298962
rect 57637 298934 57671 298962
rect 57699 298934 57747 298962
rect 57437 298900 57747 298934
rect 57437 298872 57485 298900
rect 57513 298872 57547 298900
rect 57575 298872 57609 298900
rect 57637 298872 57671 298900
rect 57699 298872 57747 298900
rect 57437 293175 57747 298872
rect 57437 293147 57485 293175
rect 57513 293147 57547 293175
rect 57575 293147 57609 293175
rect 57637 293147 57671 293175
rect 57699 293147 57747 293175
rect 57437 293113 57747 293147
rect 57437 293085 57485 293113
rect 57513 293085 57547 293113
rect 57575 293085 57609 293113
rect 57637 293085 57671 293113
rect 57699 293085 57747 293113
rect 57437 293051 57747 293085
rect 57437 293023 57485 293051
rect 57513 293023 57547 293051
rect 57575 293023 57609 293051
rect 57637 293023 57671 293051
rect 57699 293023 57747 293051
rect 57437 292989 57747 293023
rect 57437 292961 57485 292989
rect 57513 292961 57547 292989
rect 57575 292961 57609 292989
rect 57637 292961 57671 292989
rect 57699 292961 57747 292989
rect 57437 284175 57747 292961
rect 57437 284147 57485 284175
rect 57513 284147 57547 284175
rect 57575 284147 57609 284175
rect 57637 284147 57671 284175
rect 57699 284147 57747 284175
rect 57437 284113 57747 284147
rect 57437 284085 57485 284113
rect 57513 284085 57547 284113
rect 57575 284085 57609 284113
rect 57637 284085 57671 284113
rect 57699 284085 57747 284113
rect 57437 284051 57747 284085
rect 57437 284023 57485 284051
rect 57513 284023 57547 284051
rect 57575 284023 57609 284051
rect 57637 284023 57671 284051
rect 57699 284023 57747 284051
rect 57437 283989 57747 284023
rect 57437 283961 57485 283989
rect 57513 283961 57547 283989
rect 57575 283961 57609 283989
rect 57637 283961 57671 283989
rect 57699 283961 57747 283989
rect 57437 275175 57747 283961
rect 57437 275147 57485 275175
rect 57513 275147 57547 275175
rect 57575 275147 57609 275175
rect 57637 275147 57671 275175
rect 57699 275147 57747 275175
rect 57437 275113 57747 275147
rect 57437 275085 57485 275113
rect 57513 275085 57547 275113
rect 57575 275085 57609 275113
rect 57637 275085 57671 275113
rect 57699 275085 57747 275113
rect 57437 275051 57747 275085
rect 57437 275023 57485 275051
rect 57513 275023 57547 275051
rect 57575 275023 57609 275051
rect 57637 275023 57671 275051
rect 57699 275023 57747 275051
rect 57437 274989 57747 275023
rect 57437 274961 57485 274989
rect 57513 274961 57547 274989
rect 57575 274961 57609 274989
rect 57637 274961 57671 274989
rect 57699 274961 57747 274989
rect 57437 266175 57747 274961
rect 57437 266147 57485 266175
rect 57513 266147 57547 266175
rect 57575 266147 57609 266175
rect 57637 266147 57671 266175
rect 57699 266147 57747 266175
rect 57437 266113 57747 266147
rect 57437 266085 57485 266113
rect 57513 266085 57547 266113
rect 57575 266085 57609 266113
rect 57637 266085 57671 266113
rect 57699 266085 57747 266113
rect 57437 266051 57747 266085
rect 57437 266023 57485 266051
rect 57513 266023 57547 266051
rect 57575 266023 57609 266051
rect 57637 266023 57671 266051
rect 57699 266023 57747 266051
rect 57437 265989 57747 266023
rect 57437 265961 57485 265989
rect 57513 265961 57547 265989
rect 57575 265961 57609 265989
rect 57637 265961 57671 265989
rect 57699 265961 57747 265989
rect 57437 260603 57747 265961
rect 64577 298606 64887 299134
rect 64577 298578 64625 298606
rect 64653 298578 64687 298606
rect 64715 298578 64749 298606
rect 64777 298578 64811 298606
rect 64839 298578 64887 298606
rect 64577 298544 64887 298578
rect 64577 298516 64625 298544
rect 64653 298516 64687 298544
rect 64715 298516 64749 298544
rect 64777 298516 64811 298544
rect 64839 298516 64887 298544
rect 64577 298482 64887 298516
rect 64577 298454 64625 298482
rect 64653 298454 64687 298482
rect 64715 298454 64749 298482
rect 64777 298454 64811 298482
rect 64839 298454 64887 298482
rect 64577 298420 64887 298454
rect 64577 298392 64625 298420
rect 64653 298392 64687 298420
rect 64715 298392 64749 298420
rect 64777 298392 64811 298420
rect 64839 298392 64887 298420
rect 64577 290175 64887 298392
rect 64577 290147 64625 290175
rect 64653 290147 64687 290175
rect 64715 290147 64749 290175
rect 64777 290147 64811 290175
rect 64839 290147 64887 290175
rect 64577 290113 64887 290147
rect 64577 290085 64625 290113
rect 64653 290085 64687 290113
rect 64715 290085 64749 290113
rect 64777 290085 64811 290113
rect 64839 290085 64887 290113
rect 64577 290051 64887 290085
rect 64577 290023 64625 290051
rect 64653 290023 64687 290051
rect 64715 290023 64749 290051
rect 64777 290023 64811 290051
rect 64839 290023 64887 290051
rect 64577 289989 64887 290023
rect 64577 289961 64625 289989
rect 64653 289961 64687 289989
rect 64715 289961 64749 289989
rect 64777 289961 64811 289989
rect 64839 289961 64887 289989
rect 64577 281175 64887 289961
rect 64577 281147 64625 281175
rect 64653 281147 64687 281175
rect 64715 281147 64749 281175
rect 64777 281147 64811 281175
rect 64839 281147 64887 281175
rect 64577 281113 64887 281147
rect 64577 281085 64625 281113
rect 64653 281085 64687 281113
rect 64715 281085 64749 281113
rect 64777 281085 64811 281113
rect 64839 281085 64887 281113
rect 64577 281051 64887 281085
rect 64577 281023 64625 281051
rect 64653 281023 64687 281051
rect 64715 281023 64749 281051
rect 64777 281023 64811 281051
rect 64839 281023 64887 281051
rect 64577 280989 64887 281023
rect 64577 280961 64625 280989
rect 64653 280961 64687 280989
rect 64715 280961 64749 280989
rect 64777 280961 64811 280989
rect 64839 280961 64887 280989
rect 64577 272175 64887 280961
rect 64577 272147 64625 272175
rect 64653 272147 64687 272175
rect 64715 272147 64749 272175
rect 64777 272147 64811 272175
rect 64839 272147 64887 272175
rect 64577 272113 64887 272147
rect 64577 272085 64625 272113
rect 64653 272085 64687 272113
rect 64715 272085 64749 272113
rect 64777 272085 64811 272113
rect 64839 272085 64887 272113
rect 64577 272051 64887 272085
rect 64577 272023 64625 272051
rect 64653 272023 64687 272051
rect 64715 272023 64749 272051
rect 64777 272023 64811 272051
rect 64839 272023 64887 272051
rect 64577 271989 64887 272023
rect 64577 271961 64625 271989
rect 64653 271961 64687 271989
rect 64715 271961 64749 271989
rect 64777 271961 64811 271989
rect 64839 271961 64887 271989
rect 64577 263175 64887 271961
rect 64577 263147 64625 263175
rect 64653 263147 64687 263175
rect 64715 263147 64749 263175
rect 64777 263147 64811 263175
rect 64839 263147 64887 263175
rect 64577 263113 64887 263147
rect 64577 263085 64625 263113
rect 64653 263085 64687 263113
rect 64715 263085 64749 263113
rect 64777 263085 64811 263113
rect 64839 263085 64887 263113
rect 64577 263051 64887 263085
rect 64577 263023 64625 263051
rect 64653 263023 64687 263051
rect 64715 263023 64749 263051
rect 64777 263023 64811 263051
rect 64839 263023 64887 263051
rect 64577 262989 64887 263023
rect 64577 262961 64625 262989
rect 64653 262961 64687 262989
rect 64715 262961 64749 262989
rect 64777 262961 64811 262989
rect 64839 262961 64887 262989
rect 64577 260603 64887 262961
rect 66437 299086 66747 299134
rect 66437 299058 66485 299086
rect 66513 299058 66547 299086
rect 66575 299058 66609 299086
rect 66637 299058 66671 299086
rect 66699 299058 66747 299086
rect 66437 299024 66747 299058
rect 66437 298996 66485 299024
rect 66513 298996 66547 299024
rect 66575 298996 66609 299024
rect 66637 298996 66671 299024
rect 66699 298996 66747 299024
rect 66437 298962 66747 298996
rect 66437 298934 66485 298962
rect 66513 298934 66547 298962
rect 66575 298934 66609 298962
rect 66637 298934 66671 298962
rect 66699 298934 66747 298962
rect 66437 298900 66747 298934
rect 66437 298872 66485 298900
rect 66513 298872 66547 298900
rect 66575 298872 66609 298900
rect 66637 298872 66671 298900
rect 66699 298872 66747 298900
rect 66437 293175 66747 298872
rect 66437 293147 66485 293175
rect 66513 293147 66547 293175
rect 66575 293147 66609 293175
rect 66637 293147 66671 293175
rect 66699 293147 66747 293175
rect 66437 293113 66747 293147
rect 66437 293085 66485 293113
rect 66513 293085 66547 293113
rect 66575 293085 66609 293113
rect 66637 293085 66671 293113
rect 66699 293085 66747 293113
rect 66437 293051 66747 293085
rect 66437 293023 66485 293051
rect 66513 293023 66547 293051
rect 66575 293023 66609 293051
rect 66637 293023 66671 293051
rect 66699 293023 66747 293051
rect 66437 292989 66747 293023
rect 66437 292961 66485 292989
rect 66513 292961 66547 292989
rect 66575 292961 66609 292989
rect 66637 292961 66671 292989
rect 66699 292961 66747 292989
rect 66437 284175 66747 292961
rect 66437 284147 66485 284175
rect 66513 284147 66547 284175
rect 66575 284147 66609 284175
rect 66637 284147 66671 284175
rect 66699 284147 66747 284175
rect 66437 284113 66747 284147
rect 66437 284085 66485 284113
rect 66513 284085 66547 284113
rect 66575 284085 66609 284113
rect 66637 284085 66671 284113
rect 66699 284085 66747 284113
rect 66437 284051 66747 284085
rect 66437 284023 66485 284051
rect 66513 284023 66547 284051
rect 66575 284023 66609 284051
rect 66637 284023 66671 284051
rect 66699 284023 66747 284051
rect 66437 283989 66747 284023
rect 66437 283961 66485 283989
rect 66513 283961 66547 283989
rect 66575 283961 66609 283989
rect 66637 283961 66671 283989
rect 66699 283961 66747 283989
rect 66437 275175 66747 283961
rect 66437 275147 66485 275175
rect 66513 275147 66547 275175
rect 66575 275147 66609 275175
rect 66637 275147 66671 275175
rect 66699 275147 66747 275175
rect 66437 275113 66747 275147
rect 66437 275085 66485 275113
rect 66513 275085 66547 275113
rect 66575 275085 66609 275113
rect 66637 275085 66671 275113
rect 66699 275085 66747 275113
rect 66437 275051 66747 275085
rect 66437 275023 66485 275051
rect 66513 275023 66547 275051
rect 66575 275023 66609 275051
rect 66637 275023 66671 275051
rect 66699 275023 66747 275051
rect 66437 274989 66747 275023
rect 66437 274961 66485 274989
rect 66513 274961 66547 274989
rect 66575 274961 66609 274989
rect 66637 274961 66671 274989
rect 66699 274961 66747 274989
rect 66437 266175 66747 274961
rect 66437 266147 66485 266175
rect 66513 266147 66547 266175
rect 66575 266147 66609 266175
rect 66637 266147 66671 266175
rect 66699 266147 66747 266175
rect 66437 266113 66747 266147
rect 66437 266085 66485 266113
rect 66513 266085 66547 266113
rect 66575 266085 66609 266113
rect 66637 266085 66671 266113
rect 66699 266085 66747 266113
rect 66437 266051 66747 266085
rect 66437 266023 66485 266051
rect 66513 266023 66547 266051
rect 66575 266023 66609 266051
rect 66637 266023 66671 266051
rect 66699 266023 66747 266051
rect 66437 265989 66747 266023
rect 66437 265961 66485 265989
rect 66513 265961 66547 265989
rect 66575 265961 66609 265989
rect 66637 265961 66671 265989
rect 66699 265961 66747 265989
rect 66437 260603 66747 265961
rect 73577 298606 73887 299134
rect 73577 298578 73625 298606
rect 73653 298578 73687 298606
rect 73715 298578 73749 298606
rect 73777 298578 73811 298606
rect 73839 298578 73887 298606
rect 73577 298544 73887 298578
rect 73577 298516 73625 298544
rect 73653 298516 73687 298544
rect 73715 298516 73749 298544
rect 73777 298516 73811 298544
rect 73839 298516 73887 298544
rect 73577 298482 73887 298516
rect 73577 298454 73625 298482
rect 73653 298454 73687 298482
rect 73715 298454 73749 298482
rect 73777 298454 73811 298482
rect 73839 298454 73887 298482
rect 73577 298420 73887 298454
rect 73577 298392 73625 298420
rect 73653 298392 73687 298420
rect 73715 298392 73749 298420
rect 73777 298392 73811 298420
rect 73839 298392 73887 298420
rect 73577 290175 73887 298392
rect 73577 290147 73625 290175
rect 73653 290147 73687 290175
rect 73715 290147 73749 290175
rect 73777 290147 73811 290175
rect 73839 290147 73887 290175
rect 73577 290113 73887 290147
rect 73577 290085 73625 290113
rect 73653 290085 73687 290113
rect 73715 290085 73749 290113
rect 73777 290085 73811 290113
rect 73839 290085 73887 290113
rect 73577 290051 73887 290085
rect 73577 290023 73625 290051
rect 73653 290023 73687 290051
rect 73715 290023 73749 290051
rect 73777 290023 73811 290051
rect 73839 290023 73887 290051
rect 73577 289989 73887 290023
rect 73577 289961 73625 289989
rect 73653 289961 73687 289989
rect 73715 289961 73749 289989
rect 73777 289961 73811 289989
rect 73839 289961 73887 289989
rect 73577 281175 73887 289961
rect 73577 281147 73625 281175
rect 73653 281147 73687 281175
rect 73715 281147 73749 281175
rect 73777 281147 73811 281175
rect 73839 281147 73887 281175
rect 73577 281113 73887 281147
rect 73577 281085 73625 281113
rect 73653 281085 73687 281113
rect 73715 281085 73749 281113
rect 73777 281085 73811 281113
rect 73839 281085 73887 281113
rect 73577 281051 73887 281085
rect 73577 281023 73625 281051
rect 73653 281023 73687 281051
rect 73715 281023 73749 281051
rect 73777 281023 73811 281051
rect 73839 281023 73887 281051
rect 73577 280989 73887 281023
rect 73577 280961 73625 280989
rect 73653 280961 73687 280989
rect 73715 280961 73749 280989
rect 73777 280961 73811 280989
rect 73839 280961 73887 280989
rect 73577 272175 73887 280961
rect 73577 272147 73625 272175
rect 73653 272147 73687 272175
rect 73715 272147 73749 272175
rect 73777 272147 73811 272175
rect 73839 272147 73887 272175
rect 73577 272113 73887 272147
rect 73577 272085 73625 272113
rect 73653 272085 73687 272113
rect 73715 272085 73749 272113
rect 73777 272085 73811 272113
rect 73839 272085 73887 272113
rect 73577 272051 73887 272085
rect 73577 272023 73625 272051
rect 73653 272023 73687 272051
rect 73715 272023 73749 272051
rect 73777 272023 73811 272051
rect 73839 272023 73887 272051
rect 73577 271989 73887 272023
rect 73577 271961 73625 271989
rect 73653 271961 73687 271989
rect 73715 271961 73749 271989
rect 73777 271961 73811 271989
rect 73839 271961 73887 271989
rect 73577 263175 73887 271961
rect 73577 263147 73625 263175
rect 73653 263147 73687 263175
rect 73715 263147 73749 263175
rect 73777 263147 73811 263175
rect 73839 263147 73887 263175
rect 73577 263113 73887 263147
rect 73577 263085 73625 263113
rect 73653 263085 73687 263113
rect 73715 263085 73749 263113
rect 73777 263085 73811 263113
rect 73839 263085 73887 263113
rect 73577 263051 73887 263085
rect 73577 263023 73625 263051
rect 73653 263023 73687 263051
rect 73715 263023 73749 263051
rect 73777 263023 73811 263051
rect 73839 263023 73887 263051
rect 73577 262989 73887 263023
rect 73577 262961 73625 262989
rect 73653 262961 73687 262989
rect 73715 262961 73749 262989
rect 73777 262961 73811 262989
rect 73839 262961 73887 262989
rect 73577 260603 73887 262961
rect 75437 299086 75747 299134
rect 75437 299058 75485 299086
rect 75513 299058 75547 299086
rect 75575 299058 75609 299086
rect 75637 299058 75671 299086
rect 75699 299058 75747 299086
rect 75437 299024 75747 299058
rect 75437 298996 75485 299024
rect 75513 298996 75547 299024
rect 75575 298996 75609 299024
rect 75637 298996 75671 299024
rect 75699 298996 75747 299024
rect 75437 298962 75747 298996
rect 75437 298934 75485 298962
rect 75513 298934 75547 298962
rect 75575 298934 75609 298962
rect 75637 298934 75671 298962
rect 75699 298934 75747 298962
rect 75437 298900 75747 298934
rect 75437 298872 75485 298900
rect 75513 298872 75547 298900
rect 75575 298872 75609 298900
rect 75637 298872 75671 298900
rect 75699 298872 75747 298900
rect 75437 293175 75747 298872
rect 75437 293147 75485 293175
rect 75513 293147 75547 293175
rect 75575 293147 75609 293175
rect 75637 293147 75671 293175
rect 75699 293147 75747 293175
rect 75437 293113 75747 293147
rect 75437 293085 75485 293113
rect 75513 293085 75547 293113
rect 75575 293085 75609 293113
rect 75637 293085 75671 293113
rect 75699 293085 75747 293113
rect 75437 293051 75747 293085
rect 75437 293023 75485 293051
rect 75513 293023 75547 293051
rect 75575 293023 75609 293051
rect 75637 293023 75671 293051
rect 75699 293023 75747 293051
rect 75437 292989 75747 293023
rect 75437 292961 75485 292989
rect 75513 292961 75547 292989
rect 75575 292961 75609 292989
rect 75637 292961 75671 292989
rect 75699 292961 75747 292989
rect 75437 284175 75747 292961
rect 75437 284147 75485 284175
rect 75513 284147 75547 284175
rect 75575 284147 75609 284175
rect 75637 284147 75671 284175
rect 75699 284147 75747 284175
rect 75437 284113 75747 284147
rect 75437 284085 75485 284113
rect 75513 284085 75547 284113
rect 75575 284085 75609 284113
rect 75637 284085 75671 284113
rect 75699 284085 75747 284113
rect 75437 284051 75747 284085
rect 75437 284023 75485 284051
rect 75513 284023 75547 284051
rect 75575 284023 75609 284051
rect 75637 284023 75671 284051
rect 75699 284023 75747 284051
rect 75437 283989 75747 284023
rect 75437 283961 75485 283989
rect 75513 283961 75547 283989
rect 75575 283961 75609 283989
rect 75637 283961 75671 283989
rect 75699 283961 75747 283989
rect 75437 275175 75747 283961
rect 75437 275147 75485 275175
rect 75513 275147 75547 275175
rect 75575 275147 75609 275175
rect 75637 275147 75671 275175
rect 75699 275147 75747 275175
rect 75437 275113 75747 275147
rect 75437 275085 75485 275113
rect 75513 275085 75547 275113
rect 75575 275085 75609 275113
rect 75637 275085 75671 275113
rect 75699 275085 75747 275113
rect 75437 275051 75747 275085
rect 75437 275023 75485 275051
rect 75513 275023 75547 275051
rect 75575 275023 75609 275051
rect 75637 275023 75671 275051
rect 75699 275023 75747 275051
rect 75437 274989 75747 275023
rect 75437 274961 75485 274989
rect 75513 274961 75547 274989
rect 75575 274961 75609 274989
rect 75637 274961 75671 274989
rect 75699 274961 75747 274989
rect 75437 266175 75747 274961
rect 75437 266147 75485 266175
rect 75513 266147 75547 266175
rect 75575 266147 75609 266175
rect 75637 266147 75671 266175
rect 75699 266147 75747 266175
rect 75437 266113 75747 266147
rect 75437 266085 75485 266113
rect 75513 266085 75547 266113
rect 75575 266085 75609 266113
rect 75637 266085 75671 266113
rect 75699 266085 75747 266113
rect 75437 266051 75747 266085
rect 75437 266023 75485 266051
rect 75513 266023 75547 266051
rect 75575 266023 75609 266051
rect 75637 266023 75671 266051
rect 75699 266023 75747 266051
rect 75437 265989 75747 266023
rect 75437 265961 75485 265989
rect 75513 265961 75547 265989
rect 75575 265961 75609 265989
rect 75637 265961 75671 265989
rect 75699 265961 75747 265989
rect 75437 260603 75747 265961
rect 82577 298606 82887 299134
rect 82577 298578 82625 298606
rect 82653 298578 82687 298606
rect 82715 298578 82749 298606
rect 82777 298578 82811 298606
rect 82839 298578 82887 298606
rect 82577 298544 82887 298578
rect 82577 298516 82625 298544
rect 82653 298516 82687 298544
rect 82715 298516 82749 298544
rect 82777 298516 82811 298544
rect 82839 298516 82887 298544
rect 82577 298482 82887 298516
rect 82577 298454 82625 298482
rect 82653 298454 82687 298482
rect 82715 298454 82749 298482
rect 82777 298454 82811 298482
rect 82839 298454 82887 298482
rect 82577 298420 82887 298454
rect 82577 298392 82625 298420
rect 82653 298392 82687 298420
rect 82715 298392 82749 298420
rect 82777 298392 82811 298420
rect 82839 298392 82887 298420
rect 82577 290175 82887 298392
rect 82577 290147 82625 290175
rect 82653 290147 82687 290175
rect 82715 290147 82749 290175
rect 82777 290147 82811 290175
rect 82839 290147 82887 290175
rect 82577 290113 82887 290147
rect 82577 290085 82625 290113
rect 82653 290085 82687 290113
rect 82715 290085 82749 290113
rect 82777 290085 82811 290113
rect 82839 290085 82887 290113
rect 82577 290051 82887 290085
rect 82577 290023 82625 290051
rect 82653 290023 82687 290051
rect 82715 290023 82749 290051
rect 82777 290023 82811 290051
rect 82839 290023 82887 290051
rect 82577 289989 82887 290023
rect 82577 289961 82625 289989
rect 82653 289961 82687 289989
rect 82715 289961 82749 289989
rect 82777 289961 82811 289989
rect 82839 289961 82887 289989
rect 82577 281175 82887 289961
rect 82577 281147 82625 281175
rect 82653 281147 82687 281175
rect 82715 281147 82749 281175
rect 82777 281147 82811 281175
rect 82839 281147 82887 281175
rect 82577 281113 82887 281147
rect 82577 281085 82625 281113
rect 82653 281085 82687 281113
rect 82715 281085 82749 281113
rect 82777 281085 82811 281113
rect 82839 281085 82887 281113
rect 82577 281051 82887 281085
rect 82577 281023 82625 281051
rect 82653 281023 82687 281051
rect 82715 281023 82749 281051
rect 82777 281023 82811 281051
rect 82839 281023 82887 281051
rect 82577 280989 82887 281023
rect 82577 280961 82625 280989
rect 82653 280961 82687 280989
rect 82715 280961 82749 280989
rect 82777 280961 82811 280989
rect 82839 280961 82887 280989
rect 82577 272175 82887 280961
rect 82577 272147 82625 272175
rect 82653 272147 82687 272175
rect 82715 272147 82749 272175
rect 82777 272147 82811 272175
rect 82839 272147 82887 272175
rect 82577 272113 82887 272147
rect 82577 272085 82625 272113
rect 82653 272085 82687 272113
rect 82715 272085 82749 272113
rect 82777 272085 82811 272113
rect 82839 272085 82887 272113
rect 82577 272051 82887 272085
rect 82577 272023 82625 272051
rect 82653 272023 82687 272051
rect 82715 272023 82749 272051
rect 82777 272023 82811 272051
rect 82839 272023 82887 272051
rect 82577 271989 82887 272023
rect 82577 271961 82625 271989
rect 82653 271961 82687 271989
rect 82715 271961 82749 271989
rect 82777 271961 82811 271989
rect 82839 271961 82887 271989
rect 82577 263175 82887 271961
rect 82577 263147 82625 263175
rect 82653 263147 82687 263175
rect 82715 263147 82749 263175
rect 82777 263147 82811 263175
rect 82839 263147 82887 263175
rect 82577 263113 82887 263147
rect 82577 263085 82625 263113
rect 82653 263085 82687 263113
rect 82715 263085 82749 263113
rect 82777 263085 82811 263113
rect 82839 263085 82887 263113
rect 82577 263051 82887 263085
rect 82577 263023 82625 263051
rect 82653 263023 82687 263051
rect 82715 263023 82749 263051
rect 82777 263023 82811 263051
rect 82839 263023 82887 263051
rect 82577 262989 82887 263023
rect 82577 262961 82625 262989
rect 82653 262961 82687 262989
rect 82715 262961 82749 262989
rect 82777 262961 82811 262989
rect 82839 262961 82887 262989
rect 82577 260603 82887 262961
rect 84437 299086 84747 299134
rect 84437 299058 84485 299086
rect 84513 299058 84547 299086
rect 84575 299058 84609 299086
rect 84637 299058 84671 299086
rect 84699 299058 84747 299086
rect 84437 299024 84747 299058
rect 84437 298996 84485 299024
rect 84513 298996 84547 299024
rect 84575 298996 84609 299024
rect 84637 298996 84671 299024
rect 84699 298996 84747 299024
rect 84437 298962 84747 298996
rect 84437 298934 84485 298962
rect 84513 298934 84547 298962
rect 84575 298934 84609 298962
rect 84637 298934 84671 298962
rect 84699 298934 84747 298962
rect 84437 298900 84747 298934
rect 84437 298872 84485 298900
rect 84513 298872 84547 298900
rect 84575 298872 84609 298900
rect 84637 298872 84671 298900
rect 84699 298872 84747 298900
rect 84437 293175 84747 298872
rect 84437 293147 84485 293175
rect 84513 293147 84547 293175
rect 84575 293147 84609 293175
rect 84637 293147 84671 293175
rect 84699 293147 84747 293175
rect 84437 293113 84747 293147
rect 84437 293085 84485 293113
rect 84513 293085 84547 293113
rect 84575 293085 84609 293113
rect 84637 293085 84671 293113
rect 84699 293085 84747 293113
rect 84437 293051 84747 293085
rect 84437 293023 84485 293051
rect 84513 293023 84547 293051
rect 84575 293023 84609 293051
rect 84637 293023 84671 293051
rect 84699 293023 84747 293051
rect 84437 292989 84747 293023
rect 84437 292961 84485 292989
rect 84513 292961 84547 292989
rect 84575 292961 84609 292989
rect 84637 292961 84671 292989
rect 84699 292961 84747 292989
rect 84437 284175 84747 292961
rect 84437 284147 84485 284175
rect 84513 284147 84547 284175
rect 84575 284147 84609 284175
rect 84637 284147 84671 284175
rect 84699 284147 84747 284175
rect 84437 284113 84747 284147
rect 84437 284085 84485 284113
rect 84513 284085 84547 284113
rect 84575 284085 84609 284113
rect 84637 284085 84671 284113
rect 84699 284085 84747 284113
rect 84437 284051 84747 284085
rect 84437 284023 84485 284051
rect 84513 284023 84547 284051
rect 84575 284023 84609 284051
rect 84637 284023 84671 284051
rect 84699 284023 84747 284051
rect 84437 283989 84747 284023
rect 84437 283961 84485 283989
rect 84513 283961 84547 283989
rect 84575 283961 84609 283989
rect 84637 283961 84671 283989
rect 84699 283961 84747 283989
rect 84437 275175 84747 283961
rect 84437 275147 84485 275175
rect 84513 275147 84547 275175
rect 84575 275147 84609 275175
rect 84637 275147 84671 275175
rect 84699 275147 84747 275175
rect 84437 275113 84747 275147
rect 84437 275085 84485 275113
rect 84513 275085 84547 275113
rect 84575 275085 84609 275113
rect 84637 275085 84671 275113
rect 84699 275085 84747 275113
rect 84437 275051 84747 275085
rect 84437 275023 84485 275051
rect 84513 275023 84547 275051
rect 84575 275023 84609 275051
rect 84637 275023 84671 275051
rect 84699 275023 84747 275051
rect 84437 274989 84747 275023
rect 84437 274961 84485 274989
rect 84513 274961 84547 274989
rect 84575 274961 84609 274989
rect 84637 274961 84671 274989
rect 84699 274961 84747 274989
rect 84437 266175 84747 274961
rect 84437 266147 84485 266175
rect 84513 266147 84547 266175
rect 84575 266147 84609 266175
rect 84637 266147 84671 266175
rect 84699 266147 84747 266175
rect 84437 266113 84747 266147
rect 84437 266085 84485 266113
rect 84513 266085 84547 266113
rect 84575 266085 84609 266113
rect 84637 266085 84671 266113
rect 84699 266085 84747 266113
rect 84437 266051 84747 266085
rect 84437 266023 84485 266051
rect 84513 266023 84547 266051
rect 84575 266023 84609 266051
rect 84637 266023 84671 266051
rect 84699 266023 84747 266051
rect 84437 265989 84747 266023
rect 84437 265961 84485 265989
rect 84513 265961 84547 265989
rect 84575 265961 84609 265989
rect 84637 265961 84671 265989
rect 84699 265961 84747 265989
rect 84437 260603 84747 265961
rect 91577 298606 91887 299134
rect 91577 298578 91625 298606
rect 91653 298578 91687 298606
rect 91715 298578 91749 298606
rect 91777 298578 91811 298606
rect 91839 298578 91887 298606
rect 91577 298544 91887 298578
rect 91577 298516 91625 298544
rect 91653 298516 91687 298544
rect 91715 298516 91749 298544
rect 91777 298516 91811 298544
rect 91839 298516 91887 298544
rect 91577 298482 91887 298516
rect 91577 298454 91625 298482
rect 91653 298454 91687 298482
rect 91715 298454 91749 298482
rect 91777 298454 91811 298482
rect 91839 298454 91887 298482
rect 91577 298420 91887 298454
rect 91577 298392 91625 298420
rect 91653 298392 91687 298420
rect 91715 298392 91749 298420
rect 91777 298392 91811 298420
rect 91839 298392 91887 298420
rect 91577 290175 91887 298392
rect 91577 290147 91625 290175
rect 91653 290147 91687 290175
rect 91715 290147 91749 290175
rect 91777 290147 91811 290175
rect 91839 290147 91887 290175
rect 91577 290113 91887 290147
rect 91577 290085 91625 290113
rect 91653 290085 91687 290113
rect 91715 290085 91749 290113
rect 91777 290085 91811 290113
rect 91839 290085 91887 290113
rect 91577 290051 91887 290085
rect 91577 290023 91625 290051
rect 91653 290023 91687 290051
rect 91715 290023 91749 290051
rect 91777 290023 91811 290051
rect 91839 290023 91887 290051
rect 91577 289989 91887 290023
rect 91577 289961 91625 289989
rect 91653 289961 91687 289989
rect 91715 289961 91749 289989
rect 91777 289961 91811 289989
rect 91839 289961 91887 289989
rect 91577 281175 91887 289961
rect 91577 281147 91625 281175
rect 91653 281147 91687 281175
rect 91715 281147 91749 281175
rect 91777 281147 91811 281175
rect 91839 281147 91887 281175
rect 91577 281113 91887 281147
rect 91577 281085 91625 281113
rect 91653 281085 91687 281113
rect 91715 281085 91749 281113
rect 91777 281085 91811 281113
rect 91839 281085 91887 281113
rect 91577 281051 91887 281085
rect 91577 281023 91625 281051
rect 91653 281023 91687 281051
rect 91715 281023 91749 281051
rect 91777 281023 91811 281051
rect 91839 281023 91887 281051
rect 91577 280989 91887 281023
rect 91577 280961 91625 280989
rect 91653 280961 91687 280989
rect 91715 280961 91749 280989
rect 91777 280961 91811 280989
rect 91839 280961 91887 280989
rect 91577 272175 91887 280961
rect 91577 272147 91625 272175
rect 91653 272147 91687 272175
rect 91715 272147 91749 272175
rect 91777 272147 91811 272175
rect 91839 272147 91887 272175
rect 91577 272113 91887 272147
rect 91577 272085 91625 272113
rect 91653 272085 91687 272113
rect 91715 272085 91749 272113
rect 91777 272085 91811 272113
rect 91839 272085 91887 272113
rect 91577 272051 91887 272085
rect 91577 272023 91625 272051
rect 91653 272023 91687 272051
rect 91715 272023 91749 272051
rect 91777 272023 91811 272051
rect 91839 272023 91887 272051
rect 91577 271989 91887 272023
rect 91577 271961 91625 271989
rect 91653 271961 91687 271989
rect 91715 271961 91749 271989
rect 91777 271961 91811 271989
rect 91839 271961 91887 271989
rect 91577 263175 91887 271961
rect 91577 263147 91625 263175
rect 91653 263147 91687 263175
rect 91715 263147 91749 263175
rect 91777 263147 91811 263175
rect 91839 263147 91887 263175
rect 91577 263113 91887 263147
rect 91577 263085 91625 263113
rect 91653 263085 91687 263113
rect 91715 263085 91749 263113
rect 91777 263085 91811 263113
rect 91839 263085 91887 263113
rect 91577 263051 91887 263085
rect 91577 263023 91625 263051
rect 91653 263023 91687 263051
rect 91715 263023 91749 263051
rect 91777 263023 91811 263051
rect 91839 263023 91887 263051
rect 91577 262989 91887 263023
rect 91577 262961 91625 262989
rect 91653 262961 91687 262989
rect 91715 262961 91749 262989
rect 91777 262961 91811 262989
rect 91839 262961 91887 262989
rect 91577 260603 91887 262961
rect 93437 299086 93747 299134
rect 93437 299058 93485 299086
rect 93513 299058 93547 299086
rect 93575 299058 93609 299086
rect 93637 299058 93671 299086
rect 93699 299058 93747 299086
rect 93437 299024 93747 299058
rect 93437 298996 93485 299024
rect 93513 298996 93547 299024
rect 93575 298996 93609 299024
rect 93637 298996 93671 299024
rect 93699 298996 93747 299024
rect 93437 298962 93747 298996
rect 93437 298934 93485 298962
rect 93513 298934 93547 298962
rect 93575 298934 93609 298962
rect 93637 298934 93671 298962
rect 93699 298934 93747 298962
rect 93437 298900 93747 298934
rect 93437 298872 93485 298900
rect 93513 298872 93547 298900
rect 93575 298872 93609 298900
rect 93637 298872 93671 298900
rect 93699 298872 93747 298900
rect 93437 293175 93747 298872
rect 93437 293147 93485 293175
rect 93513 293147 93547 293175
rect 93575 293147 93609 293175
rect 93637 293147 93671 293175
rect 93699 293147 93747 293175
rect 93437 293113 93747 293147
rect 93437 293085 93485 293113
rect 93513 293085 93547 293113
rect 93575 293085 93609 293113
rect 93637 293085 93671 293113
rect 93699 293085 93747 293113
rect 93437 293051 93747 293085
rect 93437 293023 93485 293051
rect 93513 293023 93547 293051
rect 93575 293023 93609 293051
rect 93637 293023 93671 293051
rect 93699 293023 93747 293051
rect 93437 292989 93747 293023
rect 93437 292961 93485 292989
rect 93513 292961 93547 292989
rect 93575 292961 93609 292989
rect 93637 292961 93671 292989
rect 93699 292961 93747 292989
rect 93437 284175 93747 292961
rect 93437 284147 93485 284175
rect 93513 284147 93547 284175
rect 93575 284147 93609 284175
rect 93637 284147 93671 284175
rect 93699 284147 93747 284175
rect 93437 284113 93747 284147
rect 93437 284085 93485 284113
rect 93513 284085 93547 284113
rect 93575 284085 93609 284113
rect 93637 284085 93671 284113
rect 93699 284085 93747 284113
rect 93437 284051 93747 284085
rect 93437 284023 93485 284051
rect 93513 284023 93547 284051
rect 93575 284023 93609 284051
rect 93637 284023 93671 284051
rect 93699 284023 93747 284051
rect 93437 283989 93747 284023
rect 93437 283961 93485 283989
rect 93513 283961 93547 283989
rect 93575 283961 93609 283989
rect 93637 283961 93671 283989
rect 93699 283961 93747 283989
rect 93437 275175 93747 283961
rect 93437 275147 93485 275175
rect 93513 275147 93547 275175
rect 93575 275147 93609 275175
rect 93637 275147 93671 275175
rect 93699 275147 93747 275175
rect 93437 275113 93747 275147
rect 93437 275085 93485 275113
rect 93513 275085 93547 275113
rect 93575 275085 93609 275113
rect 93637 275085 93671 275113
rect 93699 275085 93747 275113
rect 93437 275051 93747 275085
rect 93437 275023 93485 275051
rect 93513 275023 93547 275051
rect 93575 275023 93609 275051
rect 93637 275023 93671 275051
rect 93699 275023 93747 275051
rect 93437 274989 93747 275023
rect 93437 274961 93485 274989
rect 93513 274961 93547 274989
rect 93575 274961 93609 274989
rect 93637 274961 93671 274989
rect 93699 274961 93747 274989
rect 93437 266175 93747 274961
rect 93437 266147 93485 266175
rect 93513 266147 93547 266175
rect 93575 266147 93609 266175
rect 93637 266147 93671 266175
rect 93699 266147 93747 266175
rect 93437 266113 93747 266147
rect 93437 266085 93485 266113
rect 93513 266085 93547 266113
rect 93575 266085 93609 266113
rect 93637 266085 93671 266113
rect 93699 266085 93747 266113
rect 93437 266051 93747 266085
rect 93437 266023 93485 266051
rect 93513 266023 93547 266051
rect 93575 266023 93609 266051
rect 93637 266023 93671 266051
rect 93699 266023 93747 266051
rect 93437 265989 93747 266023
rect 93437 265961 93485 265989
rect 93513 265961 93547 265989
rect 93575 265961 93609 265989
rect 93637 265961 93671 265989
rect 93699 265961 93747 265989
rect 93437 260603 93747 265961
rect 100577 298606 100887 299134
rect 100577 298578 100625 298606
rect 100653 298578 100687 298606
rect 100715 298578 100749 298606
rect 100777 298578 100811 298606
rect 100839 298578 100887 298606
rect 100577 298544 100887 298578
rect 100577 298516 100625 298544
rect 100653 298516 100687 298544
rect 100715 298516 100749 298544
rect 100777 298516 100811 298544
rect 100839 298516 100887 298544
rect 100577 298482 100887 298516
rect 100577 298454 100625 298482
rect 100653 298454 100687 298482
rect 100715 298454 100749 298482
rect 100777 298454 100811 298482
rect 100839 298454 100887 298482
rect 100577 298420 100887 298454
rect 100577 298392 100625 298420
rect 100653 298392 100687 298420
rect 100715 298392 100749 298420
rect 100777 298392 100811 298420
rect 100839 298392 100887 298420
rect 100577 290175 100887 298392
rect 100577 290147 100625 290175
rect 100653 290147 100687 290175
rect 100715 290147 100749 290175
rect 100777 290147 100811 290175
rect 100839 290147 100887 290175
rect 100577 290113 100887 290147
rect 100577 290085 100625 290113
rect 100653 290085 100687 290113
rect 100715 290085 100749 290113
rect 100777 290085 100811 290113
rect 100839 290085 100887 290113
rect 100577 290051 100887 290085
rect 100577 290023 100625 290051
rect 100653 290023 100687 290051
rect 100715 290023 100749 290051
rect 100777 290023 100811 290051
rect 100839 290023 100887 290051
rect 100577 289989 100887 290023
rect 100577 289961 100625 289989
rect 100653 289961 100687 289989
rect 100715 289961 100749 289989
rect 100777 289961 100811 289989
rect 100839 289961 100887 289989
rect 100577 281175 100887 289961
rect 100577 281147 100625 281175
rect 100653 281147 100687 281175
rect 100715 281147 100749 281175
rect 100777 281147 100811 281175
rect 100839 281147 100887 281175
rect 100577 281113 100887 281147
rect 100577 281085 100625 281113
rect 100653 281085 100687 281113
rect 100715 281085 100749 281113
rect 100777 281085 100811 281113
rect 100839 281085 100887 281113
rect 100577 281051 100887 281085
rect 100577 281023 100625 281051
rect 100653 281023 100687 281051
rect 100715 281023 100749 281051
rect 100777 281023 100811 281051
rect 100839 281023 100887 281051
rect 100577 280989 100887 281023
rect 100577 280961 100625 280989
rect 100653 280961 100687 280989
rect 100715 280961 100749 280989
rect 100777 280961 100811 280989
rect 100839 280961 100887 280989
rect 100577 272175 100887 280961
rect 100577 272147 100625 272175
rect 100653 272147 100687 272175
rect 100715 272147 100749 272175
rect 100777 272147 100811 272175
rect 100839 272147 100887 272175
rect 100577 272113 100887 272147
rect 100577 272085 100625 272113
rect 100653 272085 100687 272113
rect 100715 272085 100749 272113
rect 100777 272085 100811 272113
rect 100839 272085 100887 272113
rect 100577 272051 100887 272085
rect 100577 272023 100625 272051
rect 100653 272023 100687 272051
rect 100715 272023 100749 272051
rect 100777 272023 100811 272051
rect 100839 272023 100887 272051
rect 100577 271989 100887 272023
rect 100577 271961 100625 271989
rect 100653 271961 100687 271989
rect 100715 271961 100749 271989
rect 100777 271961 100811 271989
rect 100839 271961 100887 271989
rect 100577 263175 100887 271961
rect 100577 263147 100625 263175
rect 100653 263147 100687 263175
rect 100715 263147 100749 263175
rect 100777 263147 100811 263175
rect 100839 263147 100887 263175
rect 100577 263113 100887 263147
rect 100577 263085 100625 263113
rect 100653 263085 100687 263113
rect 100715 263085 100749 263113
rect 100777 263085 100811 263113
rect 100839 263085 100887 263113
rect 100577 263051 100887 263085
rect 100577 263023 100625 263051
rect 100653 263023 100687 263051
rect 100715 263023 100749 263051
rect 100777 263023 100811 263051
rect 100839 263023 100887 263051
rect 100577 262989 100887 263023
rect 100577 262961 100625 262989
rect 100653 262961 100687 262989
rect 100715 262961 100749 262989
rect 100777 262961 100811 262989
rect 100839 262961 100887 262989
rect 100577 260603 100887 262961
rect 102437 299086 102747 299134
rect 102437 299058 102485 299086
rect 102513 299058 102547 299086
rect 102575 299058 102609 299086
rect 102637 299058 102671 299086
rect 102699 299058 102747 299086
rect 102437 299024 102747 299058
rect 102437 298996 102485 299024
rect 102513 298996 102547 299024
rect 102575 298996 102609 299024
rect 102637 298996 102671 299024
rect 102699 298996 102747 299024
rect 102437 298962 102747 298996
rect 102437 298934 102485 298962
rect 102513 298934 102547 298962
rect 102575 298934 102609 298962
rect 102637 298934 102671 298962
rect 102699 298934 102747 298962
rect 102437 298900 102747 298934
rect 102437 298872 102485 298900
rect 102513 298872 102547 298900
rect 102575 298872 102609 298900
rect 102637 298872 102671 298900
rect 102699 298872 102747 298900
rect 102437 293175 102747 298872
rect 102437 293147 102485 293175
rect 102513 293147 102547 293175
rect 102575 293147 102609 293175
rect 102637 293147 102671 293175
rect 102699 293147 102747 293175
rect 102437 293113 102747 293147
rect 102437 293085 102485 293113
rect 102513 293085 102547 293113
rect 102575 293085 102609 293113
rect 102637 293085 102671 293113
rect 102699 293085 102747 293113
rect 102437 293051 102747 293085
rect 102437 293023 102485 293051
rect 102513 293023 102547 293051
rect 102575 293023 102609 293051
rect 102637 293023 102671 293051
rect 102699 293023 102747 293051
rect 102437 292989 102747 293023
rect 102437 292961 102485 292989
rect 102513 292961 102547 292989
rect 102575 292961 102609 292989
rect 102637 292961 102671 292989
rect 102699 292961 102747 292989
rect 102437 284175 102747 292961
rect 102437 284147 102485 284175
rect 102513 284147 102547 284175
rect 102575 284147 102609 284175
rect 102637 284147 102671 284175
rect 102699 284147 102747 284175
rect 102437 284113 102747 284147
rect 102437 284085 102485 284113
rect 102513 284085 102547 284113
rect 102575 284085 102609 284113
rect 102637 284085 102671 284113
rect 102699 284085 102747 284113
rect 102437 284051 102747 284085
rect 102437 284023 102485 284051
rect 102513 284023 102547 284051
rect 102575 284023 102609 284051
rect 102637 284023 102671 284051
rect 102699 284023 102747 284051
rect 102437 283989 102747 284023
rect 102437 283961 102485 283989
rect 102513 283961 102547 283989
rect 102575 283961 102609 283989
rect 102637 283961 102671 283989
rect 102699 283961 102747 283989
rect 102437 275175 102747 283961
rect 102437 275147 102485 275175
rect 102513 275147 102547 275175
rect 102575 275147 102609 275175
rect 102637 275147 102671 275175
rect 102699 275147 102747 275175
rect 102437 275113 102747 275147
rect 102437 275085 102485 275113
rect 102513 275085 102547 275113
rect 102575 275085 102609 275113
rect 102637 275085 102671 275113
rect 102699 275085 102747 275113
rect 102437 275051 102747 275085
rect 102437 275023 102485 275051
rect 102513 275023 102547 275051
rect 102575 275023 102609 275051
rect 102637 275023 102671 275051
rect 102699 275023 102747 275051
rect 102437 274989 102747 275023
rect 102437 274961 102485 274989
rect 102513 274961 102547 274989
rect 102575 274961 102609 274989
rect 102637 274961 102671 274989
rect 102699 274961 102747 274989
rect 102437 266175 102747 274961
rect 102437 266147 102485 266175
rect 102513 266147 102547 266175
rect 102575 266147 102609 266175
rect 102637 266147 102671 266175
rect 102699 266147 102747 266175
rect 102437 266113 102747 266147
rect 102437 266085 102485 266113
rect 102513 266085 102547 266113
rect 102575 266085 102609 266113
rect 102637 266085 102671 266113
rect 102699 266085 102747 266113
rect 102437 266051 102747 266085
rect 102437 266023 102485 266051
rect 102513 266023 102547 266051
rect 102575 266023 102609 266051
rect 102637 266023 102671 266051
rect 102699 266023 102747 266051
rect 102437 265989 102747 266023
rect 102437 265961 102485 265989
rect 102513 265961 102547 265989
rect 102575 265961 102609 265989
rect 102637 265961 102671 265989
rect 102699 265961 102747 265989
rect 102437 260603 102747 265961
rect 109577 298606 109887 299134
rect 109577 298578 109625 298606
rect 109653 298578 109687 298606
rect 109715 298578 109749 298606
rect 109777 298578 109811 298606
rect 109839 298578 109887 298606
rect 109577 298544 109887 298578
rect 109577 298516 109625 298544
rect 109653 298516 109687 298544
rect 109715 298516 109749 298544
rect 109777 298516 109811 298544
rect 109839 298516 109887 298544
rect 109577 298482 109887 298516
rect 109577 298454 109625 298482
rect 109653 298454 109687 298482
rect 109715 298454 109749 298482
rect 109777 298454 109811 298482
rect 109839 298454 109887 298482
rect 109577 298420 109887 298454
rect 109577 298392 109625 298420
rect 109653 298392 109687 298420
rect 109715 298392 109749 298420
rect 109777 298392 109811 298420
rect 109839 298392 109887 298420
rect 109577 290175 109887 298392
rect 109577 290147 109625 290175
rect 109653 290147 109687 290175
rect 109715 290147 109749 290175
rect 109777 290147 109811 290175
rect 109839 290147 109887 290175
rect 109577 290113 109887 290147
rect 109577 290085 109625 290113
rect 109653 290085 109687 290113
rect 109715 290085 109749 290113
rect 109777 290085 109811 290113
rect 109839 290085 109887 290113
rect 109577 290051 109887 290085
rect 109577 290023 109625 290051
rect 109653 290023 109687 290051
rect 109715 290023 109749 290051
rect 109777 290023 109811 290051
rect 109839 290023 109887 290051
rect 109577 289989 109887 290023
rect 109577 289961 109625 289989
rect 109653 289961 109687 289989
rect 109715 289961 109749 289989
rect 109777 289961 109811 289989
rect 109839 289961 109887 289989
rect 109577 281175 109887 289961
rect 109577 281147 109625 281175
rect 109653 281147 109687 281175
rect 109715 281147 109749 281175
rect 109777 281147 109811 281175
rect 109839 281147 109887 281175
rect 109577 281113 109887 281147
rect 109577 281085 109625 281113
rect 109653 281085 109687 281113
rect 109715 281085 109749 281113
rect 109777 281085 109811 281113
rect 109839 281085 109887 281113
rect 109577 281051 109887 281085
rect 109577 281023 109625 281051
rect 109653 281023 109687 281051
rect 109715 281023 109749 281051
rect 109777 281023 109811 281051
rect 109839 281023 109887 281051
rect 109577 280989 109887 281023
rect 109577 280961 109625 280989
rect 109653 280961 109687 280989
rect 109715 280961 109749 280989
rect 109777 280961 109811 280989
rect 109839 280961 109887 280989
rect 109577 272175 109887 280961
rect 109577 272147 109625 272175
rect 109653 272147 109687 272175
rect 109715 272147 109749 272175
rect 109777 272147 109811 272175
rect 109839 272147 109887 272175
rect 109577 272113 109887 272147
rect 109577 272085 109625 272113
rect 109653 272085 109687 272113
rect 109715 272085 109749 272113
rect 109777 272085 109811 272113
rect 109839 272085 109887 272113
rect 109577 272051 109887 272085
rect 109577 272023 109625 272051
rect 109653 272023 109687 272051
rect 109715 272023 109749 272051
rect 109777 272023 109811 272051
rect 109839 272023 109887 272051
rect 109577 271989 109887 272023
rect 109577 271961 109625 271989
rect 109653 271961 109687 271989
rect 109715 271961 109749 271989
rect 109777 271961 109811 271989
rect 109839 271961 109887 271989
rect 109577 263175 109887 271961
rect 109577 263147 109625 263175
rect 109653 263147 109687 263175
rect 109715 263147 109749 263175
rect 109777 263147 109811 263175
rect 109839 263147 109887 263175
rect 109577 263113 109887 263147
rect 109577 263085 109625 263113
rect 109653 263085 109687 263113
rect 109715 263085 109749 263113
rect 109777 263085 109811 263113
rect 109839 263085 109887 263113
rect 109577 263051 109887 263085
rect 109577 263023 109625 263051
rect 109653 263023 109687 263051
rect 109715 263023 109749 263051
rect 109777 263023 109811 263051
rect 109839 263023 109887 263051
rect 109577 262989 109887 263023
rect 109577 262961 109625 262989
rect 109653 262961 109687 262989
rect 109715 262961 109749 262989
rect 109777 262961 109811 262989
rect 109839 262961 109887 262989
rect 109577 260603 109887 262961
rect 111437 299086 111747 299134
rect 111437 299058 111485 299086
rect 111513 299058 111547 299086
rect 111575 299058 111609 299086
rect 111637 299058 111671 299086
rect 111699 299058 111747 299086
rect 111437 299024 111747 299058
rect 111437 298996 111485 299024
rect 111513 298996 111547 299024
rect 111575 298996 111609 299024
rect 111637 298996 111671 299024
rect 111699 298996 111747 299024
rect 111437 298962 111747 298996
rect 111437 298934 111485 298962
rect 111513 298934 111547 298962
rect 111575 298934 111609 298962
rect 111637 298934 111671 298962
rect 111699 298934 111747 298962
rect 111437 298900 111747 298934
rect 111437 298872 111485 298900
rect 111513 298872 111547 298900
rect 111575 298872 111609 298900
rect 111637 298872 111671 298900
rect 111699 298872 111747 298900
rect 111437 293175 111747 298872
rect 111437 293147 111485 293175
rect 111513 293147 111547 293175
rect 111575 293147 111609 293175
rect 111637 293147 111671 293175
rect 111699 293147 111747 293175
rect 111437 293113 111747 293147
rect 111437 293085 111485 293113
rect 111513 293085 111547 293113
rect 111575 293085 111609 293113
rect 111637 293085 111671 293113
rect 111699 293085 111747 293113
rect 111437 293051 111747 293085
rect 111437 293023 111485 293051
rect 111513 293023 111547 293051
rect 111575 293023 111609 293051
rect 111637 293023 111671 293051
rect 111699 293023 111747 293051
rect 111437 292989 111747 293023
rect 111437 292961 111485 292989
rect 111513 292961 111547 292989
rect 111575 292961 111609 292989
rect 111637 292961 111671 292989
rect 111699 292961 111747 292989
rect 111437 284175 111747 292961
rect 111437 284147 111485 284175
rect 111513 284147 111547 284175
rect 111575 284147 111609 284175
rect 111637 284147 111671 284175
rect 111699 284147 111747 284175
rect 111437 284113 111747 284147
rect 111437 284085 111485 284113
rect 111513 284085 111547 284113
rect 111575 284085 111609 284113
rect 111637 284085 111671 284113
rect 111699 284085 111747 284113
rect 111437 284051 111747 284085
rect 111437 284023 111485 284051
rect 111513 284023 111547 284051
rect 111575 284023 111609 284051
rect 111637 284023 111671 284051
rect 111699 284023 111747 284051
rect 111437 283989 111747 284023
rect 111437 283961 111485 283989
rect 111513 283961 111547 283989
rect 111575 283961 111609 283989
rect 111637 283961 111671 283989
rect 111699 283961 111747 283989
rect 111437 275175 111747 283961
rect 111437 275147 111485 275175
rect 111513 275147 111547 275175
rect 111575 275147 111609 275175
rect 111637 275147 111671 275175
rect 111699 275147 111747 275175
rect 111437 275113 111747 275147
rect 111437 275085 111485 275113
rect 111513 275085 111547 275113
rect 111575 275085 111609 275113
rect 111637 275085 111671 275113
rect 111699 275085 111747 275113
rect 111437 275051 111747 275085
rect 111437 275023 111485 275051
rect 111513 275023 111547 275051
rect 111575 275023 111609 275051
rect 111637 275023 111671 275051
rect 111699 275023 111747 275051
rect 111437 274989 111747 275023
rect 111437 274961 111485 274989
rect 111513 274961 111547 274989
rect 111575 274961 111609 274989
rect 111637 274961 111671 274989
rect 111699 274961 111747 274989
rect 111437 266175 111747 274961
rect 111437 266147 111485 266175
rect 111513 266147 111547 266175
rect 111575 266147 111609 266175
rect 111637 266147 111671 266175
rect 111699 266147 111747 266175
rect 111437 266113 111747 266147
rect 111437 266085 111485 266113
rect 111513 266085 111547 266113
rect 111575 266085 111609 266113
rect 111637 266085 111671 266113
rect 111699 266085 111747 266113
rect 111437 266051 111747 266085
rect 111437 266023 111485 266051
rect 111513 266023 111547 266051
rect 111575 266023 111609 266051
rect 111637 266023 111671 266051
rect 111699 266023 111747 266051
rect 111437 265989 111747 266023
rect 111437 265961 111485 265989
rect 111513 265961 111547 265989
rect 111575 265961 111609 265989
rect 111637 265961 111671 265989
rect 111699 265961 111747 265989
rect 111437 260603 111747 265961
rect 118577 298606 118887 299134
rect 118577 298578 118625 298606
rect 118653 298578 118687 298606
rect 118715 298578 118749 298606
rect 118777 298578 118811 298606
rect 118839 298578 118887 298606
rect 118577 298544 118887 298578
rect 118577 298516 118625 298544
rect 118653 298516 118687 298544
rect 118715 298516 118749 298544
rect 118777 298516 118811 298544
rect 118839 298516 118887 298544
rect 118577 298482 118887 298516
rect 118577 298454 118625 298482
rect 118653 298454 118687 298482
rect 118715 298454 118749 298482
rect 118777 298454 118811 298482
rect 118839 298454 118887 298482
rect 118577 298420 118887 298454
rect 118577 298392 118625 298420
rect 118653 298392 118687 298420
rect 118715 298392 118749 298420
rect 118777 298392 118811 298420
rect 118839 298392 118887 298420
rect 118577 290175 118887 298392
rect 118577 290147 118625 290175
rect 118653 290147 118687 290175
rect 118715 290147 118749 290175
rect 118777 290147 118811 290175
rect 118839 290147 118887 290175
rect 118577 290113 118887 290147
rect 118577 290085 118625 290113
rect 118653 290085 118687 290113
rect 118715 290085 118749 290113
rect 118777 290085 118811 290113
rect 118839 290085 118887 290113
rect 118577 290051 118887 290085
rect 118577 290023 118625 290051
rect 118653 290023 118687 290051
rect 118715 290023 118749 290051
rect 118777 290023 118811 290051
rect 118839 290023 118887 290051
rect 118577 289989 118887 290023
rect 118577 289961 118625 289989
rect 118653 289961 118687 289989
rect 118715 289961 118749 289989
rect 118777 289961 118811 289989
rect 118839 289961 118887 289989
rect 118577 281175 118887 289961
rect 118577 281147 118625 281175
rect 118653 281147 118687 281175
rect 118715 281147 118749 281175
rect 118777 281147 118811 281175
rect 118839 281147 118887 281175
rect 118577 281113 118887 281147
rect 118577 281085 118625 281113
rect 118653 281085 118687 281113
rect 118715 281085 118749 281113
rect 118777 281085 118811 281113
rect 118839 281085 118887 281113
rect 118577 281051 118887 281085
rect 118577 281023 118625 281051
rect 118653 281023 118687 281051
rect 118715 281023 118749 281051
rect 118777 281023 118811 281051
rect 118839 281023 118887 281051
rect 118577 280989 118887 281023
rect 118577 280961 118625 280989
rect 118653 280961 118687 280989
rect 118715 280961 118749 280989
rect 118777 280961 118811 280989
rect 118839 280961 118887 280989
rect 118577 272175 118887 280961
rect 118577 272147 118625 272175
rect 118653 272147 118687 272175
rect 118715 272147 118749 272175
rect 118777 272147 118811 272175
rect 118839 272147 118887 272175
rect 118577 272113 118887 272147
rect 118577 272085 118625 272113
rect 118653 272085 118687 272113
rect 118715 272085 118749 272113
rect 118777 272085 118811 272113
rect 118839 272085 118887 272113
rect 118577 272051 118887 272085
rect 118577 272023 118625 272051
rect 118653 272023 118687 272051
rect 118715 272023 118749 272051
rect 118777 272023 118811 272051
rect 118839 272023 118887 272051
rect 118577 271989 118887 272023
rect 118577 271961 118625 271989
rect 118653 271961 118687 271989
rect 118715 271961 118749 271989
rect 118777 271961 118811 271989
rect 118839 271961 118887 271989
rect 118577 263175 118887 271961
rect 118577 263147 118625 263175
rect 118653 263147 118687 263175
rect 118715 263147 118749 263175
rect 118777 263147 118811 263175
rect 118839 263147 118887 263175
rect 118577 263113 118887 263147
rect 118577 263085 118625 263113
rect 118653 263085 118687 263113
rect 118715 263085 118749 263113
rect 118777 263085 118811 263113
rect 118839 263085 118887 263113
rect 118577 263051 118887 263085
rect 118577 263023 118625 263051
rect 118653 263023 118687 263051
rect 118715 263023 118749 263051
rect 118777 263023 118811 263051
rect 118839 263023 118887 263051
rect 118577 262989 118887 263023
rect 118577 262961 118625 262989
rect 118653 262961 118687 262989
rect 118715 262961 118749 262989
rect 118777 262961 118811 262989
rect 118839 262961 118887 262989
rect 118577 260603 118887 262961
rect 120437 299086 120747 299134
rect 120437 299058 120485 299086
rect 120513 299058 120547 299086
rect 120575 299058 120609 299086
rect 120637 299058 120671 299086
rect 120699 299058 120747 299086
rect 120437 299024 120747 299058
rect 120437 298996 120485 299024
rect 120513 298996 120547 299024
rect 120575 298996 120609 299024
rect 120637 298996 120671 299024
rect 120699 298996 120747 299024
rect 120437 298962 120747 298996
rect 120437 298934 120485 298962
rect 120513 298934 120547 298962
rect 120575 298934 120609 298962
rect 120637 298934 120671 298962
rect 120699 298934 120747 298962
rect 120437 298900 120747 298934
rect 120437 298872 120485 298900
rect 120513 298872 120547 298900
rect 120575 298872 120609 298900
rect 120637 298872 120671 298900
rect 120699 298872 120747 298900
rect 120437 293175 120747 298872
rect 120437 293147 120485 293175
rect 120513 293147 120547 293175
rect 120575 293147 120609 293175
rect 120637 293147 120671 293175
rect 120699 293147 120747 293175
rect 120437 293113 120747 293147
rect 120437 293085 120485 293113
rect 120513 293085 120547 293113
rect 120575 293085 120609 293113
rect 120637 293085 120671 293113
rect 120699 293085 120747 293113
rect 120437 293051 120747 293085
rect 120437 293023 120485 293051
rect 120513 293023 120547 293051
rect 120575 293023 120609 293051
rect 120637 293023 120671 293051
rect 120699 293023 120747 293051
rect 120437 292989 120747 293023
rect 120437 292961 120485 292989
rect 120513 292961 120547 292989
rect 120575 292961 120609 292989
rect 120637 292961 120671 292989
rect 120699 292961 120747 292989
rect 120437 284175 120747 292961
rect 120437 284147 120485 284175
rect 120513 284147 120547 284175
rect 120575 284147 120609 284175
rect 120637 284147 120671 284175
rect 120699 284147 120747 284175
rect 120437 284113 120747 284147
rect 120437 284085 120485 284113
rect 120513 284085 120547 284113
rect 120575 284085 120609 284113
rect 120637 284085 120671 284113
rect 120699 284085 120747 284113
rect 120437 284051 120747 284085
rect 120437 284023 120485 284051
rect 120513 284023 120547 284051
rect 120575 284023 120609 284051
rect 120637 284023 120671 284051
rect 120699 284023 120747 284051
rect 120437 283989 120747 284023
rect 120437 283961 120485 283989
rect 120513 283961 120547 283989
rect 120575 283961 120609 283989
rect 120637 283961 120671 283989
rect 120699 283961 120747 283989
rect 120437 275175 120747 283961
rect 120437 275147 120485 275175
rect 120513 275147 120547 275175
rect 120575 275147 120609 275175
rect 120637 275147 120671 275175
rect 120699 275147 120747 275175
rect 120437 275113 120747 275147
rect 120437 275085 120485 275113
rect 120513 275085 120547 275113
rect 120575 275085 120609 275113
rect 120637 275085 120671 275113
rect 120699 275085 120747 275113
rect 120437 275051 120747 275085
rect 120437 275023 120485 275051
rect 120513 275023 120547 275051
rect 120575 275023 120609 275051
rect 120637 275023 120671 275051
rect 120699 275023 120747 275051
rect 120437 274989 120747 275023
rect 120437 274961 120485 274989
rect 120513 274961 120547 274989
rect 120575 274961 120609 274989
rect 120637 274961 120671 274989
rect 120699 274961 120747 274989
rect 120437 266175 120747 274961
rect 120437 266147 120485 266175
rect 120513 266147 120547 266175
rect 120575 266147 120609 266175
rect 120637 266147 120671 266175
rect 120699 266147 120747 266175
rect 120437 266113 120747 266147
rect 120437 266085 120485 266113
rect 120513 266085 120547 266113
rect 120575 266085 120609 266113
rect 120637 266085 120671 266113
rect 120699 266085 120747 266113
rect 120437 266051 120747 266085
rect 120437 266023 120485 266051
rect 120513 266023 120547 266051
rect 120575 266023 120609 266051
rect 120637 266023 120671 266051
rect 120699 266023 120747 266051
rect 120437 265989 120747 266023
rect 120437 265961 120485 265989
rect 120513 265961 120547 265989
rect 120575 265961 120609 265989
rect 120637 265961 120671 265989
rect 120699 265961 120747 265989
rect 120437 260603 120747 265961
rect 127577 298606 127887 299134
rect 127577 298578 127625 298606
rect 127653 298578 127687 298606
rect 127715 298578 127749 298606
rect 127777 298578 127811 298606
rect 127839 298578 127887 298606
rect 127577 298544 127887 298578
rect 127577 298516 127625 298544
rect 127653 298516 127687 298544
rect 127715 298516 127749 298544
rect 127777 298516 127811 298544
rect 127839 298516 127887 298544
rect 127577 298482 127887 298516
rect 127577 298454 127625 298482
rect 127653 298454 127687 298482
rect 127715 298454 127749 298482
rect 127777 298454 127811 298482
rect 127839 298454 127887 298482
rect 127577 298420 127887 298454
rect 127577 298392 127625 298420
rect 127653 298392 127687 298420
rect 127715 298392 127749 298420
rect 127777 298392 127811 298420
rect 127839 298392 127887 298420
rect 127577 290175 127887 298392
rect 127577 290147 127625 290175
rect 127653 290147 127687 290175
rect 127715 290147 127749 290175
rect 127777 290147 127811 290175
rect 127839 290147 127887 290175
rect 127577 290113 127887 290147
rect 127577 290085 127625 290113
rect 127653 290085 127687 290113
rect 127715 290085 127749 290113
rect 127777 290085 127811 290113
rect 127839 290085 127887 290113
rect 127577 290051 127887 290085
rect 127577 290023 127625 290051
rect 127653 290023 127687 290051
rect 127715 290023 127749 290051
rect 127777 290023 127811 290051
rect 127839 290023 127887 290051
rect 127577 289989 127887 290023
rect 127577 289961 127625 289989
rect 127653 289961 127687 289989
rect 127715 289961 127749 289989
rect 127777 289961 127811 289989
rect 127839 289961 127887 289989
rect 127577 281175 127887 289961
rect 127577 281147 127625 281175
rect 127653 281147 127687 281175
rect 127715 281147 127749 281175
rect 127777 281147 127811 281175
rect 127839 281147 127887 281175
rect 127577 281113 127887 281147
rect 127577 281085 127625 281113
rect 127653 281085 127687 281113
rect 127715 281085 127749 281113
rect 127777 281085 127811 281113
rect 127839 281085 127887 281113
rect 127577 281051 127887 281085
rect 127577 281023 127625 281051
rect 127653 281023 127687 281051
rect 127715 281023 127749 281051
rect 127777 281023 127811 281051
rect 127839 281023 127887 281051
rect 127577 280989 127887 281023
rect 127577 280961 127625 280989
rect 127653 280961 127687 280989
rect 127715 280961 127749 280989
rect 127777 280961 127811 280989
rect 127839 280961 127887 280989
rect 127577 272175 127887 280961
rect 127577 272147 127625 272175
rect 127653 272147 127687 272175
rect 127715 272147 127749 272175
rect 127777 272147 127811 272175
rect 127839 272147 127887 272175
rect 127577 272113 127887 272147
rect 127577 272085 127625 272113
rect 127653 272085 127687 272113
rect 127715 272085 127749 272113
rect 127777 272085 127811 272113
rect 127839 272085 127887 272113
rect 127577 272051 127887 272085
rect 127577 272023 127625 272051
rect 127653 272023 127687 272051
rect 127715 272023 127749 272051
rect 127777 272023 127811 272051
rect 127839 272023 127887 272051
rect 127577 271989 127887 272023
rect 127577 271961 127625 271989
rect 127653 271961 127687 271989
rect 127715 271961 127749 271989
rect 127777 271961 127811 271989
rect 127839 271961 127887 271989
rect 127577 263175 127887 271961
rect 127577 263147 127625 263175
rect 127653 263147 127687 263175
rect 127715 263147 127749 263175
rect 127777 263147 127811 263175
rect 127839 263147 127887 263175
rect 127577 263113 127887 263147
rect 127577 263085 127625 263113
rect 127653 263085 127687 263113
rect 127715 263085 127749 263113
rect 127777 263085 127811 263113
rect 127839 263085 127887 263113
rect 127577 263051 127887 263085
rect 127577 263023 127625 263051
rect 127653 263023 127687 263051
rect 127715 263023 127749 263051
rect 127777 263023 127811 263051
rect 127839 263023 127887 263051
rect 127577 262989 127887 263023
rect 127577 262961 127625 262989
rect 127653 262961 127687 262989
rect 127715 262961 127749 262989
rect 127777 262961 127811 262989
rect 127839 262961 127887 262989
rect 127577 260603 127887 262961
rect 129437 299086 129747 299134
rect 129437 299058 129485 299086
rect 129513 299058 129547 299086
rect 129575 299058 129609 299086
rect 129637 299058 129671 299086
rect 129699 299058 129747 299086
rect 129437 299024 129747 299058
rect 129437 298996 129485 299024
rect 129513 298996 129547 299024
rect 129575 298996 129609 299024
rect 129637 298996 129671 299024
rect 129699 298996 129747 299024
rect 129437 298962 129747 298996
rect 129437 298934 129485 298962
rect 129513 298934 129547 298962
rect 129575 298934 129609 298962
rect 129637 298934 129671 298962
rect 129699 298934 129747 298962
rect 129437 298900 129747 298934
rect 129437 298872 129485 298900
rect 129513 298872 129547 298900
rect 129575 298872 129609 298900
rect 129637 298872 129671 298900
rect 129699 298872 129747 298900
rect 129437 293175 129747 298872
rect 129437 293147 129485 293175
rect 129513 293147 129547 293175
rect 129575 293147 129609 293175
rect 129637 293147 129671 293175
rect 129699 293147 129747 293175
rect 129437 293113 129747 293147
rect 129437 293085 129485 293113
rect 129513 293085 129547 293113
rect 129575 293085 129609 293113
rect 129637 293085 129671 293113
rect 129699 293085 129747 293113
rect 129437 293051 129747 293085
rect 129437 293023 129485 293051
rect 129513 293023 129547 293051
rect 129575 293023 129609 293051
rect 129637 293023 129671 293051
rect 129699 293023 129747 293051
rect 129437 292989 129747 293023
rect 129437 292961 129485 292989
rect 129513 292961 129547 292989
rect 129575 292961 129609 292989
rect 129637 292961 129671 292989
rect 129699 292961 129747 292989
rect 129437 284175 129747 292961
rect 129437 284147 129485 284175
rect 129513 284147 129547 284175
rect 129575 284147 129609 284175
rect 129637 284147 129671 284175
rect 129699 284147 129747 284175
rect 129437 284113 129747 284147
rect 129437 284085 129485 284113
rect 129513 284085 129547 284113
rect 129575 284085 129609 284113
rect 129637 284085 129671 284113
rect 129699 284085 129747 284113
rect 129437 284051 129747 284085
rect 129437 284023 129485 284051
rect 129513 284023 129547 284051
rect 129575 284023 129609 284051
rect 129637 284023 129671 284051
rect 129699 284023 129747 284051
rect 129437 283989 129747 284023
rect 129437 283961 129485 283989
rect 129513 283961 129547 283989
rect 129575 283961 129609 283989
rect 129637 283961 129671 283989
rect 129699 283961 129747 283989
rect 129437 275175 129747 283961
rect 129437 275147 129485 275175
rect 129513 275147 129547 275175
rect 129575 275147 129609 275175
rect 129637 275147 129671 275175
rect 129699 275147 129747 275175
rect 129437 275113 129747 275147
rect 129437 275085 129485 275113
rect 129513 275085 129547 275113
rect 129575 275085 129609 275113
rect 129637 275085 129671 275113
rect 129699 275085 129747 275113
rect 129437 275051 129747 275085
rect 129437 275023 129485 275051
rect 129513 275023 129547 275051
rect 129575 275023 129609 275051
rect 129637 275023 129671 275051
rect 129699 275023 129747 275051
rect 129437 274989 129747 275023
rect 129437 274961 129485 274989
rect 129513 274961 129547 274989
rect 129575 274961 129609 274989
rect 129637 274961 129671 274989
rect 129699 274961 129747 274989
rect 129437 266175 129747 274961
rect 129437 266147 129485 266175
rect 129513 266147 129547 266175
rect 129575 266147 129609 266175
rect 129637 266147 129671 266175
rect 129699 266147 129747 266175
rect 129437 266113 129747 266147
rect 129437 266085 129485 266113
rect 129513 266085 129547 266113
rect 129575 266085 129609 266113
rect 129637 266085 129671 266113
rect 129699 266085 129747 266113
rect 129437 266051 129747 266085
rect 129437 266023 129485 266051
rect 129513 266023 129547 266051
rect 129575 266023 129609 266051
rect 129637 266023 129671 266051
rect 129699 266023 129747 266051
rect 129437 265989 129747 266023
rect 129437 265961 129485 265989
rect 129513 265961 129547 265989
rect 129575 265961 129609 265989
rect 129637 265961 129671 265989
rect 129699 265961 129747 265989
rect 129437 260603 129747 265961
rect 136577 298606 136887 299134
rect 136577 298578 136625 298606
rect 136653 298578 136687 298606
rect 136715 298578 136749 298606
rect 136777 298578 136811 298606
rect 136839 298578 136887 298606
rect 136577 298544 136887 298578
rect 136577 298516 136625 298544
rect 136653 298516 136687 298544
rect 136715 298516 136749 298544
rect 136777 298516 136811 298544
rect 136839 298516 136887 298544
rect 136577 298482 136887 298516
rect 136577 298454 136625 298482
rect 136653 298454 136687 298482
rect 136715 298454 136749 298482
rect 136777 298454 136811 298482
rect 136839 298454 136887 298482
rect 136577 298420 136887 298454
rect 136577 298392 136625 298420
rect 136653 298392 136687 298420
rect 136715 298392 136749 298420
rect 136777 298392 136811 298420
rect 136839 298392 136887 298420
rect 136577 290175 136887 298392
rect 136577 290147 136625 290175
rect 136653 290147 136687 290175
rect 136715 290147 136749 290175
rect 136777 290147 136811 290175
rect 136839 290147 136887 290175
rect 136577 290113 136887 290147
rect 136577 290085 136625 290113
rect 136653 290085 136687 290113
rect 136715 290085 136749 290113
rect 136777 290085 136811 290113
rect 136839 290085 136887 290113
rect 136577 290051 136887 290085
rect 136577 290023 136625 290051
rect 136653 290023 136687 290051
rect 136715 290023 136749 290051
rect 136777 290023 136811 290051
rect 136839 290023 136887 290051
rect 136577 289989 136887 290023
rect 136577 289961 136625 289989
rect 136653 289961 136687 289989
rect 136715 289961 136749 289989
rect 136777 289961 136811 289989
rect 136839 289961 136887 289989
rect 136577 281175 136887 289961
rect 136577 281147 136625 281175
rect 136653 281147 136687 281175
rect 136715 281147 136749 281175
rect 136777 281147 136811 281175
rect 136839 281147 136887 281175
rect 136577 281113 136887 281147
rect 136577 281085 136625 281113
rect 136653 281085 136687 281113
rect 136715 281085 136749 281113
rect 136777 281085 136811 281113
rect 136839 281085 136887 281113
rect 136577 281051 136887 281085
rect 136577 281023 136625 281051
rect 136653 281023 136687 281051
rect 136715 281023 136749 281051
rect 136777 281023 136811 281051
rect 136839 281023 136887 281051
rect 136577 280989 136887 281023
rect 136577 280961 136625 280989
rect 136653 280961 136687 280989
rect 136715 280961 136749 280989
rect 136777 280961 136811 280989
rect 136839 280961 136887 280989
rect 136577 272175 136887 280961
rect 136577 272147 136625 272175
rect 136653 272147 136687 272175
rect 136715 272147 136749 272175
rect 136777 272147 136811 272175
rect 136839 272147 136887 272175
rect 136577 272113 136887 272147
rect 136577 272085 136625 272113
rect 136653 272085 136687 272113
rect 136715 272085 136749 272113
rect 136777 272085 136811 272113
rect 136839 272085 136887 272113
rect 136577 272051 136887 272085
rect 136577 272023 136625 272051
rect 136653 272023 136687 272051
rect 136715 272023 136749 272051
rect 136777 272023 136811 272051
rect 136839 272023 136887 272051
rect 136577 271989 136887 272023
rect 136577 271961 136625 271989
rect 136653 271961 136687 271989
rect 136715 271961 136749 271989
rect 136777 271961 136811 271989
rect 136839 271961 136887 271989
rect 136577 263175 136887 271961
rect 136577 263147 136625 263175
rect 136653 263147 136687 263175
rect 136715 263147 136749 263175
rect 136777 263147 136811 263175
rect 136839 263147 136887 263175
rect 136577 263113 136887 263147
rect 136577 263085 136625 263113
rect 136653 263085 136687 263113
rect 136715 263085 136749 263113
rect 136777 263085 136811 263113
rect 136839 263085 136887 263113
rect 136577 263051 136887 263085
rect 136577 263023 136625 263051
rect 136653 263023 136687 263051
rect 136715 263023 136749 263051
rect 136777 263023 136811 263051
rect 136839 263023 136887 263051
rect 136577 262989 136887 263023
rect 136577 262961 136625 262989
rect 136653 262961 136687 262989
rect 136715 262961 136749 262989
rect 136777 262961 136811 262989
rect 136839 262961 136887 262989
rect 136577 260603 136887 262961
rect 138437 299086 138747 299134
rect 138437 299058 138485 299086
rect 138513 299058 138547 299086
rect 138575 299058 138609 299086
rect 138637 299058 138671 299086
rect 138699 299058 138747 299086
rect 138437 299024 138747 299058
rect 138437 298996 138485 299024
rect 138513 298996 138547 299024
rect 138575 298996 138609 299024
rect 138637 298996 138671 299024
rect 138699 298996 138747 299024
rect 138437 298962 138747 298996
rect 138437 298934 138485 298962
rect 138513 298934 138547 298962
rect 138575 298934 138609 298962
rect 138637 298934 138671 298962
rect 138699 298934 138747 298962
rect 138437 298900 138747 298934
rect 138437 298872 138485 298900
rect 138513 298872 138547 298900
rect 138575 298872 138609 298900
rect 138637 298872 138671 298900
rect 138699 298872 138747 298900
rect 138437 293175 138747 298872
rect 138437 293147 138485 293175
rect 138513 293147 138547 293175
rect 138575 293147 138609 293175
rect 138637 293147 138671 293175
rect 138699 293147 138747 293175
rect 138437 293113 138747 293147
rect 138437 293085 138485 293113
rect 138513 293085 138547 293113
rect 138575 293085 138609 293113
rect 138637 293085 138671 293113
rect 138699 293085 138747 293113
rect 138437 293051 138747 293085
rect 138437 293023 138485 293051
rect 138513 293023 138547 293051
rect 138575 293023 138609 293051
rect 138637 293023 138671 293051
rect 138699 293023 138747 293051
rect 138437 292989 138747 293023
rect 138437 292961 138485 292989
rect 138513 292961 138547 292989
rect 138575 292961 138609 292989
rect 138637 292961 138671 292989
rect 138699 292961 138747 292989
rect 138437 284175 138747 292961
rect 138437 284147 138485 284175
rect 138513 284147 138547 284175
rect 138575 284147 138609 284175
rect 138637 284147 138671 284175
rect 138699 284147 138747 284175
rect 138437 284113 138747 284147
rect 138437 284085 138485 284113
rect 138513 284085 138547 284113
rect 138575 284085 138609 284113
rect 138637 284085 138671 284113
rect 138699 284085 138747 284113
rect 138437 284051 138747 284085
rect 138437 284023 138485 284051
rect 138513 284023 138547 284051
rect 138575 284023 138609 284051
rect 138637 284023 138671 284051
rect 138699 284023 138747 284051
rect 138437 283989 138747 284023
rect 138437 283961 138485 283989
rect 138513 283961 138547 283989
rect 138575 283961 138609 283989
rect 138637 283961 138671 283989
rect 138699 283961 138747 283989
rect 138437 275175 138747 283961
rect 138437 275147 138485 275175
rect 138513 275147 138547 275175
rect 138575 275147 138609 275175
rect 138637 275147 138671 275175
rect 138699 275147 138747 275175
rect 138437 275113 138747 275147
rect 138437 275085 138485 275113
rect 138513 275085 138547 275113
rect 138575 275085 138609 275113
rect 138637 275085 138671 275113
rect 138699 275085 138747 275113
rect 138437 275051 138747 275085
rect 138437 275023 138485 275051
rect 138513 275023 138547 275051
rect 138575 275023 138609 275051
rect 138637 275023 138671 275051
rect 138699 275023 138747 275051
rect 138437 274989 138747 275023
rect 138437 274961 138485 274989
rect 138513 274961 138547 274989
rect 138575 274961 138609 274989
rect 138637 274961 138671 274989
rect 138699 274961 138747 274989
rect 138437 266175 138747 274961
rect 138437 266147 138485 266175
rect 138513 266147 138547 266175
rect 138575 266147 138609 266175
rect 138637 266147 138671 266175
rect 138699 266147 138747 266175
rect 138437 266113 138747 266147
rect 138437 266085 138485 266113
rect 138513 266085 138547 266113
rect 138575 266085 138609 266113
rect 138637 266085 138671 266113
rect 138699 266085 138747 266113
rect 138437 266051 138747 266085
rect 138437 266023 138485 266051
rect 138513 266023 138547 266051
rect 138575 266023 138609 266051
rect 138637 266023 138671 266051
rect 138699 266023 138747 266051
rect 138437 265989 138747 266023
rect 138437 265961 138485 265989
rect 138513 265961 138547 265989
rect 138575 265961 138609 265989
rect 138637 265961 138671 265989
rect 138699 265961 138747 265989
rect 138437 260603 138747 265961
rect 145577 298606 145887 299134
rect 145577 298578 145625 298606
rect 145653 298578 145687 298606
rect 145715 298578 145749 298606
rect 145777 298578 145811 298606
rect 145839 298578 145887 298606
rect 145577 298544 145887 298578
rect 145577 298516 145625 298544
rect 145653 298516 145687 298544
rect 145715 298516 145749 298544
rect 145777 298516 145811 298544
rect 145839 298516 145887 298544
rect 145577 298482 145887 298516
rect 145577 298454 145625 298482
rect 145653 298454 145687 298482
rect 145715 298454 145749 298482
rect 145777 298454 145811 298482
rect 145839 298454 145887 298482
rect 145577 298420 145887 298454
rect 145577 298392 145625 298420
rect 145653 298392 145687 298420
rect 145715 298392 145749 298420
rect 145777 298392 145811 298420
rect 145839 298392 145887 298420
rect 145577 290175 145887 298392
rect 145577 290147 145625 290175
rect 145653 290147 145687 290175
rect 145715 290147 145749 290175
rect 145777 290147 145811 290175
rect 145839 290147 145887 290175
rect 145577 290113 145887 290147
rect 145577 290085 145625 290113
rect 145653 290085 145687 290113
rect 145715 290085 145749 290113
rect 145777 290085 145811 290113
rect 145839 290085 145887 290113
rect 145577 290051 145887 290085
rect 145577 290023 145625 290051
rect 145653 290023 145687 290051
rect 145715 290023 145749 290051
rect 145777 290023 145811 290051
rect 145839 290023 145887 290051
rect 145577 289989 145887 290023
rect 145577 289961 145625 289989
rect 145653 289961 145687 289989
rect 145715 289961 145749 289989
rect 145777 289961 145811 289989
rect 145839 289961 145887 289989
rect 145577 281175 145887 289961
rect 145577 281147 145625 281175
rect 145653 281147 145687 281175
rect 145715 281147 145749 281175
rect 145777 281147 145811 281175
rect 145839 281147 145887 281175
rect 145577 281113 145887 281147
rect 145577 281085 145625 281113
rect 145653 281085 145687 281113
rect 145715 281085 145749 281113
rect 145777 281085 145811 281113
rect 145839 281085 145887 281113
rect 145577 281051 145887 281085
rect 145577 281023 145625 281051
rect 145653 281023 145687 281051
rect 145715 281023 145749 281051
rect 145777 281023 145811 281051
rect 145839 281023 145887 281051
rect 145577 280989 145887 281023
rect 145577 280961 145625 280989
rect 145653 280961 145687 280989
rect 145715 280961 145749 280989
rect 145777 280961 145811 280989
rect 145839 280961 145887 280989
rect 145577 272175 145887 280961
rect 145577 272147 145625 272175
rect 145653 272147 145687 272175
rect 145715 272147 145749 272175
rect 145777 272147 145811 272175
rect 145839 272147 145887 272175
rect 145577 272113 145887 272147
rect 145577 272085 145625 272113
rect 145653 272085 145687 272113
rect 145715 272085 145749 272113
rect 145777 272085 145811 272113
rect 145839 272085 145887 272113
rect 145577 272051 145887 272085
rect 145577 272023 145625 272051
rect 145653 272023 145687 272051
rect 145715 272023 145749 272051
rect 145777 272023 145811 272051
rect 145839 272023 145887 272051
rect 145577 271989 145887 272023
rect 145577 271961 145625 271989
rect 145653 271961 145687 271989
rect 145715 271961 145749 271989
rect 145777 271961 145811 271989
rect 145839 271961 145887 271989
rect 145577 263175 145887 271961
rect 145577 263147 145625 263175
rect 145653 263147 145687 263175
rect 145715 263147 145749 263175
rect 145777 263147 145811 263175
rect 145839 263147 145887 263175
rect 145577 263113 145887 263147
rect 145577 263085 145625 263113
rect 145653 263085 145687 263113
rect 145715 263085 145749 263113
rect 145777 263085 145811 263113
rect 145839 263085 145887 263113
rect 145577 263051 145887 263085
rect 145577 263023 145625 263051
rect 145653 263023 145687 263051
rect 145715 263023 145749 263051
rect 145777 263023 145811 263051
rect 145839 263023 145887 263051
rect 145577 262989 145887 263023
rect 145577 262961 145625 262989
rect 145653 262961 145687 262989
rect 145715 262961 145749 262989
rect 145777 262961 145811 262989
rect 145839 262961 145887 262989
rect 145577 260603 145887 262961
rect 147437 299086 147747 299134
rect 147437 299058 147485 299086
rect 147513 299058 147547 299086
rect 147575 299058 147609 299086
rect 147637 299058 147671 299086
rect 147699 299058 147747 299086
rect 147437 299024 147747 299058
rect 147437 298996 147485 299024
rect 147513 298996 147547 299024
rect 147575 298996 147609 299024
rect 147637 298996 147671 299024
rect 147699 298996 147747 299024
rect 147437 298962 147747 298996
rect 147437 298934 147485 298962
rect 147513 298934 147547 298962
rect 147575 298934 147609 298962
rect 147637 298934 147671 298962
rect 147699 298934 147747 298962
rect 147437 298900 147747 298934
rect 147437 298872 147485 298900
rect 147513 298872 147547 298900
rect 147575 298872 147609 298900
rect 147637 298872 147671 298900
rect 147699 298872 147747 298900
rect 147437 293175 147747 298872
rect 147437 293147 147485 293175
rect 147513 293147 147547 293175
rect 147575 293147 147609 293175
rect 147637 293147 147671 293175
rect 147699 293147 147747 293175
rect 147437 293113 147747 293147
rect 147437 293085 147485 293113
rect 147513 293085 147547 293113
rect 147575 293085 147609 293113
rect 147637 293085 147671 293113
rect 147699 293085 147747 293113
rect 147437 293051 147747 293085
rect 147437 293023 147485 293051
rect 147513 293023 147547 293051
rect 147575 293023 147609 293051
rect 147637 293023 147671 293051
rect 147699 293023 147747 293051
rect 147437 292989 147747 293023
rect 147437 292961 147485 292989
rect 147513 292961 147547 292989
rect 147575 292961 147609 292989
rect 147637 292961 147671 292989
rect 147699 292961 147747 292989
rect 147437 284175 147747 292961
rect 147437 284147 147485 284175
rect 147513 284147 147547 284175
rect 147575 284147 147609 284175
rect 147637 284147 147671 284175
rect 147699 284147 147747 284175
rect 147437 284113 147747 284147
rect 147437 284085 147485 284113
rect 147513 284085 147547 284113
rect 147575 284085 147609 284113
rect 147637 284085 147671 284113
rect 147699 284085 147747 284113
rect 147437 284051 147747 284085
rect 147437 284023 147485 284051
rect 147513 284023 147547 284051
rect 147575 284023 147609 284051
rect 147637 284023 147671 284051
rect 147699 284023 147747 284051
rect 147437 283989 147747 284023
rect 147437 283961 147485 283989
rect 147513 283961 147547 283989
rect 147575 283961 147609 283989
rect 147637 283961 147671 283989
rect 147699 283961 147747 283989
rect 147437 275175 147747 283961
rect 147437 275147 147485 275175
rect 147513 275147 147547 275175
rect 147575 275147 147609 275175
rect 147637 275147 147671 275175
rect 147699 275147 147747 275175
rect 147437 275113 147747 275147
rect 147437 275085 147485 275113
rect 147513 275085 147547 275113
rect 147575 275085 147609 275113
rect 147637 275085 147671 275113
rect 147699 275085 147747 275113
rect 147437 275051 147747 275085
rect 147437 275023 147485 275051
rect 147513 275023 147547 275051
rect 147575 275023 147609 275051
rect 147637 275023 147671 275051
rect 147699 275023 147747 275051
rect 147437 274989 147747 275023
rect 147437 274961 147485 274989
rect 147513 274961 147547 274989
rect 147575 274961 147609 274989
rect 147637 274961 147671 274989
rect 147699 274961 147747 274989
rect 147437 266175 147747 274961
rect 147437 266147 147485 266175
rect 147513 266147 147547 266175
rect 147575 266147 147609 266175
rect 147637 266147 147671 266175
rect 147699 266147 147747 266175
rect 147437 266113 147747 266147
rect 147437 266085 147485 266113
rect 147513 266085 147547 266113
rect 147575 266085 147609 266113
rect 147637 266085 147671 266113
rect 147699 266085 147747 266113
rect 147437 266051 147747 266085
rect 147437 266023 147485 266051
rect 147513 266023 147547 266051
rect 147575 266023 147609 266051
rect 147637 266023 147671 266051
rect 147699 266023 147747 266051
rect 147437 265989 147747 266023
rect 147437 265961 147485 265989
rect 147513 265961 147547 265989
rect 147575 265961 147609 265989
rect 147637 265961 147671 265989
rect 147699 265961 147747 265989
rect 147437 260603 147747 265961
rect 154577 298606 154887 299134
rect 154577 298578 154625 298606
rect 154653 298578 154687 298606
rect 154715 298578 154749 298606
rect 154777 298578 154811 298606
rect 154839 298578 154887 298606
rect 154577 298544 154887 298578
rect 154577 298516 154625 298544
rect 154653 298516 154687 298544
rect 154715 298516 154749 298544
rect 154777 298516 154811 298544
rect 154839 298516 154887 298544
rect 154577 298482 154887 298516
rect 154577 298454 154625 298482
rect 154653 298454 154687 298482
rect 154715 298454 154749 298482
rect 154777 298454 154811 298482
rect 154839 298454 154887 298482
rect 154577 298420 154887 298454
rect 154577 298392 154625 298420
rect 154653 298392 154687 298420
rect 154715 298392 154749 298420
rect 154777 298392 154811 298420
rect 154839 298392 154887 298420
rect 154577 290175 154887 298392
rect 154577 290147 154625 290175
rect 154653 290147 154687 290175
rect 154715 290147 154749 290175
rect 154777 290147 154811 290175
rect 154839 290147 154887 290175
rect 154577 290113 154887 290147
rect 154577 290085 154625 290113
rect 154653 290085 154687 290113
rect 154715 290085 154749 290113
rect 154777 290085 154811 290113
rect 154839 290085 154887 290113
rect 154577 290051 154887 290085
rect 154577 290023 154625 290051
rect 154653 290023 154687 290051
rect 154715 290023 154749 290051
rect 154777 290023 154811 290051
rect 154839 290023 154887 290051
rect 154577 289989 154887 290023
rect 154577 289961 154625 289989
rect 154653 289961 154687 289989
rect 154715 289961 154749 289989
rect 154777 289961 154811 289989
rect 154839 289961 154887 289989
rect 154577 281175 154887 289961
rect 154577 281147 154625 281175
rect 154653 281147 154687 281175
rect 154715 281147 154749 281175
rect 154777 281147 154811 281175
rect 154839 281147 154887 281175
rect 154577 281113 154887 281147
rect 154577 281085 154625 281113
rect 154653 281085 154687 281113
rect 154715 281085 154749 281113
rect 154777 281085 154811 281113
rect 154839 281085 154887 281113
rect 154577 281051 154887 281085
rect 154577 281023 154625 281051
rect 154653 281023 154687 281051
rect 154715 281023 154749 281051
rect 154777 281023 154811 281051
rect 154839 281023 154887 281051
rect 154577 280989 154887 281023
rect 154577 280961 154625 280989
rect 154653 280961 154687 280989
rect 154715 280961 154749 280989
rect 154777 280961 154811 280989
rect 154839 280961 154887 280989
rect 154577 272175 154887 280961
rect 154577 272147 154625 272175
rect 154653 272147 154687 272175
rect 154715 272147 154749 272175
rect 154777 272147 154811 272175
rect 154839 272147 154887 272175
rect 154577 272113 154887 272147
rect 154577 272085 154625 272113
rect 154653 272085 154687 272113
rect 154715 272085 154749 272113
rect 154777 272085 154811 272113
rect 154839 272085 154887 272113
rect 154577 272051 154887 272085
rect 154577 272023 154625 272051
rect 154653 272023 154687 272051
rect 154715 272023 154749 272051
rect 154777 272023 154811 272051
rect 154839 272023 154887 272051
rect 154577 271989 154887 272023
rect 154577 271961 154625 271989
rect 154653 271961 154687 271989
rect 154715 271961 154749 271989
rect 154777 271961 154811 271989
rect 154839 271961 154887 271989
rect 154577 263175 154887 271961
rect 154577 263147 154625 263175
rect 154653 263147 154687 263175
rect 154715 263147 154749 263175
rect 154777 263147 154811 263175
rect 154839 263147 154887 263175
rect 154577 263113 154887 263147
rect 154577 263085 154625 263113
rect 154653 263085 154687 263113
rect 154715 263085 154749 263113
rect 154777 263085 154811 263113
rect 154839 263085 154887 263113
rect 154577 263051 154887 263085
rect 154577 263023 154625 263051
rect 154653 263023 154687 263051
rect 154715 263023 154749 263051
rect 154777 263023 154811 263051
rect 154839 263023 154887 263051
rect 154577 262989 154887 263023
rect 154577 262961 154625 262989
rect 154653 262961 154687 262989
rect 154715 262961 154749 262989
rect 154777 262961 154811 262989
rect 154839 262961 154887 262989
rect 48437 257147 48485 257175
rect 48513 257147 48547 257175
rect 48575 257147 48609 257175
rect 48637 257147 48671 257175
rect 48699 257147 48747 257175
rect 48437 257113 48747 257147
rect 48437 257085 48485 257113
rect 48513 257085 48547 257113
rect 48575 257085 48609 257113
rect 48637 257085 48671 257113
rect 48699 257085 48747 257113
rect 48437 257051 48747 257085
rect 48437 257023 48485 257051
rect 48513 257023 48547 257051
rect 48575 257023 48609 257051
rect 48637 257023 48671 257051
rect 48699 257023 48747 257051
rect 48437 256989 48747 257023
rect 48437 256961 48485 256989
rect 48513 256961 48547 256989
rect 48575 256961 48609 256989
rect 48637 256961 48671 256989
rect 48699 256961 48747 256989
rect 48437 248175 48747 256961
rect 59904 257175 60064 257192
rect 59904 257147 59939 257175
rect 59967 257147 60001 257175
rect 60029 257147 60064 257175
rect 59904 257113 60064 257147
rect 59904 257085 59939 257113
rect 59967 257085 60001 257113
rect 60029 257085 60064 257113
rect 59904 257051 60064 257085
rect 59904 257023 59939 257051
rect 59967 257023 60001 257051
rect 60029 257023 60064 257051
rect 59904 256989 60064 257023
rect 59904 256961 59939 256989
rect 59967 256961 60001 256989
rect 60029 256961 60064 256989
rect 59904 256944 60064 256961
rect 75264 257175 75424 257192
rect 75264 257147 75299 257175
rect 75327 257147 75361 257175
rect 75389 257147 75424 257175
rect 75264 257113 75424 257147
rect 75264 257085 75299 257113
rect 75327 257085 75361 257113
rect 75389 257085 75424 257113
rect 75264 257051 75424 257085
rect 75264 257023 75299 257051
rect 75327 257023 75361 257051
rect 75389 257023 75424 257051
rect 75264 256989 75424 257023
rect 75264 256961 75299 256989
rect 75327 256961 75361 256989
rect 75389 256961 75424 256989
rect 75264 256944 75424 256961
rect 90624 257175 90784 257192
rect 90624 257147 90659 257175
rect 90687 257147 90721 257175
rect 90749 257147 90784 257175
rect 90624 257113 90784 257147
rect 90624 257085 90659 257113
rect 90687 257085 90721 257113
rect 90749 257085 90784 257113
rect 90624 257051 90784 257085
rect 90624 257023 90659 257051
rect 90687 257023 90721 257051
rect 90749 257023 90784 257051
rect 90624 256989 90784 257023
rect 90624 256961 90659 256989
rect 90687 256961 90721 256989
rect 90749 256961 90784 256989
rect 90624 256944 90784 256961
rect 105984 257175 106144 257192
rect 105984 257147 106019 257175
rect 106047 257147 106081 257175
rect 106109 257147 106144 257175
rect 105984 257113 106144 257147
rect 105984 257085 106019 257113
rect 106047 257085 106081 257113
rect 106109 257085 106144 257113
rect 105984 257051 106144 257085
rect 105984 257023 106019 257051
rect 106047 257023 106081 257051
rect 106109 257023 106144 257051
rect 105984 256989 106144 257023
rect 105984 256961 106019 256989
rect 106047 256961 106081 256989
rect 106109 256961 106144 256989
rect 105984 256944 106144 256961
rect 121344 257175 121504 257192
rect 121344 257147 121379 257175
rect 121407 257147 121441 257175
rect 121469 257147 121504 257175
rect 121344 257113 121504 257147
rect 121344 257085 121379 257113
rect 121407 257085 121441 257113
rect 121469 257085 121504 257113
rect 121344 257051 121504 257085
rect 121344 257023 121379 257051
rect 121407 257023 121441 257051
rect 121469 257023 121504 257051
rect 121344 256989 121504 257023
rect 121344 256961 121379 256989
rect 121407 256961 121441 256989
rect 121469 256961 121504 256989
rect 121344 256944 121504 256961
rect 136704 257175 136864 257192
rect 136704 257147 136739 257175
rect 136767 257147 136801 257175
rect 136829 257147 136864 257175
rect 136704 257113 136864 257147
rect 136704 257085 136739 257113
rect 136767 257085 136801 257113
rect 136829 257085 136864 257113
rect 136704 257051 136864 257085
rect 136704 257023 136739 257051
rect 136767 257023 136801 257051
rect 136829 257023 136864 257051
rect 136704 256989 136864 257023
rect 136704 256961 136739 256989
rect 136767 256961 136801 256989
rect 136829 256961 136864 256989
rect 136704 256944 136864 256961
rect 52224 254175 52384 254192
rect 52224 254147 52259 254175
rect 52287 254147 52321 254175
rect 52349 254147 52384 254175
rect 52224 254113 52384 254147
rect 52224 254085 52259 254113
rect 52287 254085 52321 254113
rect 52349 254085 52384 254113
rect 52224 254051 52384 254085
rect 52224 254023 52259 254051
rect 52287 254023 52321 254051
rect 52349 254023 52384 254051
rect 52224 253989 52384 254023
rect 52224 253961 52259 253989
rect 52287 253961 52321 253989
rect 52349 253961 52384 253989
rect 52224 253944 52384 253961
rect 67584 254175 67744 254192
rect 67584 254147 67619 254175
rect 67647 254147 67681 254175
rect 67709 254147 67744 254175
rect 67584 254113 67744 254147
rect 67584 254085 67619 254113
rect 67647 254085 67681 254113
rect 67709 254085 67744 254113
rect 67584 254051 67744 254085
rect 67584 254023 67619 254051
rect 67647 254023 67681 254051
rect 67709 254023 67744 254051
rect 67584 253989 67744 254023
rect 67584 253961 67619 253989
rect 67647 253961 67681 253989
rect 67709 253961 67744 253989
rect 67584 253944 67744 253961
rect 82944 254175 83104 254192
rect 82944 254147 82979 254175
rect 83007 254147 83041 254175
rect 83069 254147 83104 254175
rect 82944 254113 83104 254147
rect 82944 254085 82979 254113
rect 83007 254085 83041 254113
rect 83069 254085 83104 254113
rect 82944 254051 83104 254085
rect 82944 254023 82979 254051
rect 83007 254023 83041 254051
rect 83069 254023 83104 254051
rect 82944 253989 83104 254023
rect 82944 253961 82979 253989
rect 83007 253961 83041 253989
rect 83069 253961 83104 253989
rect 82944 253944 83104 253961
rect 98304 254175 98464 254192
rect 98304 254147 98339 254175
rect 98367 254147 98401 254175
rect 98429 254147 98464 254175
rect 98304 254113 98464 254147
rect 98304 254085 98339 254113
rect 98367 254085 98401 254113
rect 98429 254085 98464 254113
rect 98304 254051 98464 254085
rect 98304 254023 98339 254051
rect 98367 254023 98401 254051
rect 98429 254023 98464 254051
rect 98304 253989 98464 254023
rect 98304 253961 98339 253989
rect 98367 253961 98401 253989
rect 98429 253961 98464 253989
rect 98304 253944 98464 253961
rect 113664 254175 113824 254192
rect 113664 254147 113699 254175
rect 113727 254147 113761 254175
rect 113789 254147 113824 254175
rect 113664 254113 113824 254147
rect 113664 254085 113699 254113
rect 113727 254085 113761 254113
rect 113789 254085 113824 254113
rect 113664 254051 113824 254085
rect 113664 254023 113699 254051
rect 113727 254023 113761 254051
rect 113789 254023 113824 254051
rect 113664 253989 113824 254023
rect 113664 253961 113699 253989
rect 113727 253961 113761 253989
rect 113789 253961 113824 253989
rect 113664 253944 113824 253961
rect 129024 254175 129184 254192
rect 129024 254147 129059 254175
rect 129087 254147 129121 254175
rect 129149 254147 129184 254175
rect 129024 254113 129184 254147
rect 129024 254085 129059 254113
rect 129087 254085 129121 254113
rect 129149 254085 129184 254113
rect 129024 254051 129184 254085
rect 129024 254023 129059 254051
rect 129087 254023 129121 254051
rect 129149 254023 129184 254051
rect 129024 253989 129184 254023
rect 129024 253961 129059 253989
rect 129087 253961 129121 253989
rect 129149 253961 129184 253989
rect 129024 253944 129184 253961
rect 144384 254175 144544 254192
rect 144384 254147 144419 254175
rect 144447 254147 144481 254175
rect 144509 254147 144544 254175
rect 144384 254113 144544 254147
rect 144384 254085 144419 254113
rect 144447 254085 144481 254113
rect 144509 254085 144544 254113
rect 144384 254051 144544 254085
rect 144384 254023 144419 254051
rect 144447 254023 144481 254051
rect 144509 254023 144544 254051
rect 144384 253989 144544 254023
rect 144384 253961 144419 253989
rect 144447 253961 144481 253989
rect 144509 253961 144544 253989
rect 144384 253944 144544 253961
rect 154577 254175 154887 262961
rect 154577 254147 154625 254175
rect 154653 254147 154687 254175
rect 154715 254147 154749 254175
rect 154777 254147 154811 254175
rect 154839 254147 154887 254175
rect 154577 254113 154887 254147
rect 154577 254085 154625 254113
rect 154653 254085 154687 254113
rect 154715 254085 154749 254113
rect 154777 254085 154811 254113
rect 154839 254085 154887 254113
rect 154577 254051 154887 254085
rect 154577 254023 154625 254051
rect 154653 254023 154687 254051
rect 154715 254023 154749 254051
rect 154777 254023 154811 254051
rect 154839 254023 154887 254051
rect 154577 253989 154887 254023
rect 154577 253961 154625 253989
rect 154653 253961 154687 253989
rect 154715 253961 154749 253989
rect 154777 253961 154811 253989
rect 154839 253961 154887 253989
rect 48437 248147 48485 248175
rect 48513 248147 48547 248175
rect 48575 248147 48609 248175
rect 48637 248147 48671 248175
rect 48699 248147 48747 248175
rect 48437 248113 48747 248147
rect 48437 248085 48485 248113
rect 48513 248085 48547 248113
rect 48575 248085 48609 248113
rect 48637 248085 48671 248113
rect 48699 248085 48747 248113
rect 48437 248051 48747 248085
rect 48437 248023 48485 248051
rect 48513 248023 48547 248051
rect 48575 248023 48609 248051
rect 48637 248023 48671 248051
rect 48699 248023 48747 248051
rect 48437 247989 48747 248023
rect 48437 247961 48485 247989
rect 48513 247961 48547 247989
rect 48575 247961 48609 247989
rect 48637 247961 48671 247989
rect 48699 247961 48747 247989
rect 48437 239175 48747 247961
rect 59904 248175 60064 248192
rect 59904 248147 59939 248175
rect 59967 248147 60001 248175
rect 60029 248147 60064 248175
rect 59904 248113 60064 248147
rect 59904 248085 59939 248113
rect 59967 248085 60001 248113
rect 60029 248085 60064 248113
rect 59904 248051 60064 248085
rect 59904 248023 59939 248051
rect 59967 248023 60001 248051
rect 60029 248023 60064 248051
rect 59904 247989 60064 248023
rect 59904 247961 59939 247989
rect 59967 247961 60001 247989
rect 60029 247961 60064 247989
rect 59904 247944 60064 247961
rect 75264 248175 75424 248192
rect 75264 248147 75299 248175
rect 75327 248147 75361 248175
rect 75389 248147 75424 248175
rect 75264 248113 75424 248147
rect 75264 248085 75299 248113
rect 75327 248085 75361 248113
rect 75389 248085 75424 248113
rect 75264 248051 75424 248085
rect 75264 248023 75299 248051
rect 75327 248023 75361 248051
rect 75389 248023 75424 248051
rect 75264 247989 75424 248023
rect 75264 247961 75299 247989
rect 75327 247961 75361 247989
rect 75389 247961 75424 247989
rect 75264 247944 75424 247961
rect 90624 248175 90784 248192
rect 90624 248147 90659 248175
rect 90687 248147 90721 248175
rect 90749 248147 90784 248175
rect 90624 248113 90784 248147
rect 90624 248085 90659 248113
rect 90687 248085 90721 248113
rect 90749 248085 90784 248113
rect 90624 248051 90784 248085
rect 90624 248023 90659 248051
rect 90687 248023 90721 248051
rect 90749 248023 90784 248051
rect 90624 247989 90784 248023
rect 90624 247961 90659 247989
rect 90687 247961 90721 247989
rect 90749 247961 90784 247989
rect 90624 247944 90784 247961
rect 105984 248175 106144 248192
rect 105984 248147 106019 248175
rect 106047 248147 106081 248175
rect 106109 248147 106144 248175
rect 105984 248113 106144 248147
rect 105984 248085 106019 248113
rect 106047 248085 106081 248113
rect 106109 248085 106144 248113
rect 105984 248051 106144 248085
rect 105984 248023 106019 248051
rect 106047 248023 106081 248051
rect 106109 248023 106144 248051
rect 105984 247989 106144 248023
rect 105984 247961 106019 247989
rect 106047 247961 106081 247989
rect 106109 247961 106144 247989
rect 105984 247944 106144 247961
rect 121344 248175 121504 248192
rect 121344 248147 121379 248175
rect 121407 248147 121441 248175
rect 121469 248147 121504 248175
rect 121344 248113 121504 248147
rect 121344 248085 121379 248113
rect 121407 248085 121441 248113
rect 121469 248085 121504 248113
rect 121344 248051 121504 248085
rect 121344 248023 121379 248051
rect 121407 248023 121441 248051
rect 121469 248023 121504 248051
rect 121344 247989 121504 248023
rect 121344 247961 121379 247989
rect 121407 247961 121441 247989
rect 121469 247961 121504 247989
rect 121344 247944 121504 247961
rect 136704 248175 136864 248192
rect 136704 248147 136739 248175
rect 136767 248147 136801 248175
rect 136829 248147 136864 248175
rect 136704 248113 136864 248147
rect 136704 248085 136739 248113
rect 136767 248085 136801 248113
rect 136829 248085 136864 248113
rect 136704 248051 136864 248085
rect 136704 248023 136739 248051
rect 136767 248023 136801 248051
rect 136829 248023 136864 248051
rect 136704 247989 136864 248023
rect 136704 247961 136739 247989
rect 136767 247961 136801 247989
rect 136829 247961 136864 247989
rect 136704 247944 136864 247961
rect 52224 245175 52384 245192
rect 52224 245147 52259 245175
rect 52287 245147 52321 245175
rect 52349 245147 52384 245175
rect 52224 245113 52384 245147
rect 52224 245085 52259 245113
rect 52287 245085 52321 245113
rect 52349 245085 52384 245113
rect 52224 245051 52384 245085
rect 52224 245023 52259 245051
rect 52287 245023 52321 245051
rect 52349 245023 52384 245051
rect 52224 244989 52384 245023
rect 52224 244961 52259 244989
rect 52287 244961 52321 244989
rect 52349 244961 52384 244989
rect 52224 244944 52384 244961
rect 67584 245175 67744 245192
rect 67584 245147 67619 245175
rect 67647 245147 67681 245175
rect 67709 245147 67744 245175
rect 67584 245113 67744 245147
rect 67584 245085 67619 245113
rect 67647 245085 67681 245113
rect 67709 245085 67744 245113
rect 67584 245051 67744 245085
rect 67584 245023 67619 245051
rect 67647 245023 67681 245051
rect 67709 245023 67744 245051
rect 67584 244989 67744 245023
rect 67584 244961 67619 244989
rect 67647 244961 67681 244989
rect 67709 244961 67744 244989
rect 67584 244944 67744 244961
rect 82944 245175 83104 245192
rect 82944 245147 82979 245175
rect 83007 245147 83041 245175
rect 83069 245147 83104 245175
rect 82944 245113 83104 245147
rect 82944 245085 82979 245113
rect 83007 245085 83041 245113
rect 83069 245085 83104 245113
rect 82944 245051 83104 245085
rect 82944 245023 82979 245051
rect 83007 245023 83041 245051
rect 83069 245023 83104 245051
rect 82944 244989 83104 245023
rect 82944 244961 82979 244989
rect 83007 244961 83041 244989
rect 83069 244961 83104 244989
rect 82944 244944 83104 244961
rect 98304 245175 98464 245192
rect 98304 245147 98339 245175
rect 98367 245147 98401 245175
rect 98429 245147 98464 245175
rect 98304 245113 98464 245147
rect 98304 245085 98339 245113
rect 98367 245085 98401 245113
rect 98429 245085 98464 245113
rect 98304 245051 98464 245085
rect 98304 245023 98339 245051
rect 98367 245023 98401 245051
rect 98429 245023 98464 245051
rect 98304 244989 98464 245023
rect 98304 244961 98339 244989
rect 98367 244961 98401 244989
rect 98429 244961 98464 244989
rect 98304 244944 98464 244961
rect 113664 245175 113824 245192
rect 113664 245147 113699 245175
rect 113727 245147 113761 245175
rect 113789 245147 113824 245175
rect 113664 245113 113824 245147
rect 113664 245085 113699 245113
rect 113727 245085 113761 245113
rect 113789 245085 113824 245113
rect 113664 245051 113824 245085
rect 113664 245023 113699 245051
rect 113727 245023 113761 245051
rect 113789 245023 113824 245051
rect 113664 244989 113824 245023
rect 113664 244961 113699 244989
rect 113727 244961 113761 244989
rect 113789 244961 113824 244989
rect 113664 244944 113824 244961
rect 129024 245175 129184 245192
rect 129024 245147 129059 245175
rect 129087 245147 129121 245175
rect 129149 245147 129184 245175
rect 129024 245113 129184 245147
rect 129024 245085 129059 245113
rect 129087 245085 129121 245113
rect 129149 245085 129184 245113
rect 129024 245051 129184 245085
rect 129024 245023 129059 245051
rect 129087 245023 129121 245051
rect 129149 245023 129184 245051
rect 129024 244989 129184 245023
rect 129024 244961 129059 244989
rect 129087 244961 129121 244989
rect 129149 244961 129184 244989
rect 129024 244944 129184 244961
rect 144384 245175 144544 245192
rect 144384 245147 144419 245175
rect 144447 245147 144481 245175
rect 144509 245147 144544 245175
rect 144384 245113 144544 245147
rect 144384 245085 144419 245113
rect 144447 245085 144481 245113
rect 144509 245085 144544 245113
rect 144384 245051 144544 245085
rect 144384 245023 144419 245051
rect 144447 245023 144481 245051
rect 144509 245023 144544 245051
rect 144384 244989 144544 245023
rect 144384 244961 144419 244989
rect 144447 244961 144481 244989
rect 144509 244961 144544 244989
rect 144384 244944 144544 244961
rect 154577 245175 154887 253961
rect 154577 245147 154625 245175
rect 154653 245147 154687 245175
rect 154715 245147 154749 245175
rect 154777 245147 154811 245175
rect 154839 245147 154887 245175
rect 154577 245113 154887 245147
rect 154577 245085 154625 245113
rect 154653 245085 154687 245113
rect 154715 245085 154749 245113
rect 154777 245085 154811 245113
rect 154839 245085 154887 245113
rect 154577 245051 154887 245085
rect 154577 245023 154625 245051
rect 154653 245023 154687 245051
rect 154715 245023 154749 245051
rect 154777 245023 154811 245051
rect 154839 245023 154887 245051
rect 154577 244989 154887 245023
rect 154577 244961 154625 244989
rect 154653 244961 154687 244989
rect 154715 244961 154749 244989
rect 154777 244961 154811 244989
rect 154839 244961 154887 244989
rect 48437 239147 48485 239175
rect 48513 239147 48547 239175
rect 48575 239147 48609 239175
rect 48637 239147 48671 239175
rect 48699 239147 48747 239175
rect 48437 239113 48747 239147
rect 48437 239085 48485 239113
rect 48513 239085 48547 239113
rect 48575 239085 48609 239113
rect 48637 239085 48671 239113
rect 48699 239085 48747 239113
rect 48437 239051 48747 239085
rect 48437 239023 48485 239051
rect 48513 239023 48547 239051
rect 48575 239023 48609 239051
rect 48637 239023 48671 239051
rect 48699 239023 48747 239051
rect 48437 238989 48747 239023
rect 48437 238961 48485 238989
rect 48513 238961 48547 238989
rect 48575 238961 48609 238989
rect 48637 238961 48671 238989
rect 48699 238961 48747 238989
rect 48437 230175 48747 238961
rect 59904 239175 60064 239192
rect 59904 239147 59939 239175
rect 59967 239147 60001 239175
rect 60029 239147 60064 239175
rect 59904 239113 60064 239147
rect 59904 239085 59939 239113
rect 59967 239085 60001 239113
rect 60029 239085 60064 239113
rect 59904 239051 60064 239085
rect 59904 239023 59939 239051
rect 59967 239023 60001 239051
rect 60029 239023 60064 239051
rect 59904 238989 60064 239023
rect 59904 238961 59939 238989
rect 59967 238961 60001 238989
rect 60029 238961 60064 238989
rect 59904 238944 60064 238961
rect 75264 239175 75424 239192
rect 75264 239147 75299 239175
rect 75327 239147 75361 239175
rect 75389 239147 75424 239175
rect 75264 239113 75424 239147
rect 75264 239085 75299 239113
rect 75327 239085 75361 239113
rect 75389 239085 75424 239113
rect 75264 239051 75424 239085
rect 75264 239023 75299 239051
rect 75327 239023 75361 239051
rect 75389 239023 75424 239051
rect 75264 238989 75424 239023
rect 75264 238961 75299 238989
rect 75327 238961 75361 238989
rect 75389 238961 75424 238989
rect 75264 238944 75424 238961
rect 90624 239175 90784 239192
rect 90624 239147 90659 239175
rect 90687 239147 90721 239175
rect 90749 239147 90784 239175
rect 90624 239113 90784 239147
rect 90624 239085 90659 239113
rect 90687 239085 90721 239113
rect 90749 239085 90784 239113
rect 90624 239051 90784 239085
rect 90624 239023 90659 239051
rect 90687 239023 90721 239051
rect 90749 239023 90784 239051
rect 90624 238989 90784 239023
rect 90624 238961 90659 238989
rect 90687 238961 90721 238989
rect 90749 238961 90784 238989
rect 90624 238944 90784 238961
rect 105984 239175 106144 239192
rect 105984 239147 106019 239175
rect 106047 239147 106081 239175
rect 106109 239147 106144 239175
rect 105984 239113 106144 239147
rect 105984 239085 106019 239113
rect 106047 239085 106081 239113
rect 106109 239085 106144 239113
rect 105984 239051 106144 239085
rect 105984 239023 106019 239051
rect 106047 239023 106081 239051
rect 106109 239023 106144 239051
rect 105984 238989 106144 239023
rect 105984 238961 106019 238989
rect 106047 238961 106081 238989
rect 106109 238961 106144 238989
rect 105984 238944 106144 238961
rect 121344 239175 121504 239192
rect 121344 239147 121379 239175
rect 121407 239147 121441 239175
rect 121469 239147 121504 239175
rect 121344 239113 121504 239147
rect 121344 239085 121379 239113
rect 121407 239085 121441 239113
rect 121469 239085 121504 239113
rect 121344 239051 121504 239085
rect 121344 239023 121379 239051
rect 121407 239023 121441 239051
rect 121469 239023 121504 239051
rect 121344 238989 121504 239023
rect 121344 238961 121379 238989
rect 121407 238961 121441 238989
rect 121469 238961 121504 238989
rect 121344 238944 121504 238961
rect 136704 239175 136864 239192
rect 136704 239147 136739 239175
rect 136767 239147 136801 239175
rect 136829 239147 136864 239175
rect 136704 239113 136864 239147
rect 136704 239085 136739 239113
rect 136767 239085 136801 239113
rect 136829 239085 136864 239113
rect 136704 239051 136864 239085
rect 136704 239023 136739 239051
rect 136767 239023 136801 239051
rect 136829 239023 136864 239051
rect 136704 238989 136864 239023
rect 136704 238961 136739 238989
rect 136767 238961 136801 238989
rect 136829 238961 136864 238989
rect 136704 238944 136864 238961
rect 52224 236175 52384 236192
rect 52224 236147 52259 236175
rect 52287 236147 52321 236175
rect 52349 236147 52384 236175
rect 52224 236113 52384 236147
rect 52224 236085 52259 236113
rect 52287 236085 52321 236113
rect 52349 236085 52384 236113
rect 52224 236051 52384 236085
rect 52224 236023 52259 236051
rect 52287 236023 52321 236051
rect 52349 236023 52384 236051
rect 52224 235989 52384 236023
rect 52224 235961 52259 235989
rect 52287 235961 52321 235989
rect 52349 235961 52384 235989
rect 52224 235944 52384 235961
rect 67584 236175 67744 236192
rect 67584 236147 67619 236175
rect 67647 236147 67681 236175
rect 67709 236147 67744 236175
rect 67584 236113 67744 236147
rect 67584 236085 67619 236113
rect 67647 236085 67681 236113
rect 67709 236085 67744 236113
rect 67584 236051 67744 236085
rect 67584 236023 67619 236051
rect 67647 236023 67681 236051
rect 67709 236023 67744 236051
rect 67584 235989 67744 236023
rect 67584 235961 67619 235989
rect 67647 235961 67681 235989
rect 67709 235961 67744 235989
rect 67584 235944 67744 235961
rect 82944 236175 83104 236192
rect 82944 236147 82979 236175
rect 83007 236147 83041 236175
rect 83069 236147 83104 236175
rect 82944 236113 83104 236147
rect 82944 236085 82979 236113
rect 83007 236085 83041 236113
rect 83069 236085 83104 236113
rect 82944 236051 83104 236085
rect 82944 236023 82979 236051
rect 83007 236023 83041 236051
rect 83069 236023 83104 236051
rect 82944 235989 83104 236023
rect 82944 235961 82979 235989
rect 83007 235961 83041 235989
rect 83069 235961 83104 235989
rect 82944 235944 83104 235961
rect 98304 236175 98464 236192
rect 98304 236147 98339 236175
rect 98367 236147 98401 236175
rect 98429 236147 98464 236175
rect 98304 236113 98464 236147
rect 98304 236085 98339 236113
rect 98367 236085 98401 236113
rect 98429 236085 98464 236113
rect 98304 236051 98464 236085
rect 98304 236023 98339 236051
rect 98367 236023 98401 236051
rect 98429 236023 98464 236051
rect 98304 235989 98464 236023
rect 98304 235961 98339 235989
rect 98367 235961 98401 235989
rect 98429 235961 98464 235989
rect 98304 235944 98464 235961
rect 113664 236175 113824 236192
rect 113664 236147 113699 236175
rect 113727 236147 113761 236175
rect 113789 236147 113824 236175
rect 113664 236113 113824 236147
rect 113664 236085 113699 236113
rect 113727 236085 113761 236113
rect 113789 236085 113824 236113
rect 113664 236051 113824 236085
rect 113664 236023 113699 236051
rect 113727 236023 113761 236051
rect 113789 236023 113824 236051
rect 113664 235989 113824 236023
rect 113664 235961 113699 235989
rect 113727 235961 113761 235989
rect 113789 235961 113824 235989
rect 113664 235944 113824 235961
rect 129024 236175 129184 236192
rect 129024 236147 129059 236175
rect 129087 236147 129121 236175
rect 129149 236147 129184 236175
rect 129024 236113 129184 236147
rect 129024 236085 129059 236113
rect 129087 236085 129121 236113
rect 129149 236085 129184 236113
rect 129024 236051 129184 236085
rect 129024 236023 129059 236051
rect 129087 236023 129121 236051
rect 129149 236023 129184 236051
rect 129024 235989 129184 236023
rect 129024 235961 129059 235989
rect 129087 235961 129121 235989
rect 129149 235961 129184 235989
rect 129024 235944 129184 235961
rect 144384 236175 144544 236192
rect 144384 236147 144419 236175
rect 144447 236147 144481 236175
rect 144509 236147 144544 236175
rect 144384 236113 144544 236147
rect 144384 236085 144419 236113
rect 144447 236085 144481 236113
rect 144509 236085 144544 236113
rect 144384 236051 144544 236085
rect 144384 236023 144419 236051
rect 144447 236023 144481 236051
rect 144509 236023 144544 236051
rect 144384 235989 144544 236023
rect 144384 235961 144419 235989
rect 144447 235961 144481 235989
rect 144509 235961 144544 235989
rect 144384 235944 144544 235961
rect 154577 236175 154887 244961
rect 154577 236147 154625 236175
rect 154653 236147 154687 236175
rect 154715 236147 154749 236175
rect 154777 236147 154811 236175
rect 154839 236147 154887 236175
rect 154577 236113 154887 236147
rect 154577 236085 154625 236113
rect 154653 236085 154687 236113
rect 154715 236085 154749 236113
rect 154777 236085 154811 236113
rect 154839 236085 154887 236113
rect 154577 236051 154887 236085
rect 154577 236023 154625 236051
rect 154653 236023 154687 236051
rect 154715 236023 154749 236051
rect 154777 236023 154811 236051
rect 154839 236023 154887 236051
rect 154577 235989 154887 236023
rect 154577 235961 154625 235989
rect 154653 235961 154687 235989
rect 154715 235961 154749 235989
rect 154777 235961 154811 235989
rect 154839 235961 154887 235989
rect 48437 230147 48485 230175
rect 48513 230147 48547 230175
rect 48575 230147 48609 230175
rect 48637 230147 48671 230175
rect 48699 230147 48747 230175
rect 48437 230113 48747 230147
rect 48437 230085 48485 230113
rect 48513 230085 48547 230113
rect 48575 230085 48609 230113
rect 48637 230085 48671 230113
rect 48699 230085 48747 230113
rect 48437 230051 48747 230085
rect 48437 230023 48485 230051
rect 48513 230023 48547 230051
rect 48575 230023 48609 230051
rect 48637 230023 48671 230051
rect 48699 230023 48747 230051
rect 48437 229989 48747 230023
rect 48437 229961 48485 229989
rect 48513 229961 48547 229989
rect 48575 229961 48609 229989
rect 48637 229961 48671 229989
rect 48699 229961 48747 229989
rect 48437 221175 48747 229961
rect 59904 230175 60064 230192
rect 59904 230147 59939 230175
rect 59967 230147 60001 230175
rect 60029 230147 60064 230175
rect 59904 230113 60064 230147
rect 59904 230085 59939 230113
rect 59967 230085 60001 230113
rect 60029 230085 60064 230113
rect 59904 230051 60064 230085
rect 59904 230023 59939 230051
rect 59967 230023 60001 230051
rect 60029 230023 60064 230051
rect 59904 229989 60064 230023
rect 59904 229961 59939 229989
rect 59967 229961 60001 229989
rect 60029 229961 60064 229989
rect 59904 229944 60064 229961
rect 75264 230175 75424 230192
rect 75264 230147 75299 230175
rect 75327 230147 75361 230175
rect 75389 230147 75424 230175
rect 75264 230113 75424 230147
rect 75264 230085 75299 230113
rect 75327 230085 75361 230113
rect 75389 230085 75424 230113
rect 75264 230051 75424 230085
rect 75264 230023 75299 230051
rect 75327 230023 75361 230051
rect 75389 230023 75424 230051
rect 75264 229989 75424 230023
rect 75264 229961 75299 229989
rect 75327 229961 75361 229989
rect 75389 229961 75424 229989
rect 75264 229944 75424 229961
rect 90624 230175 90784 230192
rect 90624 230147 90659 230175
rect 90687 230147 90721 230175
rect 90749 230147 90784 230175
rect 90624 230113 90784 230147
rect 90624 230085 90659 230113
rect 90687 230085 90721 230113
rect 90749 230085 90784 230113
rect 90624 230051 90784 230085
rect 90624 230023 90659 230051
rect 90687 230023 90721 230051
rect 90749 230023 90784 230051
rect 90624 229989 90784 230023
rect 90624 229961 90659 229989
rect 90687 229961 90721 229989
rect 90749 229961 90784 229989
rect 90624 229944 90784 229961
rect 105984 230175 106144 230192
rect 105984 230147 106019 230175
rect 106047 230147 106081 230175
rect 106109 230147 106144 230175
rect 105984 230113 106144 230147
rect 105984 230085 106019 230113
rect 106047 230085 106081 230113
rect 106109 230085 106144 230113
rect 105984 230051 106144 230085
rect 105984 230023 106019 230051
rect 106047 230023 106081 230051
rect 106109 230023 106144 230051
rect 105984 229989 106144 230023
rect 105984 229961 106019 229989
rect 106047 229961 106081 229989
rect 106109 229961 106144 229989
rect 105984 229944 106144 229961
rect 121344 230175 121504 230192
rect 121344 230147 121379 230175
rect 121407 230147 121441 230175
rect 121469 230147 121504 230175
rect 121344 230113 121504 230147
rect 121344 230085 121379 230113
rect 121407 230085 121441 230113
rect 121469 230085 121504 230113
rect 121344 230051 121504 230085
rect 121344 230023 121379 230051
rect 121407 230023 121441 230051
rect 121469 230023 121504 230051
rect 121344 229989 121504 230023
rect 121344 229961 121379 229989
rect 121407 229961 121441 229989
rect 121469 229961 121504 229989
rect 121344 229944 121504 229961
rect 136704 230175 136864 230192
rect 136704 230147 136739 230175
rect 136767 230147 136801 230175
rect 136829 230147 136864 230175
rect 136704 230113 136864 230147
rect 136704 230085 136739 230113
rect 136767 230085 136801 230113
rect 136829 230085 136864 230113
rect 136704 230051 136864 230085
rect 136704 230023 136739 230051
rect 136767 230023 136801 230051
rect 136829 230023 136864 230051
rect 136704 229989 136864 230023
rect 136704 229961 136739 229989
rect 136767 229961 136801 229989
rect 136829 229961 136864 229989
rect 136704 229944 136864 229961
rect 52224 227175 52384 227192
rect 52224 227147 52259 227175
rect 52287 227147 52321 227175
rect 52349 227147 52384 227175
rect 52224 227113 52384 227147
rect 52224 227085 52259 227113
rect 52287 227085 52321 227113
rect 52349 227085 52384 227113
rect 52224 227051 52384 227085
rect 52224 227023 52259 227051
rect 52287 227023 52321 227051
rect 52349 227023 52384 227051
rect 52224 226989 52384 227023
rect 52224 226961 52259 226989
rect 52287 226961 52321 226989
rect 52349 226961 52384 226989
rect 52224 226944 52384 226961
rect 67584 227175 67744 227192
rect 67584 227147 67619 227175
rect 67647 227147 67681 227175
rect 67709 227147 67744 227175
rect 67584 227113 67744 227147
rect 67584 227085 67619 227113
rect 67647 227085 67681 227113
rect 67709 227085 67744 227113
rect 67584 227051 67744 227085
rect 67584 227023 67619 227051
rect 67647 227023 67681 227051
rect 67709 227023 67744 227051
rect 67584 226989 67744 227023
rect 67584 226961 67619 226989
rect 67647 226961 67681 226989
rect 67709 226961 67744 226989
rect 67584 226944 67744 226961
rect 82944 227175 83104 227192
rect 82944 227147 82979 227175
rect 83007 227147 83041 227175
rect 83069 227147 83104 227175
rect 82944 227113 83104 227147
rect 82944 227085 82979 227113
rect 83007 227085 83041 227113
rect 83069 227085 83104 227113
rect 82944 227051 83104 227085
rect 82944 227023 82979 227051
rect 83007 227023 83041 227051
rect 83069 227023 83104 227051
rect 82944 226989 83104 227023
rect 82944 226961 82979 226989
rect 83007 226961 83041 226989
rect 83069 226961 83104 226989
rect 82944 226944 83104 226961
rect 98304 227175 98464 227192
rect 98304 227147 98339 227175
rect 98367 227147 98401 227175
rect 98429 227147 98464 227175
rect 98304 227113 98464 227147
rect 98304 227085 98339 227113
rect 98367 227085 98401 227113
rect 98429 227085 98464 227113
rect 98304 227051 98464 227085
rect 98304 227023 98339 227051
rect 98367 227023 98401 227051
rect 98429 227023 98464 227051
rect 98304 226989 98464 227023
rect 98304 226961 98339 226989
rect 98367 226961 98401 226989
rect 98429 226961 98464 226989
rect 98304 226944 98464 226961
rect 113664 227175 113824 227192
rect 113664 227147 113699 227175
rect 113727 227147 113761 227175
rect 113789 227147 113824 227175
rect 113664 227113 113824 227147
rect 113664 227085 113699 227113
rect 113727 227085 113761 227113
rect 113789 227085 113824 227113
rect 113664 227051 113824 227085
rect 113664 227023 113699 227051
rect 113727 227023 113761 227051
rect 113789 227023 113824 227051
rect 113664 226989 113824 227023
rect 113664 226961 113699 226989
rect 113727 226961 113761 226989
rect 113789 226961 113824 226989
rect 113664 226944 113824 226961
rect 129024 227175 129184 227192
rect 129024 227147 129059 227175
rect 129087 227147 129121 227175
rect 129149 227147 129184 227175
rect 129024 227113 129184 227147
rect 129024 227085 129059 227113
rect 129087 227085 129121 227113
rect 129149 227085 129184 227113
rect 129024 227051 129184 227085
rect 129024 227023 129059 227051
rect 129087 227023 129121 227051
rect 129149 227023 129184 227051
rect 129024 226989 129184 227023
rect 129024 226961 129059 226989
rect 129087 226961 129121 226989
rect 129149 226961 129184 226989
rect 129024 226944 129184 226961
rect 144384 227175 144544 227192
rect 144384 227147 144419 227175
rect 144447 227147 144481 227175
rect 144509 227147 144544 227175
rect 144384 227113 144544 227147
rect 144384 227085 144419 227113
rect 144447 227085 144481 227113
rect 144509 227085 144544 227113
rect 144384 227051 144544 227085
rect 144384 227023 144419 227051
rect 144447 227023 144481 227051
rect 144509 227023 144544 227051
rect 144384 226989 144544 227023
rect 144384 226961 144419 226989
rect 144447 226961 144481 226989
rect 144509 226961 144544 226989
rect 144384 226944 144544 226961
rect 154577 227175 154887 235961
rect 154577 227147 154625 227175
rect 154653 227147 154687 227175
rect 154715 227147 154749 227175
rect 154777 227147 154811 227175
rect 154839 227147 154887 227175
rect 154577 227113 154887 227147
rect 154577 227085 154625 227113
rect 154653 227085 154687 227113
rect 154715 227085 154749 227113
rect 154777 227085 154811 227113
rect 154839 227085 154887 227113
rect 154577 227051 154887 227085
rect 154577 227023 154625 227051
rect 154653 227023 154687 227051
rect 154715 227023 154749 227051
rect 154777 227023 154811 227051
rect 154839 227023 154887 227051
rect 154577 226989 154887 227023
rect 154577 226961 154625 226989
rect 154653 226961 154687 226989
rect 154715 226961 154749 226989
rect 154777 226961 154811 226989
rect 154839 226961 154887 226989
rect 48437 221147 48485 221175
rect 48513 221147 48547 221175
rect 48575 221147 48609 221175
rect 48637 221147 48671 221175
rect 48699 221147 48747 221175
rect 48437 221113 48747 221147
rect 48437 221085 48485 221113
rect 48513 221085 48547 221113
rect 48575 221085 48609 221113
rect 48637 221085 48671 221113
rect 48699 221085 48747 221113
rect 48437 221051 48747 221085
rect 48437 221023 48485 221051
rect 48513 221023 48547 221051
rect 48575 221023 48609 221051
rect 48637 221023 48671 221051
rect 48699 221023 48747 221051
rect 48437 220989 48747 221023
rect 48437 220961 48485 220989
rect 48513 220961 48547 220989
rect 48575 220961 48609 220989
rect 48637 220961 48671 220989
rect 48699 220961 48747 220989
rect 48437 212175 48747 220961
rect 59904 221175 60064 221192
rect 59904 221147 59939 221175
rect 59967 221147 60001 221175
rect 60029 221147 60064 221175
rect 59904 221113 60064 221147
rect 59904 221085 59939 221113
rect 59967 221085 60001 221113
rect 60029 221085 60064 221113
rect 59904 221051 60064 221085
rect 59904 221023 59939 221051
rect 59967 221023 60001 221051
rect 60029 221023 60064 221051
rect 59904 220989 60064 221023
rect 59904 220961 59939 220989
rect 59967 220961 60001 220989
rect 60029 220961 60064 220989
rect 59904 220944 60064 220961
rect 75264 221175 75424 221192
rect 75264 221147 75299 221175
rect 75327 221147 75361 221175
rect 75389 221147 75424 221175
rect 75264 221113 75424 221147
rect 75264 221085 75299 221113
rect 75327 221085 75361 221113
rect 75389 221085 75424 221113
rect 75264 221051 75424 221085
rect 75264 221023 75299 221051
rect 75327 221023 75361 221051
rect 75389 221023 75424 221051
rect 75264 220989 75424 221023
rect 75264 220961 75299 220989
rect 75327 220961 75361 220989
rect 75389 220961 75424 220989
rect 75264 220944 75424 220961
rect 90624 221175 90784 221192
rect 90624 221147 90659 221175
rect 90687 221147 90721 221175
rect 90749 221147 90784 221175
rect 90624 221113 90784 221147
rect 90624 221085 90659 221113
rect 90687 221085 90721 221113
rect 90749 221085 90784 221113
rect 90624 221051 90784 221085
rect 90624 221023 90659 221051
rect 90687 221023 90721 221051
rect 90749 221023 90784 221051
rect 90624 220989 90784 221023
rect 90624 220961 90659 220989
rect 90687 220961 90721 220989
rect 90749 220961 90784 220989
rect 90624 220944 90784 220961
rect 105984 221175 106144 221192
rect 105984 221147 106019 221175
rect 106047 221147 106081 221175
rect 106109 221147 106144 221175
rect 105984 221113 106144 221147
rect 105984 221085 106019 221113
rect 106047 221085 106081 221113
rect 106109 221085 106144 221113
rect 105984 221051 106144 221085
rect 105984 221023 106019 221051
rect 106047 221023 106081 221051
rect 106109 221023 106144 221051
rect 105984 220989 106144 221023
rect 105984 220961 106019 220989
rect 106047 220961 106081 220989
rect 106109 220961 106144 220989
rect 105984 220944 106144 220961
rect 121344 221175 121504 221192
rect 121344 221147 121379 221175
rect 121407 221147 121441 221175
rect 121469 221147 121504 221175
rect 121344 221113 121504 221147
rect 121344 221085 121379 221113
rect 121407 221085 121441 221113
rect 121469 221085 121504 221113
rect 121344 221051 121504 221085
rect 121344 221023 121379 221051
rect 121407 221023 121441 221051
rect 121469 221023 121504 221051
rect 121344 220989 121504 221023
rect 121344 220961 121379 220989
rect 121407 220961 121441 220989
rect 121469 220961 121504 220989
rect 121344 220944 121504 220961
rect 136704 221175 136864 221192
rect 136704 221147 136739 221175
rect 136767 221147 136801 221175
rect 136829 221147 136864 221175
rect 136704 221113 136864 221147
rect 136704 221085 136739 221113
rect 136767 221085 136801 221113
rect 136829 221085 136864 221113
rect 136704 221051 136864 221085
rect 136704 221023 136739 221051
rect 136767 221023 136801 221051
rect 136829 221023 136864 221051
rect 136704 220989 136864 221023
rect 136704 220961 136739 220989
rect 136767 220961 136801 220989
rect 136829 220961 136864 220989
rect 136704 220944 136864 220961
rect 52224 218175 52384 218192
rect 52224 218147 52259 218175
rect 52287 218147 52321 218175
rect 52349 218147 52384 218175
rect 52224 218113 52384 218147
rect 52224 218085 52259 218113
rect 52287 218085 52321 218113
rect 52349 218085 52384 218113
rect 52224 218051 52384 218085
rect 52224 218023 52259 218051
rect 52287 218023 52321 218051
rect 52349 218023 52384 218051
rect 52224 217989 52384 218023
rect 52224 217961 52259 217989
rect 52287 217961 52321 217989
rect 52349 217961 52384 217989
rect 52224 217944 52384 217961
rect 67584 218175 67744 218192
rect 67584 218147 67619 218175
rect 67647 218147 67681 218175
rect 67709 218147 67744 218175
rect 67584 218113 67744 218147
rect 67584 218085 67619 218113
rect 67647 218085 67681 218113
rect 67709 218085 67744 218113
rect 67584 218051 67744 218085
rect 67584 218023 67619 218051
rect 67647 218023 67681 218051
rect 67709 218023 67744 218051
rect 67584 217989 67744 218023
rect 67584 217961 67619 217989
rect 67647 217961 67681 217989
rect 67709 217961 67744 217989
rect 67584 217944 67744 217961
rect 82944 218175 83104 218192
rect 82944 218147 82979 218175
rect 83007 218147 83041 218175
rect 83069 218147 83104 218175
rect 82944 218113 83104 218147
rect 82944 218085 82979 218113
rect 83007 218085 83041 218113
rect 83069 218085 83104 218113
rect 82944 218051 83104 218085
rect 82944 218023 82979 218051
rect 83007 218023 83041 218051
rect 83069 218023 83104 218051
rect 82944 217989 83104 218023
rect 82944 217961 82979 217989
rect 83007 217961 83041 217989
rect 83069 217961 83104 217989
rect 82944 217944 83104 217961
rect 98304 218175 98464 218192
rect 98304 218147 98339 218175
rect 98367 218147 98401 218175
rect 98429 218147 98464 218175
rect 98304 218113 98464 218147
rect 98304 218085 98339 218113
rect 98367 218085 98401 218113
rect 98429 218085 98464 218113
rect 98304 218051 98464 218085
rect 98304 218023 98339 218051
rect 98367 218023 98401 218051
rect 98429 218023 98464 218051
rect 98304 217989 98464 218023
rect 98304 217961 98339 217989
rect 98367 217961 98401 217989
rect 98429 217961 98464 217989
rect 98304 217944 98464 217961
rect 113664 218175 113824 218192
rect 113664 218147 113699 218175
rect 113727 218147 113761 218175
rect 113789 218147 113824 218175
rect 113664 218113 113824 218147
rect 113664 218085 113699 218113
rect 113727 218085 113761 218113
rect 113789 218085 113824 218113
rect 113664 218051 113824 218085
rect 113664 218023 113699 218051
rect 113727 218023 113761 218051
rect 113789 218023 113824 218051
rect 113664 217989 113824 218023
rect 113664 217961 113699 217989
rect 113727 217961 113761 217989
rect 113789 217961 113824 217989
rect 113664 217944 113824 217961
rect 129024 218175 129184 218192
rect 129024 218147 129059 218175
rect 129087 218147 129121 218175
rect 129149 218147 129184 218175
rect 129024 218113 129184 218147
rect 129024 218085 129059 218113
rect 129087 218085 129121 218113
rect 129149 218085 129184 218113
rect 129024 218051 129184 218085
rect 129024 218023 129059 218051
rect 129087 218023 129121 218051
rect 129149 218023 129184 218051
rect 129024 217989 129184 218023
rect 129024 217961 129059 217989
rect 129087 217961 129121 217989
rect 129149 217961 129184 217989
rect 129024 217944 129184 217961
rect 144384 218175 144544 218192
rect 144384 218147 144419 218175
rect 144447 218147 144481 218175
rect 144509 218147 144544 218175
rect 144384 218113 144544 218147
rect 144384 218085 144419 218113
rect 144447 218085 144481 218113
rect 144509 218085 144544 218113
rect 144384 218051 144544 218085
rect 144384 218023 144419 218051
rect 144447 218023 144481 218051
rect 144509 218023 144544 218051
rect 144384 217989 144544 218023
rect 144384 217961 144419 217989
rect 144447 217961 144481 217989
rect 144509 217961 144544 217989
rect 144384 217944 144544 217961
rect 154577 218175 154887 226961
rect 154577 218147 154625 218175
rect 154653 218147 154687 218175
rect 154715 218147 154749 218175
rect 154777 218147 154811 218175
rect 154839 218147 154887 218175
rect 154577 218113 154887 218147
rect 154577 218085 154625 218113
rect 154653 218085 154687 218113
rect 154715 218085 154749 218113
rect 154777 218085 154811 218113
rect 154839 218085 154887 218113
rect 154577 218051 154887 218085
rect 154577 218023 154625 218051
rect 154653 218023 154687 218051
rect 154715 218023 154749 218051
rect 154777 218023 154811 218051
rect 154839 218023 154887 218051
rect 154577 217989 154887 218023
rect 154577 217961 154625 217989
rect 154653 217961 154687 217989
rect 154715 217961 154749 217989
rect 154777 217961 154811 217989
rect 154839 217961 154887 217989
rect 48437 212147 48485 212175
rect 48513 212147 48547 212175
rect 48575 212147 48609 212175
rect 48637 212147 48671 212175
rect 48699 212147 48747 212175
rect 48437 212113 48747 212147
rect 48437 212085 48485 212113
rect 48513 212085 48547 212113
rect 48575 212085 48609 212113
rect 48637 212085 48671 212113
rect 48699 212085 48747 212113
rect 48437 212051 48747 212085
rect 48437 212023 48485 212051
rect 48513 212023 48547 212051
rect 48575 212023 48609 212051
rect 48637 212023 48671 212051
rect 48699 212023 48747 212051
rect 48437 211989 48747 212023
rect 48437 211961 48485 211989
rect 48513 211961 48547 211989
rect 48575 211961 48609 211989
rect 48637 211961 48671 211989
rect 48699 211961 48747 211989
rect 48437 203175 48747 211961
rect 59904 212175 60064 212192
rect 59904 212147 59939 212175
rect 59967 212147 60001 212175
rect 60029 212147 60064 212175
rect 59904 212113 60064 212147
rect 59904 212085 59939 212113
rect 59967 212085 60001 212113
rect 60029 212085 60064 212113
rect 59904 212051 60064 212085
rect 59904 212023 59939 212051
rect 59967 212023 60001 212051
rect 60029 212023 60064 212051
rect 59904 211989 60064 212023
rect 59904 211961 59939 211989
rect 59967 211961 60001 211989
rect 60029 211961 60064 211989
rect 59904 211944 60064 211961
rect 75264 212175 75424 212192
rect 75264 212147 75299 212175
rect 75327 212147 75361 212175
rect 75389 212147 75424 212175
rect 75264 212113 75424 212147
rect 75264 212085 75299 212113
rect 75327 212085 75361 212113
rect 75389 212085 75424 212113
rect 75264 212051 75424 212085
rect 75264 212023 75299 212051
rect 75327 212023 75361 212051
rect 75389 212023 75424 212051
rect 75264 211989 75424 212023
rect 75264 211961 75299 211989
rect 75327 211961 75361 211989
rect 75389 211961 75424 211989
rect 75264 211944 75424 211961
rect 90624 212175 90784 212192
rect 90624 212147 90659 212175
rect 90687 212147 90721 212175
rect 90749 212147 90784 212175
rect 90624 212113 90784 212147
rect 90624 212085 90659 212113
rect 90687 212085 90721 212113
rect 90749 212085 90784 212113
rect 90624 212051 90784 212085
rect 90624 212023 90659 212051
rect 90687 212023 90721 212051
rect 90749 212023 90784 212051
rect 90624 211989 90784 212023
rect 90624 211961 90659 211989
rect 90687 211961 90721 211989
rect 90749 211961 90784 211989
rect 90624 211944 90784 211961
rect 105984 212175 106144 212192
rect 105984 212147 106019 212175
rect 106047 212147 106081 212175
rect 106109 212147 106144 212175
rect 105984 212113 106144 212147
rect 105984 212085 106019 212113
rect 106047 212085 106081 212113
rect 106109 212085 106144 212113
rect 105984 212051 106144 212085
rect 105984 212023 106019 212051
rect 106047 212023 106081 212051
rect 106109 212023 106144 212051
rect 105984 211989 106144 212023
rect 105984 211961 106019 211989
rect 106047 211961 106081 211989
rect 106109 211961 106144 211989
rect 105984 211944 106144 211961
rect 121344 212175 121504 212192
rect 121344 212147 121379 212175
rect 121407 212147 121441 212175
rect 121469 212147 121504 212175
rect 121344 212113 121504 212147
rect 121344 212085 121379 212113
rect 121407 212085 121441 212113
rect 121469 212085 121504 212113
rect 121344 212051 121504 212085
rect 121344 212023 121379 212051
rect 121407 212023 121441 212051
rect 121469 212023 121504 212051
rect 121344 211989 121504 212023
rect 121344 211961 121379 211989
rect 121407 211961 121441 211989
rect 121469 211961 121504 211989
rect 121344 211944 121504 211961
rect 136704 212175 136864 212192
rect 136704 212147 136739 212175
rect 136767 212147 136801 212175
rect 136829 212147 136864 212175
rect 136704 212113 136864 212147
rect 136704 212085 136739 212113
rect 136767 212085 136801 212113
rect 136829 212085 136864 212113
rect 136704 212051 136864 212085
rect 136704 212023 136739 212051
rect 136767 212023 136801 212051
rect 136829 212023 136864 212051
rect 136704 211989 136864 212023
rect 136704 211961 136739 211989
rect 136767 211961 136801 211989
rect 136829 211961 136864 211989
rect 136704 211944 136864 211961
rect 52224 209175 52384 209192
rect 52224 209147 52259 209175
rect 52287 209147 52321 209175
rect 52349 209147 52384 209175
rect 52224 209113 52384 209147
rect 52224 209085 52259 209113
rect 52287 209085 52321 209113
rect 52349 209085 52384 209113
rect 52224 209051 52384 209085
rect 52224 209023 52259 209051
rect 52287 209023 52321 209051
rect 52349 209023 52384 209051
rect 52224 208989 52384 209023
rect 52224 208961 52259 208989
rect 52287 208961 52321 208989
rect 52349 208961 52384 208989
rect 52224 208944 52384 208961
rect 67584 209175 67744 209192
rect 67584 209147 67619 209175
rect 67647 209147 67681 209175
rect 67709 209147 67744 209175
rect 67584 209113 67744 209147
rect 67584 209085 67619 209113
rect 67647 209085 67681 209113
rect 67709 209085 67744 209113
rect 67584 209051 67744 209085
rect 67584 209023 67619 209051
rect 67647 209023 67681 209051
rect 67709 209023 67744 209051
rect 67584 208989 67744 209023
rect 67584 208961 67619 208989
rect 67647 208961 67681 208989
rect 67709 208961 67744 208989
rect 67584 208944 67744 208961
rect 82944 209175 83104 209192
rect 82944 209147 82979 209175
rect 83007 209147 83041 209175
rect 83069 209147 83104 209175
rect 82944 209113 83104 209147
rect 82944 209085 82979 209113
rect 83007 209085 83041 209113
rect 83069 209085 83104 209113
rect 82944 209051 83104 209085
rect 82944 209023 82979 209051
rect 83007 209023 83041 209051
rect 83069 209023 83104 209051
rect 82944 208989 83104 209023
rect 82944 208961 82979 208989
rect 83007 208961 83041 208989
rect 83069 208961 83104 208989
rect 82944 208944 83104 208961
rect 98304 209175 98464 209192
rect 98304 209147 98339 209175
rect 98367 209147 98401 209175
rect 98429 209147 98464 209175
rect 98304 209113 98464 209147
rect 98304 209085 98339 209113
rect 98367 209085 98401 209113
rect 98429 209085 98464 209113
rect 98304 209051 98464 209085
rect 98304 209023 98339 209051
rect 98367 209023 98401 209051
rect 98429 209023 98464 209051
rect 98304 208989 98464 209023
rect 98304 208961 98339 208989
rect 98367 208961 98401 208989
rect 98429 208961 98464 208989
rect 98304 208944 98464 208961
rect 113664 209175 113824 209192
rect 113664 209147 113699 209175
rect 113727 209147 113761 209175
rect 113789 209147 113824 209175
rect 113664 209113 113824 209147
rect 113664 209085 113699 209113
rect 113727 209085 113761 209113
rect 113789 209085 113824 209113
rect 113664 209051 113824 209085
rect 113664 209023 113699 209051
rect 113727 209023 113761 209051
rect 113789 209023 113824 209051
rect 113664 208989 113824 209023
rect 113664 208961 113699 208989
rect 113727 208961 113761 208989
rect 113789 208961 113824 208989
rect 113664 208944 113824 208961
rect 129024 209175 129184 209192
rect 129024 209147 129059 209175
rect 129087 209147 129121 209175
rect 129149 209147 129184 209175
rect 129024 209113 129184 209147
rect 129024 209085 129059 209113
rect 129087 209085 129121 209113
rect 129149 209085 129184 209113
rect 129024 209051 129184 209085
rect 129024 209023 129059 209051
rect 129087 209023 129121 209051
rect 129149 209023 129184 209051
rect 129024 208989 129184 209023
rect 129024 208961 129059 208989
rect 129087 208961 129121 208989
rect 129149 208961 129184 208989
rect 129024 208944 129184 208961
rect 144384 209175 144544 209192
rect 144384 209147 144419 209175
rect 144447 209147 144481 209175
rect 144509 209147 144544 209175
rect 144384 209113 144544 209147
rect 144384 209085 144419 209113
rect 144447 209085 144481 209113
rect 144509 209085 144544 209113
rect 144384 209051 144544 209085
rect 144384 209023 144419 209051
rect 144447 209023 144481 209051
rect 144509 209023 144544 209051
rect 144384 208989 144544 209023
rect 144384 208961 144419 208989
rect 144447 208961 144481 208989
rect 144509 208961 144544 208989
rect 144384 208944 144544 208961
rect 154577 209175 154887 217961
rect 154577 209147 154625 209175
rect 154653 209147 154687 209175
rect 154715 209147 154749 209175
rect 154777 209147 154811 209175
rect 154839 209147 154887 209175
rect 154577 209113 154887 209147
rect 154577 209085 154625 209113
rect 154653 209085 154687 209113
rect 154715 209085 154749 209113
rect 154777 209085 154811 209113
rect 154839 209085 154887 209113
rect 154577 209051 154887 209085
rect 154577 209023 154625 209051
rect 154653 209023 154687 209051
rect 154715 209023 154749 209051
rect 154777 209023 154811 209051
rect 154839 209023 154887 209051
rect 154577 208989 154887 209023
rect 154577 208961 154625 208989
rect 154653 208961 154687 208989
rect 154715 208961 154749 208989
rect 154777 208961 154811 208989
rect 154839 208961 154887 208989
rect 48437 203147 48485 203175
rect 48513 203147 48547 203175
rect 48575 203147 48609 203175
rect 48637 203147 48671 203175
rect 48699 203147 48747 203175
rect 48437 203113 48747 203147
rect 48437 203085 48485 203113
rect 48513 203085 48547 203113
rect 48575 203085 48609 203113
rect 48637 203085 48671 203113
rect 48699 203085 48747 203113
rect 48437 203051 48747 203085
rect 48437 203023 48485 203051
rect 48513 203023 48547 203051
rect 48575 203023 48609 203051
rect 48637 203023 48671 203051
rect 48699 203023 48747 203051
rect 48437 202989 48747 203023
rect 48437 202961 48485 202989
rect 48513 202961 48547 202989
rect 48575 202961 48609 202989
rect 48637 202961 48671 202989
rect 48699 202961 48747 202989
rect 48437 194175 48747 202961
rect 59904 203175 60064 203192
rect 59904 203147 59939 203175
rect 59967 203147 60001 203175
rect 60029 203147 60064 203175
rect 59904 203113 60064 203147
rect 59904 203085 59939 203113
rect 59967 203085 60001 203113
rect 60029 203085 60064 203113
rect 59904 203051 60064 203085
rect 59904 203023 59939 203051
rect 59967 203023 60001 203051
rect 60029 203023 60064 203051
rect 59904 202989 60064 203023
rect 59904 202961 59939 202989
rect 59967 202961 60001 202989
rect 60029 202961 60064 202989
rect 59904 202944 60064 202961
rect 75264 203175 75424 203192
rect 75264 203147 75299 203175
rect 75327 203147 75361 203175
rect 75389 203147 75424 203175
rect 75264 203113 75424 203147
rect 75264 203085 75299 203113
rect 75327 203085 75361 203113
rect 75389 203085 75424 203113
rect 75264 203051 75424 203085
rect 75264 203023 75299 203051
rect 75327 203023 75361 203051
rect 75389 203023 75424 203051
rect 75264 202989 75424 203023
rect 75264 202961 75299 202989
rect 75327 202961 75361 202989
rect 75389 202961 75424 202989
rect 75264 202944 75424 202961
rect 90624 203175 90784 203192
rect 90624 203147 90659 203175
rect 90687 203147 90721 203175
rect 90749 203147 90784 203175
rect 90624 203113 90784 203147
rect 90624 203085 90659 203113
rect 90687 203085 90721 203113
rect 90749 203085 90784 203113
rect 90624 203051 90784 203085
rect 90624 203023 90659 203051
rect 90687 203023 90721 203051
rect 90749 203023 90784 203051
rect 90624 202989 90784 203023
rect 90624 202961 90659 202989
rect 90687 202961 90721 202989
rect 90749 202961 90784 202989
rect 90624 202944 90784 202961
rect 105984 203175 106144 203192
rect 105984 203147 106019 203175
rect 106047 203147 106081 203175
rect 106109 203147 106144 203175
rect 105984 203113 106144 203147
rect 105984 203085 106019 203113
rect 106047 203085 106081 203113
rect 106109 203085 106144 203113
rect 105984 203051 106144 203085
rect 105984 203023 106019 203051
rect 106047 203023 106081 203051
rect 106109 203023 106144 203051
rect 105984 202989 106144 203023
rect 105984 202961 106019 202989
rect 106047 202961 106081 202989
rect 106109 202961 106144 202989
rect 105984 202944 106144 202961
rect 121344 203175 121504 203192
rect 121344 203147 121379 203175
rect 121407 203147 121441 203175
rect 121469 203147 121504 203175
rect 121344 203113 121504 203147
rect 121344 203085 121379 203113
rect 121407 203085 121441 203113
rect 121469 203085 121504 203113
rect 121344 203051 121504 203085
rect 121344 203023 121379 203051
rect 121407 203023 121441 203051
rect 121469 203023 121504 203051
rect 121344 202989 121504 203023
rect 121344 202961 121379 202989
rect 121407 202961 121441 202989
rect 121469 202961 121504 202989
rect 121344 202944 121504 202961
rect 136704 203175 136864 203192
rect 136704 203147 136739 203175
rect 136767 203147 136801 203175
rect 136829 203147 136864 203175
rect 136704 203113 136864 203147
rect 136704 203085 136739 203113
rect 136767 203085 136801 203113
rect 136829 203085 136864 203113
rect 136704 203051 136864 203085
rect 136704 203023 136739 203051
rect 136767 203023 136801 203051
rect 136829 203023 136864 203051
rect 136704 202989 136864 203023
rect 136704 202961 136739 202989
rect 136767 202961 136801 202989
rect 136829 202961 136864 202989
rect 136704 202944 136864 202961
rect 154577 200175 154887 208961
rect 154577 200147 154625 200175
rect 154653 200147 154687 200175
rect 154715 200147 154749 200175
rect 154777 200147 154811 200175
rect 154839 200147 154887 200175
rect 154577 200113 154887 200147
rect 154577 200085 154625 200113
rect 154653 200085 154687 200113
rect 154715 200085 154749 200113
rect 154777 200085 154811 200113
rect 154839 200085 154887 200113
rect 154577 200051 154887 200085
rect 154577 200023 154625 200051
rect 154653 200023 154687 200051
rect 154715 200023 154749 200051
rect 154777 200023 154811 200051
rect 154839 200023 154887 200051
rect 154577 199989 154887 200023
rect 154577 199961 154625 199989
rect 154653 199961 154687 199989
rect 154715 199961 154749 199989
rect 154777 199961 154811 199989
rect 154839 199961 154887 199989
rect 48437 194147 48485 194175
rect 48513 194147 48547 194175
rect 48575 194147 48609 194175
rect 48637 194147 48671 194175
rect 48699 194147 48747 194175
rect 48437 194113 48747 194147
rect 48437 194085 48485 194113
rect 48513 194085 48547 194113
rect 48575 194085 48609 194113
rect 48637 194085 48671 194113
rect 48699 194085 48747 194113
rect 48437 194051 48747 194085
rect 48437 194023 48485 194051
rect 48513 194023 48547 194051
rect 48575 194023 48609 194051
rect 48637 194023 48671 194051
rect 48699 194023 48747 194051
rect 48437 193989 48747 194023
rect 48437 193961 48485 193989
rect 48513 193961 48547 193989
rect 48575 193961 48609 193989
rect 48637 193961 48671 193989
rect 48699 193961 48747 193989
rect 48437 185175 48747 193961
rect 48437 185147 48485 185175
rect 48513 185147 48547 185175
rect 48575 185147 48609 185175
rect 48637 185147 48671 185175
rect 48699 185147 48747 185175
rect 48437 185113 48747 185147
rect 48437 185085 48485 185113
rect 48513 185085 48547 185113
rect 48575 185085 48609 185113
rect 48637 185085 48671 185113
rect 48699 185085 48747 185113
rect 48437 185051 48747 185085
rect 48437 185023 48485 185051
rect 48513 185023 48547 185051
rect 48575 185023 48609 185051
rect 48637 185023 48671 185051
rect 48699 185023 48747 185051
rect 48437 184989 48747 185023
rect 48437 184961 48485 184989
rect 48513 184961 48547 184989
rect 48575 184961 48609 184989
rect 48637 184961 48671 184989
rect 48699 184961 48747 184989
rect 48437 176175 48747 184961
rect 57437 194175 57747 199205
rect 57437 194147 57485 194175
rect 57513 194147 57547 194175
rect 57575 194147 57609 194175
rect 57637 194147 57671 194175
rect 57699 194147 57747 194175
rect 57437 194113 57747 194147
rect 57437 194085 57485 194113
rect 57513 194085 57547 194113
rect 57575 194085 57609 194113
rect 57637 194085 57671 194113
rect 57699 194085 57747 194113
rect 57437 194051 57747 194085
rect 57437 194023 57485 194051
rect 57513 194023 57547 194051
rect 57575 194023 57609 194051
rect 57637 194023 57671 194051
rect 57699 194023 57747 194051
rect 57437 193989 57747 194023
rect 57437 193961 57485 193989
rect 57513 193961 57547 193989
rect 57575 193961 57609 193989
rect 57637 193961 57671 193989
rect 57699 193961 57747 193989
rect 57437 185175 57747 193961
rect 57437 185147 57485 185175
rect 57513 185147 57547 185175
rect 57575 185147 57609 185175
rect 57637 185147 57671 185175
rect 57699 185147 57747 185175
rect 57437 185113 57747 185147
rect 57437 185085 57485 185113
rect 57513 185085 57547 185113
rect 57575 185085 57609 185113
rect 57637 185085 57671 185113
rect 57699 185085 57747 185113
rect 57437 185051 57747 185085
rect 57437 185023 57485 185051
rect 57513 185023 57547 185051
rect 57575 185023 57609 185051
rect 57637 185023 57671 185051
rect 57699 185023 57747 185051
rect 57437 184989 57747 185023
rect 57437 184961 57485 184989
rect 57513 184961 57547 184989
rect 57575 184961 57609 184989
rect 57637 184961 57671 184989
rect 57699 184961 57747 184989
rect 57437 182635 57747 184961
rect 66437 194175 66747 199205
rect 66437 194147 66485 194175
rect 66513 194147 66547 194175
rect 66575 194147 66609 194175
rect 66637 194147 66671 194175
rect 66699 194147 66747 194175
rect 66437 194113 66747 194147
rect 66437 194085 66485 194113
rect 66513 194085 66547 194113
rect 66575 194085 66609 194113
rect 66637 194085 66671 194113
rect 66699 194085 66747 194113
rect 66437 194051 66747 194085
rect 66437 194023 66485 194051
rect 66513 194023 66547 194051
rect 66575 194023 66609 194051
rect 66637 194023 66671 194051
rect 66699 194023 66747 194051
rect 66437 193989 66747 194023
rect 66437 193961 66485 193989
rect 66513 193961 66547 193989
rect 66575 193961 66609 193989
rect 66637 193961 66671 193989
rect 66699 193961 66747 193989
rect 66437 185175 66747 193961
rect 66437 185147 66485 185175
rect 66513 185147 66547 185175
rect 66575 185147 66609 185175
rect 66637 185147 66671 185175
rect 66699 185147 66747 185175
rect 66437 185113 66747 185147
rect 66437 185085 66485 185113
rect 66513 185085 66547 185113
rect 66575 185085 66609 185113
rect 66637 185085 66671 185113
rect 66699 185085 66747 185113
rect 66437 185051 66747 185085
rect 66437 185023 66485 185051
rect 66513 185023 66547 185051
rect 66575 185023 66609 185051
rect 66637 185023 66671 185051
rect 66699 185023 66747 185051
rect 66437 184989 66747 185023
rect 66437 184961 66485 184989
rect 66513 184961 66547 184989
rect 66575 184961 66609 184989
rect 66637 184961 66671 184989
rect 66699 184961 66747 184989
rect 66437 182635 66747 184961
rect 75437 194175 75747 199205
rect 75437 194147 75485 194175
rect 75513 194147 75547 194175
rect 75575 194147 75609 194175
rect 75637 194147 75671 194175
rect 75699 194147 75747 194175
rect 75437 194113 75747 194147
rect 75437 194085 75485 194113
rect 75513 194085 75547 194113
rect 75575 194085 75609 194113
rect 75637 194085 75671 194113
rect 75699 194085 75747 194113
rect 75437 194051 75747 194085
rect 75437 194023 75485 194051
rect 75513 194023 75547 194051
rect 75575 194023 75609 194051
rect 75637 194023 75671 194051
rect 75699 194023 75747 194051
rect 75437 193989 75747 194023
rect 75437 193961 75485 193989
rect 75513 193961 75547 193989
rect 75575 193961 75609 193989
rect 75637 193961 75671 193989
rect 75699 193961 75747 193989
rect 75437 185175 75747 193961
rect 75437 185147 75485 185175
rect 75513 185147 75547 185175
rect 75575 185147 75609 185175
rect 75637 185147 75671 185175
rect 75699 185147 75747 185175
rect 75437 185113 75747 185147
rect 75437 185085 75485 185113
rect 75513 185085 75547 185113
rect 75575 185085 75609 185113
rect 75637 185085 75671 185113
rect 75699 185085 75747 185113
rect 75437 185051 75747 185085
rect 75437 185023 75485 185051
rect 75513 185023 75547 185051
rect 75575 185023 75609 185051
rect 75637 185023 75671 185051
rect 75699 185023 75747 185051
rect 75437 184989 75747 185023
rect 75437 184961 75485 184989
rect 75513 184961 75547 184989
rect 75575 184961 75609 184989
rect 75637 184961 75671 184989
rect 75699 184961 75747 184989
rect 75437 184466 75747 184961
rect 84437 194175 84747 199205
rect 84437 194147 84485 194175
rect 84513 194147 84547 194175
rect 84575 194147 84609 194175
rect 84637 194147 84671 194175
rect 84699 194147 84747 194175
rect 84437 194113 84747 194147
rect 84437 194085 84485 194113
rect 84513 194085 84547 194113
rect 84575 194085 84609 194113
rect 84637 194085 84671 194113
rect 84699 194085 84747 194113
rect 84437 194051 84747 194085
rect 84437 194023 84485 194051
rect 84513 194023 84547 194051
rect 84575 194023 84609 194051
rect 84637 194023 84671 194051
rect 84699 194023 84747 194051
rect 84437 193989 84747 194023
rect 84437 193961 84485 193989
rect 84513 193961 84547 193989
rect 84575 193961 84609 193989
rect 84637 193961 84671 193989
rect 84699 193961 84747 193989
rect 84437 185175 84747 193961
rect 84437 185147 84485 185175
rect 84513 185147 84547 185175
rect 84575 185147 84609 185175
rect 84637 185147 84671 185175
rect 84699 185147 84747 185175
rect 84437 185113 84747 185147
rect 84437 185085 84485 185113
rect 84513 185085 84547 185113
rect 84575 185085 84609 185113
rect 84637 185085 84671 185113
rect 84699 185085 84747 185113
rect 84437 185051 84747 185085
rect 84437 185023 84485 185051
rect 84513 185023 84547 185051
rect 84575 185023 84609 185051
rect 84637 185023 84671 185051
rect 84699 185023 84747 185051
rect 84437 184989 84747 185023
rect 84437 184961 84485 184989
rect 84513 184961 84547 184989
rect 84575 184961 84609 184989
rect 84637 184961 84671 184989
rect 84699 184961 84747 184989
rect 84437 182635 84747 184961
rect 93437 194175 93747 199205
rect 93437 194147 93485 194175
rect 93513 194147 93547 194175
rect 93575 194147 93609 194175
rect 93637 194147 93671 194175
rect 93699 194147 93747 194175
rect 93437 194113 93747 194147
rect 93437 194085 93485 194113
rect 93513 194085 93547 194113
rect 93575 194085 93609 194113
rect 93637 194085 93671 194113
rect 93699 194085 93747 194113
rect 93437 194051 93747 194085
rect 93437 194023 93485 194051
rect 93513 194023 93547 194051
rect 93575 194023 93609 194051
rect 93637 194023 93671 194051
rect 93699 194023 93747 194051
rect 93437 193989 93747 194023
rect 93437 193961 93485 193989
rect 93513 193961 93547 193989
rect 93575 193961 93609 193989
rect 93637 193961 93671 193989
rect 93699 193961 93747 193989
rect 93437 185175 93747 193961
rect 93437 185147 93485 185175
rect 93513 185147 93547 185175
rect 93575 185147 93609 185175
rect 93637 185147 93671 185175
rect 93699 185147 93747 185175
rect 93437 185113 93747 185147
rect 93437 185085 93485 185113
rect 93513 185085 93547 185113
rect 93575 185085 93609 185113
rect 93637 185085 93671 185113
rect 93699 185085 93747 185113
rect 93437 185051 93747 185085
rect 93437 185023 93485 185051
rect 93513 185023 93547 185051
rect 93575 185023 93609 185051
rect 93637 185023 93671 185051
rect 93699 185023 93747 185051
rect 93437 184989 93747 185023
rect 93437 184961 93485 184989
rect 93513 184961 93547 184989
rect 93575 184961 93609 184989
rect 93637 184961 93671 184989
rect 93699 184961 93747 184989
rect 93437 182635 93747 184961
rect 102437 194175 102747 199205
rect 102437 194147 102485 194175
rect 102513 194147 102547 194175
rect 102575 194147 102609 194175
rect 102637 194147 102671 194175
rect 102699 194147 102747 194175
rect 102437 194113 102747 194147
rect 102437 194085 102485 194113
rect 102513 194085 102547 194113
rect 102575 194085 102609 194113
rect 102637 194085 102671 194113
rect 102699 194085 102747 194113
rect 102437 194051 102747 194085
rect 102437 194023 102485 194051
rect 102513 194023 102547 194051
rect 102575 194023 102609 194051
rect 102637 194023 102671 194051
rect 102699 194023 102747 194051
rect 102437 193989 102747 194023
rect 102437 193961 102485 193989
rect 102513 193961 102547 193989
rect 102575 193961 102609 193989
rect 102637 193961 102671 193989
rect 102699 193961 102747 193989
rect 102437 185175 102747 193961
rect 102437 185147 102485 185175
rect 102513 185147 102547 185175
rect 102575 185147 102609 185175
rect 102637 185147 102671 185175
rect 102699 185147 102747 185175
rect 102437 185113 102747 185147
rect 102437 185085 102485 185113
rect 102513 185085 102547 185113
rect 102575 185085 102609 185113
rect 102637 185085 102671 185113
rect 102699 185085 102747 185113
rect 102437 185051 102747 185085
rect 102437 185023 102485 185051
rect 102513 185023 102547 185051
rect 102575 185023 102609 185051
rect 102637 185023 102671 185051
rect 102699 185023 102747 185051
rect 102437 184989 102747 185023
rect 102437 184961 102485 184989
rect 102513 184961 102547 184989
rect 102575 184961 102609 184989
rect 102637 184961 102671 184989
rect 102699 184961 102747 184989
rect 102437 182635 102747 184961
rect 111437 194175 111747 199205
rect 111437 194147 111485 194175
rect 111513 194147 111547 194175
rect 111575 194147 111609 194175
rect 111637 194147 111671 194175
rect 111699 194147 111747 194175
rect 111437 194113 111747 194147
rect 111437 194085 111485 194113
rect 111513 194085 111547 194113
rect 111575 194085 111609 194113
rect 111637 194085 111671 194113
rect 111699 194085 111747 194113
rect 111437 194051 111747 194085
rect 111437 194023 111485 194051
rect 111513 194023 111547 194051
rect 111575 194023 111609 194051
rect 111637 194023 111671 194051
rect 111699 194023 111747 194051
rect 111437 193989 111747 194023
rect 111437 193961 111485 193989
rect 111513 193961 111547 193989
rect 111575 193961 111609 193989
rect 111637 193961 111671 193989
rect 111699 193961 111747 193989
rect 111437 185175 111747 193961
rect 111437 185147 111485 185175
rect 111513 185147 111547 185175
rect 111575 185147 111609 185175
rect 111637 185147 111671 185175
rect 111699 185147 111747 185175
rect 111437 185113 111747 185147
rect 111437 185085 111485 185113
rect 111513 185085 111547 185113
rect 111575 185085 111609 185113
rect 111637 185085 111671 185113
rect 111699 185085 111747 185113
rect 111437 185051 111747 185085
rect 111437 185023 111485 185051
rect 111513 185023 111547 185051
rect 111575 185023 111609 185051
rect 111637 185023 111671 185051
rect 111699 185023 111747 185051
rect 111437 184989 111747 185023
rect 111437 184961 111485 184989
rect 111513 184961 111547 184989
rect 111575 184961 111609 184989
rect 111637 184961 111671 184989
rect 111699 184961 111747 184989
rect 111437 182635 111747 184961
rect 120437 194175 120747 199205
rect 120437 194147 120485 194175
rect 120513 194147 120547 194175
rect 120575 194147 120609 194175
rect 120637 194147 120671 194175
rect 120699 194147 120747 194175
rect 120437 194113 120747 194147
rect 120437 194085 120485 194113
rect 120513 194085 120547 194113
rect 120575 194085 120609 194113
rect 120637 194085 120671 194113
rect 120699 194085 120747 194113
rect 120437 194051 120747 194085
rect 120437 194023 120485 194051
rect 120513 194023 120547 194051
rect 120575 194023 120609 194051
rect 120637 194023 120671 194051
rect 120699 194023 120747 194051
rect 120437 193989 120747 194023
rect 120437 193961 120485 193989
rect 120513 193961 120547 193989
rect 120575 193961 120609 193989
rect 120637 193961 120671 193989
rect 120699 193961 120747 193989
rect 120437 185175 120747 193961
rect 120437 185147 120485 185175
rect 120513 185147 120547 185175
rect 120575 185147 120609 185175
rect 120637 185147 120671 185175
rect 120699 185147 120747 185175
rect 120437 185113 120747 185147
rect 120437 185085 120485 185113
rect 120513 185085 120547 185113
rect 120575 185085 120609 185113
rect 120637 185085 120671 185113
rect 120699 185085 120747 185113
rect 120437 185051 120747 185085
rect 120437 185023 120485 185051
rect 120513 185023 120547 185051
rect 120575 185023 120609 185051
rect 120637 185023 120671 185051
rect 120699 185023 120747 185051
rect 120437 184989 120747 185023
rect 120437 184961 120485 184989
rect 120513 184961 120547 184989
rect 120575 184961 120609 184989
rect 120637 184961 120671 184989
rect 120699 184961 120747 184989
rect 120437 182635 120747 184961
rect 129437 194175 129747 199205
rect 129437 194147 129485 194175
rect 129513 194147 129547 194175
rect 129575 194147 129609 194175
rect 129637 194147 129671 194175
rect 129699 194147 129747 194175
rect 129437 194113 129747 194147
rect 129437 194085 129485 194113
rect 129513 194085 129547 194113
rect 129575 194085 129609 194113
rect 129637 194085 129671 194113
rect 129699 194085 129747 194113
rect 129437 194051 129747 194085
rect 129437 194023 129485 194051
rect 129513 194023 129547 194051
rect 129575 194023 129609 194051
rect 129637 194023 129671 194051
rect 129699 194023 129747 194051
rect 129437 193989 129747 194023
rect 129437 193961 129485 193989
rect 129513 193961 129547 193989
rect 129575 193961 129609 193989
rect 129637 193961 129671 193989
rect 129699 193961 129747 193989
rect 129437 185175 129747 193961
rect 129437 185147 129485 185175
rect 129513 185147 129547 185175
rect 129575 185147 129609 185175
rect 129637 185147 129671 185175
rect 129699 185147 129747 185175
rect 129437 185113 129747 185147
rect 129437 185085 129485 185113
rect 129513 185085 129547 185113
rect 129575 185085 129609 185113
rect 129637 185085 129671 185113
rect 129699 185085 129747 185113
rect 129437 185051 129747 185085
rect 129437 185023 129485 185051
rect 129513 185023 129547 185051
rect 129575 185023 129609 185051
rect 129637 185023 129671 185051
rect 129699 185023 129747 185051
rect 129437 184989 129747 185023
rect 129437 184961 129485 184989
rect 129513 184961 129547 184989
rect 129575 184961 129609 184989
rect 129637 184961 129671 184989
rect 129699 184961 129747 184989
rect 129437 182635 129747 184961
rect 138437 194175 138747 199205
rect 138437 194147 138485 194175
rect 138513 194147 138547 194175
rect 138575 194147 138609 194175
rect 138637 194147 138671 194175
rect 138699 194147 138747 194175
rect 138437 194113 138747 194147
rect 138437 194085 138485 194113
rect 138513 194085 138547 194113
rect 138575 194085 138609 194113
rect 138637 194085 138671 194113
rect 138699 194085 138747 194113
rect 138437 194051 138747 194085
rect 138437 194023 138485 194051
rect 138513 194023 138547 194051
rect 138575 194023 138609 194051
rect 138637 194023 138671 194051
rect 138699 194023 138747 194051
rect 138437 193989 138747 194023
rect 138437 193961 138485 193989
rect 138513 193961 138547 193989
rect 138575 193961 138609 193989
rect 138637 193961 138671 193989
rect 138699 193961 138747 193989
rect 138437 185175 138747 193961
rect 138437 185147 138485 185175
rect 138513 185147 138547 185175
rect 138575 185147 138609 185175
rect 138637 185147 138671 185175
rect 138699 185147 138747 185175
rect 138437 185113 138747 185147
rect 138437 185085 138485 185113
rect 138513 185085 138547 185113
rect 138575 185085 138609 185113
rect 138637 185085 138671 185113
rect 138699 185085 138747 185113
rect 138437 185051 138747 185085
rect 138437 185023 138485 185051
rect 138513 185023 138547 185051
rect 138575 185023 138609 185051
rect 138637 185023 138671 185051
rect 138699 185023 138747 185051
rect 138437 184989 138747 185023
rect 138437 184961 138485 184989
rect 138513 184961 138547 184989
rect 138575 184961 138609 184989
rect 138637 184961 138671 184989
rect 138699 184961 138747 184989
rect 138437 182635 138747 184961
rect 147437 194175 147747 199205
rect 147437 194147 147485 194175
rect 147513 194147 147547 194175
rect 147575 194147 147609 194175
rect 147637 194147 147671 194175
rect 147699 194147 147747 194175
rect 147437 194113 147747 194147
rect 147437 194085 147485 194113
rect 147513 194085 147547 194113
rect 147575 194085 147609 194113
rect 147637 194085 147671 194113
rect 147699 194085 147747 194113
rect 147437 194051 147747 194085
rect 147437 194023 147485 194051
rect 147513 194023 147547 194051
rect 147575 194023 147609 194051
rect 147637 194023 147671 194051
rect 147699 194023 147747 194051
rect 147437 193989 147747 194023
rect 147437 193961 147485 193989
rect 147513 193961 147547 193989
rect 147575 193961 147609 193989
rect 147637 193961 147671 193989
rect 147699 193961 147747 193989
rect 147437 185175 147747 193961
rect 147437 185147 147485 185175
rect 147513 185147 147547 185175
rect 147575 185147 147609 185175
rect 147637 185147 147671 185175
rect 147699 185147 147747 185175
rect 147437 185113 147747 185147
rect 147437 185085 147485 185113
rect 147513 185085 147547 185113
rect 147575 185085 147609 185113
rect 147637 185085 147671 185113
rect 147699 185085 147747 185113
rect 147437 185051 147747 185085
rect 147437 185023 147485 185051
rect 147513 185023 147547 185051
rect 147575 185023 147609 185051
rect 147637 185023 147671 185051
rect 147699 185023 147747 185051
rect 147437 184989 147747 185023
rect 147437 184961 147485 184989
rect 147513 184961 147547 184989
rect 147575 184961 147609 184989
rect 147637 184961 147671 184989
rect 147699 184961 147747 184989
rect 147437 182635 147747 184961
rect 154577 191175 154887 199961
rect 154577 191147 154625 191175
rect 154653 191147 154687 191175
rect 154715 191147 154749 191175
rect 154777 191147 154811 191175
rect 154839 191147 154887 191175
rect 154577 191113 154887 191147
rect 154577 191085 154625 191113
rect 154653 191085 154687 191113
rect 154715 191085 154749 191113
rect 154777 191085 154811 191113
rect 154839 191085 154887 191113
rect 154577 191051 154887 191085
rect 154577 191023 154625 191051
rect 154653 191023 154687 191051
rect 154715 191023 154749 191051
rect 154777 191023 154811 191051
rect 154839 191023 154887 191051
rect 154577 190989 154887 191023
rect 154577 190961 154625 190989
rect 154653 190961 154687 190989
rect 154715 190961 154749 190989
rect 154777 190961 154811 190989
rect 154839 190961 154887 190989
rect 52224 182175 52384 182192
rect 52224 182147 52259 182175
rect 52287 182147 52321 182175
rect 52349 182147 52384 182175
rect 52224 182113 52384 182147
rect 52224 182085 52259 182113
rect 52287 182085 52321 182113
rect 52349 182085 52384 182113
rect 52224 182051 52384 182085
rect 52224 182023 52259 182051
rect 52287 182023 52321 182051
rect 52349 182023 52384 182051
rect 52224 181989 52384 182023
rect 52224 181961 52259 181989
rect 52287 181961 52321 181989
rect 52349 181961 52384 181989
rect 52224 181944 52384 181961
rect 67584 182175 67744 182192
rect 67584 182147 67619 182175
rect 67647 182147 67681 182175
rect 67709 182147 67744 182175
rect 67584 182113 67744 182147
rect 67584 182085 67619 182113
rect 67647 182085 67681 182113
rect 67709 182085 67744 182113
rect 67584 182051 67744 182085
rect 67584 182023 67619 182051
rect 67647 182023 67681 182051
rect 67709 182023 67744 182051
rect 67584 181989 67744 182023
rect 67584 181961 67619 181989
rect 67647 181961 67681 181989
rect 67709 181961 67744 181989
rect 67584 181944 67744 181961
rect 82944 182175 83104 182192
rect 82944 182147 82979 182175
rect 83007 182147 83041 182175
rect 83069 182147 83104 182175
rect 82944 182113 83104 182147
rect 82944 182085 82979 182113
rect 83007 182085 83041 182113
rect 83069 182085 83104 182113
rect 82944 182051 83104 182085
rect 82944 182023 82979 182051
rect 83007 182023 83041 182051
rect 83069 182023 83104 182051
rect 82944 181989 83104 182023
rect 82944 181961 82979 181989
rect 83007 181961 83041 181989
rect 83069 181961 83104 181989
rect 82944 181944 83104 181961
rect 98304 182175 98464 182192
rect 98304 182147 98339 182175
rect 98367 182147 98401 182175
rect 98429 182147 98464 182175
rect 98304 182113 98464 182147
rect 98304 182085 98339 182113
rect 98367 182085 98401 182113
rect 98429 182085 98464 182113
rect 98304 182051 98464 182085
rect 98304 182023 98339 182051
rect 98367 182023 98401 182051
rect 98429 182023 98464 182051
rect 98304 181989 98464 182023
rect 98304 181961 98339 181989
rect 98367 181961 98401 181989
rect 98429 181961 98464 181989
rect 98304 181944 98464 181961
rect 113664 182175 113824 182192
rect 113664 182147 113699 182175
rect 113727 182147 113761 182175
rect 113789 182147 113824 182175
rect 113664 182113 113824 182147
rect 113664 182085 113699 182113
rect 113727 182085 113761 182113
rect 113789 182085 113824 182113
rect 113664 182051 113824 182085
rect 113664 182023 113699 182051
rect 113727 182023 113761 182051
rect 113789 182023 113824 182051
rect 113664 181989 113824 182023
rect 113664 181961 113699 181989
rect 113727 181961 113761 181989
rect 113789 181961 113824 181989
rect 113664 181944 113824 181961
rect 129024 182175 129184 182192
rect 129024 182147 129059 182175
rect 129087 182147 129121 182175
rect 129149 182147 129184 182175
rect 129024 182113 129184 182147
rect 129024 182085 129059 182113
rect 129087 182085 129121 182113
rect 129149 182085 129184 182113
rect 129024 182051 129184 182085
rect 129024 182023 129059 182051
rect 129087 182023 129121 182051
rect 129149 182023 129184 182051
rect 129024 181989 129184 182023
rect 129024 181961 129059 181989
rect 129087 181961 129121 181989
rect 129149 181961 129184 181989
rect 129024 181944 129184 181961
rect 144384 182175 144544 182192
rect 144384 182147 144419 182175
rect 144447 182147 144481 182175
rect 144509 182147 144544 182175
rect 144384 182113 144544 182147
rect 144384 182085 144419 182113
rect 144447 182085 144481 182113
rect 144509 182085 144544 182113
rect 144384 182051 144544 182085
rect 144384 182023 144419 182051
rect 144447 182023 144481 182051
rect 144509 182023 144544 182051
rect 144384 181989 144544 182023
rect 144384 181961 144419 181989
rect 144447 181961 144481 181989
rect 144509 181961 144544 181989
rect 144384 181944 144544 181961
rect 154577 182175 154887 190961
rect 154577 182147 154625 182175
rect 154653 182147 154687 182175
rect 154715 182147 154749 182175
rect 154777 182147 154811 182175
rect 154839 182147 154887 182175
rect 154577 182113 154887 182147
rect 154577 182085 154625 182113
rect 154653 182085 154687 182113
rect 154715 182085 154749 182113
rect 154777 182085 154811 182113
rect 154839 182085 154887 182113
rect 154577 182051 154887 182085
rect 154577 182023 154625 182051
rect 154653 182023 154687 182051
rect 154715 182023 154749 182051
rect 154777 182023 154811 182051
rect 154839 182023 154887 182051
rect 154577 181989 154887 182023
rect 154577 181961 154625 181989
rect 154653 181961 154687 181989
rect 154715 181961 154749 181989
rect 154777 181961 154811 181989
rect 154839 181961 154887 181989
rect 48437 176147 48485 176175
rect 48513 176147 48547 176175
rect 48575 176147 48609 176175
rect 48637 176147 48671 176175
rect 48699 176147 48747 176175
rect 48437 176113 48747 176147
rect 48437 176085 48485 176113
rect 48513 176085 48547 176113
rect 48575 176085 48609 176113
rect 48637 176085 48671 176113
rect 48699 176085 48747 176113
rect 48437 176051 48747 176085
rect 48437 176023 48485 176051
rect 48513 176023 48547 176051
rect 48575 176023 48609 176051
rect 48637 176023 48671 176051
rect 48699 176023 48747 176051
rect 48437 175989 48747 176023
rect 48437 175961 48485 175989
rect 48513 175961 48547 175989
rect 48575 175961 48609 175989
rect 48637 175961 48671 175989
rect 48699 175961 48747 175989
rect 48437 167175 48747 175961
rect 59904 176175 60064 176192
rect 59904 176147 59939 176175
rect 59967 176147 60001 176175
rect 60029 176147 60064 176175
rect 59904 176113 60064 176147
rect 59904 176085 59939 176113
rect 59967 176085 60001 176113
rect 60029 176085 60064 176113
rect 59904 176051 60064 176085
rect 59904 176023 59939 176051
rect 59967 176023 60001 176051
rect 60029 176023 60064 176051
rect 59904 175989 60064 176023
rect 59904 175961 59939 175989
rect 59967 175961 60001 175989
rect 60029 175961 60064 175989
rect 59904 175944 60064 175961
rect 75264 176175 75424 176192
rect 75264 176147 75299 176175
rect 75327 176147 75361 176175
rect 75389 176147 75424 176175
rect 75264 176113 75424 176147
rect 75264 176085 75299 176113
rect 75327 176085 75361 176113
rect 75389 176085 75424 176113
rect 75264 176051 75424 176085
rect 75264 176023 75299 176051
rect 75327 176023 75361 176051
rect 75389 176023 75424 176051
rect 75264 175989 75424 176023
rect 75264 175961 75299 175989
rect 75327 175961 75361 175989
rect 75389 175961 75424 175989
rect 75264 175944 75424 175961
rect 90624 176175 90784 176192
rect 90624 176147 90659 176175
rect 90687 176147 90721 176175
rect 90749 176147 90784 176175
rect 90624 176113 90784 176147
rect 90624 176085 90659 176113
rect 90687 176085 90721 176113
rect 90749 176085 90784 176113
rect 90624 176051 90784 176085
rect 90624 176023 90659 176051
rect 90687 176023 90721 176051
rect 90749 176023 90784 176051
rect 90624 175989 90784 176023
rect 90624 175961 90659 175989
rect 90687 175961 90721 175989
rect 90749 175961 90784 175989
rect 90624 175944 90784 175961
rect 105984 176175 106144 176192
rect 105984 176147 106019 176175
rect 106047 176147 106081 176175
rect 106109 176147 106144 176175
rect 105984 176113 106144 176147
rect 105984 176085 106019 176113
rect 106047 176085 106081 176113
rect 106109 176085 106144 176113
rect 105984 176051 106144 176085
rect 105984 176023 106019 176051
rect 106047 176023 106081 176051
rect 106109 176023 106144 176051
rect 105984 175989 106144 176023
rect 105984 175961 106019 175989
rect 106047 175961 106081 175989
rect 106109 175961 106144 175989
rect 105984 175944 106144 175961
rect 121344 176175 121504 176192
rect 121344 176147 121379 176175
rect 121407 176147 121441 176175
rect 121469 176147 121504 176175
rect 121344 176113 121504 176147
rect 121344 176085 121379 176113
rect 121407 176085 121441 176113
rect 121469 176085 121504 176113
rect 121344 176051 121504 176085
rect 121344 176023 121379 176051
rect 121407 176023 121441 176051
rect 121469 176023 121504 176051
rect 121344 175989 121504 176023
rect 121344 175961 121379 175989
rect 121407 175961 121441 175989
rect 121469 175961 121504 175989
rect 121344 175944 121504 175961
rect 136704 176175 136864 176192
rect 136704 176147 136739 176175
rect 136767 176147 136801 176175
rect 136829 176147 136864 176175
rect 136704 176113 136864 176147
rect 136704 176085 136739 176113
rect 136767 176085 136801 176113
rect 136829 176085 136864 176113
rect 136704 176051 136864 176085
rect 136704 176023 136739 176051
rect 136767 176023 136801 176051
rect 136829 176023 136864 176051
rect 136704 175989 136864 176023
rect 136704 175961 136739 175989
rect 136767 175961 136801 175989
rect 136829 175961 136864 175989
rect 136704 175944 136864 175961
rect 52224 173175 52384 173192
rect 52224 173147 52259 173175
rect 52287 173147 52321 173175
rect 52349 173147 52384 173175
rect 52224 173113 52384 173147
rect 52224 173085 52259 173113
rect 52287 173085 52321 173113
rect 52349 173085 52384 173113
rect 52224 173051 52384 173085
rect 52224 173023 52259 173051
rect 52287 173023 52321 173051
rect 52349 173023 52384 173051
rect 52224 172989 52384 173023
rect 52224 172961 52259 172989
rect 52287 172961 52321 172989
rect 52349 172961 52384 172989
rect 52224 172944 52384 172961
rect 67584 173175 67744 173192
rect 67584 173147 67619 173175
rect 67647 173147 67681 173175
rect 67709 173147 67744 173175
rect 67584 173113 67744 173147
rect 67584 173085 67619 173113
rect 67647 173085 67681 173113
rect 67709 173085 67744 173113
rect 67584 173051 67744 173085
rect 67584 173023 67619 173051
rect 67647 173023 67681 173051
rect 67709 173023 67744 173051
rect 67584 172989 67744 173023
rect 67584 172961 67619 172989
rect 67647 172961 67681 172989
rect 67709 172961 67744 172989
rect 67584 172944 67744 172961
rect 82944 173175 83104 173192
rect 82944 173147 82979 173175
rect 83007 173147 83041 173175
rect 83069 173147 83104 173175
rect 82944 173113 83104 173147
rect 82944 173085 82979 173113
rect 83007 173085 83041 173113
rect 83069 173085 83104 173113
rect 82944 173051 83104 173085
rect 82944 173023 82979 173051
rect 83007 173023 83041 173051
rect 83069 173023 83104 173051
rect 82944 172989 83104 173023
rect 82944 172961 82979 172989
rect 83007 172961 83041 172989
rect 83069 172961 83104 172989
rect 82944 172944 83104 172961
rect 98304 173175 98464 173192
rect 98304 173147 98339 173175
rect 98367 173147 98401 173175
rect 98429 173147 98464 173175
rect 98304 173113 98464 173147
rect 98304 173085 98339 173113
rect 98367 173085 98401 173113
rect 98429 173085 98464 173113
rect 98304 173051 98464 173085
rect 98304 173023 98339 173051
rect 98367 173023 98401 173051
rect 98429 173023 98464 173051
rect 98304 172989 98464 173023
rect 98304 172961 98339 172989
rect 98367 172961 98401 172989
rect 98429 172961 98464 172989
rect 98304 172944 98464 172961
rect 113664 173175 113824 173192
rect 113664 173147 113699 173175
rect 113727 173147 113761 173175
rect 113789 173147 113824 173175
rect 113664 173113 113824 173147
rect 113664 173085 113699 173113
rect 113727 173085 113761 173113
rect 113789 173085 113824 173113
rect 113664 173051 113824 173085
rect 113664 173023 113699 173051
rect 113727 173023 113761 173051
rect 113789 173023 113824 173051
rect 113664 172989 113824 173023
rect 113664 172961 113699 172989
rect 113727 172961 113761 172989
rect 113789 172961 113824 172989
rect 113664 172944 113824 172961
rect 129024 173175 129184 173192
rect 129024 173147 129059 173175
rect 129087 173147 129121 173175
rect 129149 173147 129184 173175
rect 129024 173113 129184 173147
rect 129024 173085 129059 173113
rect 129087 173085 129121 173113
rect 129149 173085 129184 173113
rect 129024 173051 129184 173085
rect 129024 173023 129059 173051
rect 129087 173023 129121 173051
rect 129149 173023 129184 173051
rect 129024 172989 129184 173023
rect 129024 172961 129059 172989
rect 129087 172961 129121 172989
rect 129149 172961 129184 172989
rect 129024 172944 129184 172961
rect 144384 173175 144544 173192
rect 144384 173147 144419 173175
rect 144447 173147 144481 173175
rect 144509 173147 144544 173175
rect 144384 173113 144544 173147
rect 144384 173085 144419 173113
rect 144447 173085 144481 173113
rect 144509 173085 144544 173113
rect 144384 173051 144544 173085
rect 144384 173023 144419 173051
rect 144447 173023 144481 173051
rect 144509 173023 144544 173051
rect 144384 172989 144544 173023
rect 144384 172961 144419 172989
rect 144447 172961 144481 172989
rect 144509 172961 144544 172989
rect 144384 172944 144544 172961
rect 154577 173175 154887 181961
rect 154577 173147 154625 173175
rect 154653 173147 154687 173175
rect 154715 173147 154749 173175
rect 154777 173147 154811 173175
rect 154839 173147 154887 173175
rect 154577 173113 154887 173147
rect 154577 173085 154625 173113
rect 154653 173085 154687 173113
rect 154715 173085 154749 173113
rect 154777 173085 154811 173113
rect 154839 173085 154887 173113
rect 154577 173051 154887 173085
rect 154577 173023 154625 173051
rect 154653 173023 154687 173051
rect 154715 173023 154749 173051
rect 154777 173023 154811 173051
rect 154839 173023 154887 173051
rect 154577 172989 154887 173023
rect 154577 172961 154625 172989
rect 154653 172961 154687 172989
rect 154715 172961 154749 172989
rect 154777 172961 154811 172989
rect 154839 172961 154887 172989
rect 48437 167147 48485 167175
rect 48513 167147 48547 167175
rect 48575 167147 48609 167175
rect 48637 167147 48671 167175
rect 48699 167147 48747 167175
rect 48437 167113 48747 167147
rect 48437 167085 48485 167113
rect 48513 167085 48547 167113
rect 48575 167085 48609 167113
rect 48637 167085 48671 167113
rect 48699 167085 48747 167113
rect 48437 167051 48747 167085
rect 48437 167023 48485 167051
rect 48513 167023 48547 167051
rect 48575 167023 48609 167051
rect 48637 167023 48671 167051
rect 48699 167023 48747 167051
rect 48437 166989 48747 167023
rect 48437 166961 48485 166989
rect 48513 166961 48547 166989
rect 48575 166961 48609 166989
rect 48637 166961 48671 166989
rect 48699 166961 48747 166989
rect 48437 158175 48747 166961
rect 59904 167175 60064 167192
rect 59904 167147 59939 167175
rect 59967 167147 60001 167175
rect 60029 167147 60064 167175
rect 59904 167113 60064 167147
rect 59904 167085 59939 167113
rect 59967 167085 60001 167113
rect 60029 167085 60064 167113
rect 59904 167051 60064 167085
rect 59904 167023 59939 167051
rect 59967 167023 60001 167051
rect 60029 167023 60064 167051
rect 59904 166989 60064 167023
rect 59904 166961 59939 166989
rect 59967 166961 60001 166989
rect 60029 166961 60064 166989
rect 59904 166944 60064 166961
rect 75264 167175 75424 167192
rect 75264 167147 75299 167175
rect 75327 167147 75361 167175
rect 75389 167147 75424 167175
rect 75264 167113 75424 167147
rect 75264 167085 75299 167113
rect 75327 167085 75361 167113
rect 75389 167085 75424 167113
rect 75264 167051 75424 167085
rect 75264 167023 75299 167051
rect 75327 167023 75361 167051
rect 75389 167023 75424 167051
rect 75264 166989 75424 167023
rect 75264 166961 75299 166989
rect 75327 166961 75361 166989
rect 75389 166961 75424 166989
rect 75264 166944 75424 166961
rect 90624 167175 90784 167192
rect 90624 167147 90659 167175
rect 90687 167147 90721 167175
rect 90749 167147 90784 167175
rect 90624 167113 90784 167147
rect 90624 167085 90659 167113
rect 90687 167085 90721 167113
rect 90749 167085 90784 167113
rect 90624 167051 90784 167085
rect 90624 167023 90659 167051
rect 90687 167023 90721 167051
rect 90749 167023 90784 167051
rect 90624 166989 90784 167023
rect 90624 166961 90659 166989
rect 90687 166961 90721 166989
rect 90749 166961 90784 166989
rect 90624 166944 90784 166961
rect 105984 167175 106144 167192
rect 105984 167147 106019 167175
rect 106047 167147 106081 167175
rect 106109 167147 106144 167175
rect 105984 167113 106144 167147
rect 105984 167085 106019 167113
rect 106047 167085 106081 167113
rect 106109 167085 106144 167113
rect 105984 167051 106144 167085
rect 105984 167023 106019 167051
rect 106047 167023 106081 167051
rect 106109 167023 106144 167051
rect 105984 166989 106144 167023
rect 105984 166961 106019 166989
rect 106047 166961 106081 166989
rect 106109 166961 106144 166989
rect 105984 166944 106144 166961
rect 121344 167175 121504 167192
rect 121344 167147 121379 167175
rect 121407 167147 121441 167175
rect 121469 167147 121504 167175
rect 121344 167113 121504 167147
rect 121344 167085 121379 167113
rect 121407 167085 121441 167113
rect 121469 167085 121504 167113
rect 121344 167051 121504 167085
rect 121344 167023 121379 167051
rect 121407 167023 121441 167051
rect 121469 167023 121504 167051
rect 121344 166989 121504 167023
rect 121344 166961 121379 166989
rect 121407 166961 121441 166989
rect 121469 166961 121504 166989
rect 121344 166944 121504 166961
rect 136704 167175 136864 167192
rect 136704 167147 136739 167175
rect 136767 167147 136801 167175
rect 136829 167147 136864 167175
rect 136704 167113 136864 167147
rect 136704 167085 136739 167113
rect 136767 167085 136801 167113
rect 136829 167085 136864 167113
rect 136704 167051 136864 167085
rect 136704 167023 136739 167051
rect 136767 167023 136801 167051
rect 136829 167023 136864 167051
rect 136704 166989 136864 167023
rect 136704 166961 136739 166989
rect 136767 166961 136801 166989
rect 136829 166961 136864 166989
rect 136704 166944 136864 166961
rect 52224 164175 52384 164192
rect 52224 164147 52259 164175
rect 52287 164147 52321 164175
rect 52349 164147 52384 164175
rect 52224 164113 52384 164147
rect 52224 164085 52259 164113
rect 52287 164085 52321 164113
rect 52349 164085 52384 164113
rect 52224 164051 52384 164085
rect 52224 164023 52259 164051
rect 52287 164023 52321 164051
rect 52349 164023 52384 164051
rect 52224 163989 52384 164023
rect 52224 163961 52259 163989
rect 52287 163961 52321 163989
rect 52349 163961 52384 163989
rect 52224 163944 52384 163961
rect 67584 164175 67744 164192
rect 67584 164147 67619 164175
rect 67647 164147 67681 164175
rect 67709 164147 67744 164175
rect 67584 164113 67744 164147
rect 67584 164085 67619 164113
rect 67647 164085 67681 164113
rect 67709 164085 67744 164113
rect 67584 164051 67744 164085
rect 67584 164023 67619 164051
rect 67647 164023 67681 164051
rect 67709 164023 67744 164051
rect 67584 163989 67744 164023
rect 67584 163961 67619 163989
rect 67647 163961 67681 163989
rect 67709 163961 67744 163989
rect 67584 163944 67744 163961
rect 82944 164175 83104 164192
rect 82944 164147 82979 164175
rect 83007 164147 83041 164175
rect 83069 164147 83104 164175
rect 82944 164113 83104 164147
rect 82944 164085 82979 164113
rect 83007 164085 83041 164113
rect 83069 164085 83104 164113
rect 82944 164051 83104 164085
rect 82944 164023 82979 164051
rect 83007 164023 83041 164051
rect 83069 164023 83104 164051
rect 82944 163989 83104 164023
rect 82944 163961 82979 163989
rect 83007 163961 83041 163989
rect 83069 163961 83104 163989
rect 82944 163944 83104 163961
rect 98304 164175 98464 164192
rect 98304 164147 98339 164175
rect 98367 164147 98401 164175
rect 98429 164147 98464 164175
rect 98304 164113 98464 164147
rect 98304 164085 98339 164113
rect 98367 164085 98401 164113
rect 98429 164085 98464 164113
rect 98304 164051 98464 164085
rect 98304 164023 98339 164051
rect 98367 164023 98401 164051
rect 98429 164023 98464 164051
rect 98304 163989 98464 164023
rect 98304 163961 98339 163989
rect 98367 163961 98401 163989
rect 98429 163961 98464 163989
rect 98304 163944 98464 163961
rect 113664 164175 113824 164192
rect 113664 164147 113699 164175
rect 113727 164147 113761 164175
rect 113789 164147 113824 164175
rect 113664 164113 113824 164147
rect 113664 164085 113699 164113
rect 113727 164085 113761 164113
rect 113789 164085 113824 164113
rect 113664 164051 113824 164085
rect 113664 164023 113699 164051
rect 113727 164023 113761 164051
rect 113789 164023 113824 164051
rect 113664 163989 113824 164023
rect 113664 163961 113699 163989
rect 113727 163961 113761 163989
rect 113789 163961 113824 163989
rect 113664 163944 113824 163961
rect 129024 164175 129184 164192
rect 129024 164147 129059 164175
rect 129087 164147 129121 164175
rect 129149 164147 129184 164175
rect 129024 164113 129184 164147
rect 129024 164085 129059 164113
rect 129087 164085 129121 164113
rect 129149 164085 129184 164113
rect 129024 164051 129184 164085
rect 129024 164023 129059 164051
rect 129087 164023 129121 164051
rect 129149 164023 129184 164051
rect 129024 163989 129184 164023
rect 129024 163961 129059 163989
rect 129087 163961 129121 163989
rect 129149 163961 129184 163989
rect 129024 163944 129184 163961
rect 144384 164175 144544 164192
rect 144384 164147 144419 164175
rect 144447 164147 144481 164175
rect 144509 164147 144544 164175
rect 144384 164113 144544 164147
rect 144384 164085 144419 164113
rect 144447 164085 144481 164113
rect 144509 164085 144544 164113
rect 144384 164051 144544 164085
rect 144384 164023 144419 164051
rect 144447 164023 144481 164051
rect 144509 164023 144544 164051
rect 144384 163989 144544 164023
rect 144384 163961 144419 163989
rect 144447 163961 144481 163989
rect 144509 163961 144544 163989
rect 144384 163944 144544 163961
rect 154577 164175 154887 172961
rect 154577 164147 154625 164175
rect 154653 164147 154687 164175
rect 154715 164147 154749 164175
rect 154777 164147 154811 164175
rect 154839 164147 154887 164175
rect 154577 164113 154887 164147
rect 154577 164085 154625 164113
rect 154653 164085 154687 164113
rect 154715 164085 154749 164113
rect 154777 164085 154811 164113
rect 154839 164085 154887 164113
rect 154577 164051 154887 164085
rect 154577 164023 154625 164051
rect 154653 164023 154687 164051
rect 154715 164023 154749 164051
rect 154777 164023 154811 164051
rect 154839 164023 154887 164051
rect 154577 163989 154887 164023
rect 154577 163961 154625 163989
rect 154653 163961 154687 163989
rect 154715 163961 154749 163989
rect 154777 163961 154811 163989
rect 154839 163961 154887 163989
rect 48437 158147 48485 158175
rect 48513 158147 48547 158175
rect 48575 158147 48609 158175
rect 48637 158147 48671 158175
rect 48699 158147 48747 158175
rect 48437 158113 48747 158147
rect 48437 158085 48485 158113
rect 48513 158085 48547 158113
rect 48575 158085 48609 158113
rect 48637 158085 48671 158113
rect 48699 158085 48747 158113
rect 48437 158051 48747 158085
rect 48437 158023 48485 158051
rect 48513 158023 48547 158051
rect 48575 158023 48609 158051
rect 48637 158023 48671 158051
rect 48699 158023 48747 158051
rect 48437 157989 48747 158023
rect 48437 157961 48485 157989
rect 48513 157961 48547 157989
rect 48575 157961 48609 157989
rect 48637 157961 48671 157989
rect 48699 157961 48747 157989
rect 48437 149175 48747 157961
rect 59904 158175 60064 158192
rect 59904 158147 59939 158175
rect 59967 158147 60001 158175
rect 60029 158147 60064 158175
rect 59904 158113 60064 158147
rect 59904 158085 59939 158113
rect 59967 158085 60001 158113
rect 60029 158085 60064 158113
rect 59904 158051 60064 158085
rect 59904 158023 59939 158051
rect 59967 158023 60001 158051
rect 60029 158023 60064 158051
rect 59904 157989 60064 158023
rect 59904 157961 59939 157989
rect 59967 157961 60001 157989
rect 60029 157961 60064 157989
rect 59904 157944 60064 157961
rect 75264 158175 75424 158192
rect 75264 158147 75299 158175
rect 75327 158147 75361 158175
rect 75389 158147 75424 158175
rect 75264 158113 75424 158147
rect 75264 158085 75299 158113
rect 75327 158085 75361 158113
rect 75389 158085 75424 158113
rect 75264 158051 75424 158085
rect 75264 158023 75299 158051
rect 75327 158023 75361 158051
rect 75389 158023 75424 158051
rect 75264 157989 75424 158023
rect 75264 157961 75299 157989
rect 75327 157961 75361 157989
rect 75389 157961 75424 157989
rect 75264 157944 75424 157961
rect 90624 158175 90784 158192
rect 90624 158147 90659 158175
rect 90687 158147 90721 158175
rect 90749 158147 90784 158175
rect 90624 158113 90784 158147
rect 90624 158085 90659 158113
rect 90687 158085 90721 158113
rect 90749 158085 90784 158113
rect 90624 158051 90784 158085
rect 90624 158023 90659 158051
rect 90687 158023 90721 158051
rect 90749 158023 90784 158051
rect 90624 157989 90784 158023
rect 90624 157961 90659 157989
rect 90687 157961 90721 157989
rect 90749 157961 90784 157989
rect 90624 157944 90784 157961
rect 105984 158175 106144 158192
rect 105984 158147 106019 158175
rect 106047 158147 106081 158175
rect 106109 158147 106144 158175
rect 105984 158113 106144 158147
rect 105984 158085 106019 158113
rect 106047 158085 106081 158113
rect 106109 158085 106144 158113
rect 105984 158051 106144 158085
rect 105984 158023 106019 158051
rect 106047 158023 106081 158051
rect 106109 158023 106144 158051
rect 105984 157989 106144 158023
rect 105984 157961 106019 157989
rect 106047 157961 106081 157989
rect 106109 157961 106144 157989
rect 105984 157944 106144 157961
rect 121344 158175 121504 158192
rect 121344 158147 121379 158175
rect 121407 158147 121441 158175
rect 121469 158147 121504 158175
rect 121344 158113 121504 158147
rect 121344 158085 121379 158113
rect 121407 158085 121441 158113
rect 121469 158085 121504 158113
rect 121344 158051 121504 158085
rect 121344 158023 121379 158051
rect 121407 158023 121441 158051
rect 121469 158023 121504 158051
rect 121344 157989 121504 158023
rect 121344 157961 121379 157989
rect 121407 157961 121441 157989
rect 121469 157961 121504 157989
rect 121344 157944 121504 157961
rect 136704 158175 136864 158192
rect 136704 158147 136739 158175
rect 136767 158147 136801 158175
rect 136829 158147 136864 158175
rect 136704 158113 136864 158147
rect 136704 158085 136739 158113
rect 136767 158085 136801 158113
rect 136829 158085 136864 158113
rect 136704 158051 136864 158085
rect 136704 158023 136739 158051
rect 136767 158023 136801 158051
rect 136829 158023 136864 158051
rect 136704 157989 136864 158023
rect 136704 157961 136739 157989
rect 136767 157961 136801 157989
rect 136829 157961 136864 157989
rect 136704 157944 136864 157961
rect 52224 155175 52384 155192
rect 52224 155147 52259 155175
rect 52287 155147 52321 155175
rect 52349 155147 52384 155175
rect 52224 155113 52384 155147
rect 52224 155085 52259 155113
rect 52287 155085 52321 155113
rect 52349 155085 52384 155113
rect 52224 155051 52384 155085
rect 52224 155023 52259 155051
rect 52287 155023 52321 155051
rect 52349 155023 52384 155051
rect 52224 154989 52384 155023
rect 52224 154961 52259 154989
rect 52287 154961 52321 154989
rect 52349 154961 52384 154989
rect 52224 154944 52384 154961
rect 67584 155175 67744 155192
rect 67584 155147 67619 155175
rect 67647 155147 67681 155175
rect 67709 155147 67744 155175
rect 67584 155113 67744 155147
rect 67584 155085 67619 155113
rect 67647 155085 67681 155113
rect 67709 155085 67744 155113
rect 67584 155051 67744 155085
rect 67584 155023 67619 155051
rect 67647 155023 67681 155051
rect 67709 155023 67744 155051
rect 67584 154989 67744 155023
rect 67584 154961 67619 154989
rect 67647 154961 67681 154989
rect 67709 154961 67744 154989
rect 67584 154944 67744 154961
rect 82944 155175 83104 155192
rect 82944 155147 82979 155175
rect 83007 155147 83041 155175
rect 83069 155147 83104 155175
rect 82944 155113 83104 155147
rect 82944 155085 82979 155113
rect 83007 155085 83041 155113
rect 83069 155085 83104 155113
rect 82944 155051 83104 155085
rect 82944 155023 82979 155051
rect 83007 155023 83041 155051
rect 83069 155023 83104 155051
rect 82944 154989 83104 155023
rect 82944 154961 82979 154989
rect 83007 154961 83041 154989
rect 83069 154961 83104 154989
rect 82944 154944 83104 154961
rect 98304 155175 98464 155192
rect 98304 155147 98339 155175
rect 98367 155147 98401 155175
rect 98429 155147 98464 155175
rect 98304 155113 98464 155147
rect 98304 155085 98339 155113
rect 98367 155085 98401 155113
rect 98429 155085 98464 155113
rect 98304 155051 98464 155085
rect 98304 155023 98339 155051
rect 98367 155023 98401 155051
rect 98429 155023 98464 155051
rect 98304 154989 98464 155023
rect 98304 154961 98339 154989
rect 98367 154961 98401 154989
rect 98429 154961 98464 154989
rect 98304 154944 98464 154961
rect 113664 155175 113824 155192
rect 113664 155147 113699 155175
rect 113727 155147 113761 155175
rect 113789 155147 113824 155175
rect 113664 155113 113824 155147
rect 113664 155085 113699 155113
rect 113727 155085 113761 155113
rect 113789 155085 113824 155113
rect 113664 155051 113824 155085
rect 113664 155023 113699 155051
rect 113727 155023 113761 155051
rect 113789 155023 113824 155051
rect 113664 154989 113824 155023
rect 113664 154961 113699 154989
rect 113727 154961 113761 154989
rect 113789 154961 113824 154989
rect 113664 154944 113824 154961
rect 129024 155175 129184 155192
rect 129024 155147 129059 155175
rect 129087 155147 129121 155175
rect 129149 155147 129184 155175
rect 129024 155113 129184 155147
rect 129024 155085 129059 155113
rect 129087 155085 129121 155113
rect 129149 155085 129184 155113
rect 129024 155051 129184 155085
rect 129024 155023 129059 155051
rect 129087 155023 129121 155051
rect 129149 155023 129184 155051
rect 129024 154989 129184 155023
rect 129024 154961 129059 154989
rect 129087 154961 129121 154989
rect 129149 154961 129184 154989
rect 129024 154944 129184 154961
rect 144384 155175 144544 155192
rect 144384 155147 144419 155175
rect 144447 155147 144481 155175
rect 144509 155147 144544 155175
rect 144384 155113 144544 155147
rect 144384 155085 144419 155113
rect 144447 155085 144481 155113
rect 144509 155085 144544 155113
rect 144384 155051 144544 155085
rect 144384 155023 144419 155051
rect 144447 155023 144481 155051
rect 144509 155023 144544 155051
rect 144384 154989 144544 155023
rect 144384 154961 144419 154989
rect 144447 154961 144481 154989
rect 144509 154961 144544 154989
rect 144384 154944 144544 154961
rect 154577 155175 154887 163961
rect 154577 155147 154625 155175
rect 154653 155147 154687 155175
rect 154715 155147 154749 155175
rect 154777 155147 154811 155175
rect 154839 155147 154887 155175
rect 154577 155113 154887 155147
rect 154577 155085 154625 155113
rect 154653 155085 154687 155113
rect 154715 155085 154749 155113
rect 154777 155085 154811 155113
rect 154839 155085 154887 155113
rect 154577 155051 154887 155085
rect 154577 155023 154625 155051
rect 154653 155023 154687 155051
rect 154715 155023 154749 155051
rect 154777 155023 154811 155051
rect 154839 155023 154887 155051
rect 154577 154989 154887 155023
rect 154577 154961 154625 154989
rect 154653 154961 154687 154989
rect 154715 154961 154749 154989
rect 154777 154961 154811 154989
rect 154839 154961 154887 154989
rect 48437 149147 48485 149175
rect 48513 149147 48547 149175
rect 48575 149147 48609 149175
rect 48637 149147 48671 149175
rect 48699 149147 48747 149175
rect 48437 149113 48747 149147
rect 48437 149085 48485 149113
rect 48513 149085 48547 149113
rect 48575 149085 48609 149113
rect 48637 149085 48671 149113
rect 48699 149085 48747 149113
rect 48437 149051 48747 149085
rect 48437 149023 48485 149051
rect 48513 149023 48547 149051
rect 48575 149023 48609 149051
rect 48637 149023 48671 149051
rect 48699 149023 48747 149051
rect 48437 148989 48747 149023
rect 48437 148961 48485 148989
rect 48513 148961 48547 148989
rect 48575 148961 48609 148989
rect 48637 148961 48671 148989
rect 48699 148961 48747 148989
rect 48437 140175 48747 148961
rect 59904 149175 60064 149192
rect 59904 149147 59939 149175
rect 59967 149147 60001 149175
rect 60029 149147 60064 149175
rect 59904 149113 60064 149147
rect 59904 149085 59939 149113
rect 59967 149085 60001 149113
rect 60029 149085 60064 149113
rect 59904 149051 60064 149085
rect 59904 149023 59939 149051
rect 59967 149023 60001 149051
rect 60029 149023 60064 149051
rect 59904 148989 60064 149023
rect 59904 148961 59939 148989
rect 59967 148961 60001 148989
rect 60029 148961 60064 148989
rect 59904 148944 60064 148961
rect 75264 149175 75424 149192
rect 75264 149147 75299 149175
rect 75327 149147 75361 149175
rect 75389 149147 75424 149175
rect 75264 149113 75424 149147
rect 75264 149085 75299 149113
rect 75327 149085 75361 149113
rect 75389 149085 75424 149113
rect 75264 149051 75424 149085
rect 75264 149023 75299 149051
rect 75327 149023 75361 149051
rect 75389 149023 75424 149051
rect 75264 148989 75424 149023
rect 75264 148961 75299 148989
rect 75327 148961 75361 148989
rect 75389 148961 75424 148989
rect 75264 148944 75424 148961
rect 90624 149175 90784 149192
rect 90624 149147 90659 149175
rect 90687 149147 90721 149175
rect 90749 149147 90784 149175
rect 90624 149113 90784 149147
rect 90624 149085 90659 149113
rect 90687 149085 90721 149113
rect 90749 149085 90784 149113
rect 90624 149051 90784 149085
rect 90624 149023 90659 149051
rect 90687 149023 90721 149051
rect 90749 149023 90784 149051
rect 90624 148989 90784 149023
rect 90624 148961 90659 148989
rect 90687 148961 90721 148989
rect 90749 148961 90784 148989
rect 90624 148944 90784 148961
rect 105984 149175 106144 149192
rect 105984 149147 106019 149175
rect 106047 149147 106081 149175
rect 106109 149147 106144 149175
rect 105984 149113 106144 149147
rect 105984 149085 106019 149113
rect 106047 149085 106081 149113
rect 106109 149085 106144 149113
rect 105984 149051 106144 149085
rect 105984 149023 106019 149051
rect 106047 149023 106081 149051
rect 106109 149023 106144 149051
rect 105984 148989 106144 149023
rect 105984 148961 106019 148989
rect 106047 148961 106081 148989
rect 106109 148961 106144 148989
rect 105984 148944 106144 148961
rect 121344 149175 121504 149192
rect 121344 149147 121379 149175
rect 121407 149147 121441 149175
rect 121469 149147 121504 149175
rect 121344 149113 121504 149147
rect 121344 149085 121379 149113
rect 121407 149085 121441 149113
rect 121469 149085 121504 149113
rect 121344 149051 121504 149085
rect 121344 149023 121379 149051
rect 121407 149023 121441 149051
rect 121469 149023 121504 149051
rect 121344 148989 121504 149023
rect 121344 148961 121379 148989
rect 121407 148961 121441 148989
rect 121469 148961 121504 148989
rect 121344 148944 121504 148961
rect 136704 149175 136864 149192
rect 136704 149147 136739 149175
rect 136767 149147 136801 149175
rect 136829 149147 136864 149175
rect 136704 149113 136864 149147
rect 136704 149085 136739 149113
rect 136767 149085 136801 149113
rect 136829 149085 136864 149113
rect 136704 149051 136864 149085
rect 136704 149023 136739 149051
rect 136767 149023 136801 149051
rect 136829 149023 136864 149051
rect 136704 148989 136864 149023
rect 136704 148961 136739 148989
rect 136767 148961 136801 148989
rect 136829 148961 136864 148989
rect 136704 148944 136864 148961
rect 52224 146175 52384 146192
rect 52224 146147 52259 146175
rect 52287 146147 52321 146175
rect 52349 146147 52384 146175
rect 52224 146113 52384 146147
rect 52224 146085 52259 146113
rect 52287 146085 52321 146113
rect 52349 146085 52384 146113
rect 52224 146051 52384 146085
rect 52224 146023 52259 146051
rect 52287 146023 52321 146051
rect 52349 146023 52384 146051
rect 52224 145989 52384 146023
rect 52224 145961 52259 145989
rect 52287 145961 52321 145989
rect 52349 145961 52384 145989
rect 52224 145944 52384 145961
rect 67584 146175 67744 146192
rect 67584 146147 67619 146175
rect 67647 146147 67681 146175
rect 67709 146147 67744 146175
rect 67584 146113 67744 146147
rect 67584 146085 67619 146113
rect 67647 146085 67681 146113
rect 67709 146085 67744 146113
rect 67584 146051 67744 146085
rect 67584 146023 67619 146051
rect 67647 146023 67681 146051
rect 67709 146023 67744 146051
rect 67584 145989 67744 146023
rect 67584 145961 67619 145989
rect 67647 145961 67681 145989
rect 67709 145961 67744 145989
rect 67584 145944 67744 145961
rect 82944 146175 83104 146192
rect 82944 146147 82979 146175
rect 83007 146147 83041 146175
rect 83069 146147 83104 146175
rect 82944 146113 83104 146147
rect 82944 146085 82979 146113
rect 83007 146085 83041 146113
rect 83069 146085 83104 146113
rect 82944 146051 83104 146085
rect 82944 146023 82979 146051
rect 83007 146023 83041 146051
rect 83069 146023 83104 146051
rect 82944 145989 83104 146023
rect 82944 145961 82979 145989
rect 83007 145961 83041 145989
rect 83069 145961 83104 145989
rect 82944 145944 83104 145961
rect 98304 146175 98464 146192
rect 98304 146147 98339 146175
rect 98367 146147 98401 146175
rect 98429 146147 98464 146175
rect 98304 146113 98464 146147
rect 98304 146085 98339 146113
rect 98367 146085 98401 146113
rect 98429 146085 98464 146113
rect 98304 146051 98464 146085
rect 98304 146023 98339 146051
rect 98367 146023 98401 146051
rect 98429 146023 98464 146051
rect 98304 145989 98464 146023
rect 98304 145961 98339 145989
rect 98367 145961 98401 145989
rect 98429 145961 98464 145989
rect 98304 145944 98464 145961
rect 113664 146175 113824 146192
rect 113664 146147 113699 146175
rect 113727 146147 113761 146175
rect 113789 146147 113824 146175
rect 113664 146113 113824 146147
rect 113664 146085 113699 146113
rect 113727 146085 113761 146113
rect 113789 146085 113824 146113
rect 113664 146051 113824 146085
rect 113664 146023 113699 146051
rect 113727 146023 113761 146051
rect 113789 146023 113824 146051
rect 113664 145989 113824 146023
rect 113664 145961 113699 145989
rect 113727 145961 113761 145989
rect 113789 145961 113824 145989
rect 113664 145944 113824 145961
rect 129024 146175 129184 146192
rect 129024 146147 129059 146175
rect 129087 146147 129121 146175
rect 129149 146147 129184 146175
rect 129024 146113 129184 146147
rect 129024 146085 129059 146113
rect 129087 146085 129121 146113
rect 129149 146085 129184 146113
rect 129024 146051 129184 146085
rect 129024 146023 129059 146051
rect 129087 146023 129121 146051
rect 129149 146023 129184 146051
rect 129024 145989 129184 146023
rect 129024 145961 129059 145989
rect 129087 145961 129121 145989
rect 129149 145961 129184 145989
rect 129024 145944 129184 145961
rect 144384 146175 144544 146192
rect 144384 146147 144419 146175
rect 144447 146147 144481 146175
rect 144509 146147 144544 146175
rect 144384 146113 144544 146147
rect 144384 146085 144419 146113
rect 144447 146085 144481 146113
rect 144509 146085 144544 146113
rect 144384 146051 144544 146085
rect 144384 146023 144419 146051
rect 144447 146023 144481 146051
rect 144509 146023 144544 146051
rect 144384 145989 144544 146023
rect 144384 145961 144419 145989
rect 144447 145961 144481 145989
rect 144509 145961 144544 145989
rect 144384 145944 144544 145961
rect 154577 146175 154887 154961
rect 154577 146147 154625 146175
rect 154653 146147 154687 146175
rect 154715 146147 154749 146175
rect 154777 146147 154811 146175
rect 154839 146147 154887 146175
rect 154577 146113 154887 146147
rect 154577 146085 154625 146113
rect 154653 146085 154687 146113
rect 154715 146085 154749 146113
rect 154777 146085 154811 146113
rect 154839 146085 154887 146113
rect 154577 146051 154887 146085
rect 154577 146023 154625 146051
rect 154653 146023 154687 146051
rect 154715 146023 154749 146051
rect 154777 146023 154811 146051
rect 154839 146023 154887 146051
rect 154577 145989 154887 146023
rect 154577 145961 154625 145989
rect 154653 145961 154687 145989
rect 154715 145961 154749 145989
rect 154777 145961 154811 145989
rect 154839 145961 154887 145989
rect 48437 140147 48485 140175
rect 48513 140147 48547 140175
rect 48575 140147 48609 140175
rect 48637 140147 48671 140175
rect 48699 140147 48747 140175
rect 48437 140113 48747 140147
rect 48437 140085 48485 140113
rect 48513 140085 48547 140113
rect 48575 140085 48609 140113
rect 48637 140085 48671 140113
rect 48699 140085 48747 140113
rect 48437 140051 48747 140085
rect 48437 140023 48485 140051
rect 48513 140023 48547 140051
rect 48575 140023 48609 140051
rect 48637 140023 48671 140051
rect 48699 140023 48747 140051
rect 48437 139989 48747 140023
rect 48437 139961 48485 139989
rect 48513 139961 48547 139989
rect 48575 139961 48609 139989
rect 48637 139961 48671 139989
rect 48699 139961 48747 139989
rect 48437 131175 48747 139961
rect 59904 140175 60064 140192
rect 59904 140147 59939 140175
rect 59967 140147 60001 140175
rect 60029 140147 60064 140175
rect 59904 140113 60064 140147
rect 59904 140085 59939 140113
rect 59967 140085 60001 140113
rect 60029 140085 60064 140113
rect 59904 140051 60064 140085
rect 59904 140023 59939 140051
rect 59967 140023 60001 140051
rect 60029 140023 60064 140051
rect 59904 139989 60064 140023
rect 59904 139961 59939 139989
rect 59967 139961 60001 139989
rect 60029 139961 60064 139989
rect 59904 139944 60064 139961
rect 75264 140175 75424 140192
rect 75264 140147 75299 140175
rect 75327 140147 75361 140175
rect 75389 140147 75424 140175
rect 75264 140113 75424 140147
rect 75264 140085 75299 140113
rect 75327 140085 75361 140113
rect 75389 140085 75424 140113
rect 75264 140051 75424 140085
rect 75264 140023 75299 140051
rect 75327 140023 75361 140051
rect 75389 140023 75424 140051
rect 75264 139989 75424 140023
rect 75264 139961 75299 139989
rect 75327 139961 75361 139989
rect 75389 139961 75424 139989
rect 75264 139944 75424 139961
rect 90624 140175 90784 140192
rect 90624 140147 90659 140175
rect 90687 140147 90721 140175
rect 90749 140147 90784 140175
rect 90624 140113 90784 140147
rect 90624 140085 90659 140113
rect 90687 140085 90721 140113
rect 90749 140085 90784 140113
rect 90624 140051 90784 140085
rect 90624 140023 90659 140051
rect 90687 140023 90721 140051
rect 90749 140023 90784 140051
rect 90624 139989 90784 140023
rect 90624 139961 90659 139989
rect 90687 139961 90721 139989
rect 90749 139961 90784 139989
rect 90624 139944 90784 139961
rect 105984 140175 106144 140192
rect 105984 140147 106019 140175
rect 106047 140147 106081 140175
rect 106109 140147 106144 140175
rect 105984 140113 106144 140147
rect 105984 140085 106019 140113
rect 106047 140085 106081 140113
rect 106109 140085 106144 140113
rect 105984 140051 106144 140085
rect 105984 140023 106019 140051
rect 106047 140023 106081 140051
rect 106109 140023 106144 140051
rect 105984 139989 106144 140023
rect 105984 139961 106019 139989
rect 106047 139961 106081 139989
rect 106109 139961 106144 139989
rect 105984 139944 106144 139961
rect 121344 140175 121504 140192
rect 121344 140147 121379 140175
rect 121407 140147 121441 140175
rect 121469 140147 121504 140175
rect 121344 140113 121504 140147
rect 121344 140085 121379 140113
rect 121407 140085 121441 140113
rect 121469 140085 121504 140113
rect 121344 140051 121504 140085
rect 121344 140023 121379 140051
rect 121407 140023 121441 140051
rect 121469 140023 121504 140051
rect 121344 139989 121504 140023
rect 121344 139961 121379 139989
rect 121407 139961 121441 139989
rect 121469 139961 121504 139989
rect 121344 139944 121504 139961
rect 136704 140175 136864 140192
rect 136704 140147 136739 140175
rect 136767 140147 136801 140175
rect 136829 140147 136864 140175
rect 136704 140113 136864 140147
rect 136704 140085 136739 140113
rect 136767 140085 136801 140113
rect 136829 140085 136864 140113
rect 136704 140051 136864 140085
rect 136704 140023 136739 140051
rect 136767 140023 136801 140051
rect 136829 140023 136864 140051
rect 136704 139989 136864 140023
rect 136704 139961 136739 139989
rect 136767 139961 136801 139989
rect 136829 139961 136864 139989
rect 136704 139944 136864 139961
rect 52224 137175 52384 137192
rect 52224 137147 52259 137175
rect 52287 137147 52321 137175
rect 52349 137147 52384 137175
rect 52224 137113 52384 137147
rect 52224 137085 52259 137113
rect 52287 137085 52321 137113
rect 52349 137085 52384 137113
rect 52224 137051 52384 137085
rect 52224 137023 52259 137051
rect 52287 137023 52321 137051
rect 52349 137023 52384 137051
rect 52224 136989 52384 137023
rect 52224 136961 52259 136989
rect 52287 136961 52321 136989
rect 52349 136961 52384 136989
rect 52224 136944 52384 136961
rect 67584 137175 67744 137192
rect 67584 137147 67619 137175
rect 67647 137147 67681 137175
rect 67709 137147 67744 137175
rect 67584 137113 67744 137147
rect 67584 137085 67619 137113
rect 67647 137085 67681 137113
rect 67709 137085 67744 137113
rect 67584 137051 67744 137085
rect 67584 137023 67619 137051
rect 67647 137023 67681 137051
rect 67709 137023 67744 137051
rect 67584 136989 67744 137023
rect 67584 136961 67619 136989
rect 67647 136961 67681 136989
rect 67709 136961 67744 136989
rect 67584 136944 67744 136961
rect 82944 137175 83104 137192
rect 82944 137147 82979 137175
rect 83007 137147 83041 137175
rect 83069 137147 83104 137175
rect 82944 137113 83104 137147
rect 82944 137085 82979 137113
rect 83007 137085 83041 137113
rect 83069 137085 83104 137113
rect 82944 137051 83104 137085
rect 82944 137023 82979 137051
rect 83007 137023 83041 137051
rect 83069 137023 83104 137051
rect 82944 136989 83104 137023
rect 82944 136961 82979 136989
rect 83007 136961 83041 136989
rect 83069 136961 83104 136989
rect 82944 136944 83104 136961
rect 98304 137175 98464 137192
rect 98304 137147 98339 137175
rect 98367 137147 98401 137175
rect 98429 137147 98464 137175
rect 98304 137113 98464 137147
rect 98304 137085 98339 137113
rect 98367 137085 98401 137113
rect 98429 137085 98464 137113
rect 98304 137051 98464 137085
rect 98304 137023 98339 137051
rect 98367 137023 98401 137051
rect 98429 137023 98464 137051
rect 98304 136989 98464 137023
rect 98304 136961 98339 136989
rect 98367 136961 98401 136989
rect 98429 136961 98464 136989
rect 98304 136944 98464 136961
rect 113664 137175 113824 137192
rect 113664 137147 113699 137175
rect 113727 137147 113761 137175
rect 113789 137147 113824 137175
rect 113664 137113 113824 137147
rect 113664 137085 113699 137113
rect 113727 137085 113761 137113
rect 113789 137085 113824 137113
rect 113664 137051 113824 137085
rect 113664 137023 113699 137051
rect 113727 137023 113761 137051
rect 113789 137023 113824 137051
rect 113664 136989 113824 137023
rect 113664 136961 113699 136989
rect 113727 136961 113761 136989
rect 113789 136961 113824 136989
rect 113664 136944 113824 136961
rect 129024 137175 129184 137192
rect 129024 137147 129059 137175
rect 129087 137147 129121 137175
rect 129149 137147 129184 137175
rect 129024 137113 129184 137147
rect 129024 137085 129059 137113
rect 129087 137085 129121 137113
rect 129149 137085 129184 137113
rect 129024 137051 129184 137085
rect 129024 137023 129059 137051
rect 129087 137023 129121 137051
rect 129149 137023 129184 137051
rect 129024 136989 129184 137023
rect 129024 136961 129059 136989
rect 129087 136961 129121 136989
rect 129149 136961 129184 136989
rect 129024 136944 129184 136961
rect 144384 137175 144544 137192
rect 144384 137147 144419 137175
rect 144447 137147 144481 137175
rect 144509 137147 144544 137175
rect 144384 137113 144544 137147
rect 144384 137085 144419 137113
rect 144447 137085 144481 137113
rect 144509 137085 144544 137113
rect 144384 137051 144544 137085
rect 144384 137023 144419 137051
rect 144447 137023 144481 137051
rect 144509 137023 144544 137051
rect 144384 136989 144544 137023
rect 144384 136961 144419 136989
rect 144447 136961 144481 136989
rect 144509 136961 144544 136989
rect 144384 136944 144544 136961
rect 154577 137175 154887 145961
rect 154577 137147 154625 137175
rect 154653 137147 154687 137175
rect 154715 137147 154749 137175
rect 154777 137147 154811 137175
rect 154839 137147 154887 137175
rect 154577 137113 154887 137147
rect 154577 137085 154625 137113
rect 154653 137085 154687 137113
rect 154715 137085 154749 137113
rect 154777 137085 154811 137113
rect 154839 137085 154887 137113
rect 154577 137051 154887 137085
rect 154577 137023 154625 137051
rect 154653 137023 154687 137051
rect 154715 137023 154749 137051
rect 154777 137023 154811 137051
rect 154839 137023 154887 137051
rect 154577 136989 154887 137023
rect 154577 136961 154625 136989
rect 154653 136961 154687 136989
rect 154715 136961 154749 136989
rect 154777 136961 154811 136989
rect 154839 136961 154887 136989
rect 48437 131147 48485 131175
rect 48513 131147 48547 131175
rect 48575 131147 48609 131175
rect 48637 131147 48671 131175
rect 48699 131147 48747 131175
rect 48437 131113 48747 131147
rect 48437 131085 48485 131113
rect 48513 131085 48547 131113
rect 48575 131085 48609 131113
rect 48637 131085 48671 131113
rect 48699 131085 48747 131113
rect 48437 131051 48747 131085
rect 48437 131023 48485 131051
rect 48513 131023 48547 131051
rect 48575 131023 48609 131051
rect 48637 131023 48671 131051
rect 48699 131023 48747 131051
rect 48437 130989 48747 131023
rect 48437 130961 48485 130989
rect 48513 130961 48547 130989
rect 48575 130961 48609 130989
rect 48637 130961 48671 130989
rect 48699 130961 48747 130989
rect 48437 122175 48747 130961
rect 59904 131175 60064 131192
rect 59904 131147 59939 131175
rect 59967 131147 60001 131175
rect 60029 131147 60064 131175
rect 59904 131113 60064 131147
rect 59904 131085 59939 131113
rect 59967 131085 60001 131113
rect 60029 131085 60064 131113
rect 59904 131051 60064 131085
rect 59904 131023 59939 131051
rect 59967 131023 60001 131051
rect 60029 131023 60064 131051
rect 59904 130989 60064 131023
rect 59904 130961 59939 130989
rect 59967 130961 60001 130989
rect 60029 130961 60064 130989
rect 59904 130944 60064 130961
rect 75264 131175 75424 131192
rect 75264 131147 75299 131175
rect 75327 131147 75361 131175
rect 75389 131147 75424 131175
rect 75264 131113 75424 131147
rect 75264 131085 75299 131113
rect 75327 131085 75361 131113
rect 75389 131085 75424 131113
rect 75264 131051 75424 131085
rect 75264 131023 75299 131051
rect 75327 131023 75361 131051
rect 75389 131023 75424 131051
rect 75264 130989 75424 131023
rect 75264 130961 75299 130989
rect 75327 130961 75361 130989
rect 75389 130961 75424 130989
rect 75264 130944 75424 130961
rect 90624 131175 90784 131192
rect 90624 131147 90659 131175
rect 90687 131147 90721 131175
rect 90749 131147 90784 131175
rect 90624 131113 90784 131147
rect 90624 131085 90659 131113
rect 90687 131085 90721 131113
rect 90749 131085 90784 131113
rect 90624 131051 90784 131085
rect 90624 131023 90659 131051
rect 90687 131023 90721 131051
rect 90749 131023 90784 131051
rect 90624 130989 90784 131023
rect 90624 130961 90659 130989
rect 90687 130961 90721 130989
rect 90749 130961 90784 130989
rect 90624 130944 90784 130961
rect 105984 131175 106144 131192
rect 105984 131147 106019 131175
rect 106047 131147 106081 131175
rect 106109 131147 106144 131175
rect 105984 131113 106144 131147
rect 105984 131085 106019 131113
rect 106047 131085 106081 131113
rect 106109 131085 106144 131113
rect 105984 131051 106144 131085
rect 105984 131023 106019 131051
rect 106047 131023 106081 131051
rect 106109 131023 106144 131051
rect 105984 130989 106144 131023
rect 105984 130961 106019 130989
rect 106047 130961 106081 130989
rect 106109 130961 106144 130989
rect 105984 130944 106144 130961
rect 121344 131175 121504 131192
rect 121344 131147 121379 131175
rect 121407 131147 121441 131175
rect 121469 131147 121504 131175
rect 121344 131113 121504 131147
rect 121344 131085 121379 131113
rect 121407 131085 121441 131113
rect 121469 131085 121504 131113
rect 121344 131051 121504 131085
rect 121344 131023 121379 131051
rect 121407 131023 121441 131051
rect 121469 131023 121504 131051
rect 121344 130989 121504 131023
rect 121344 130961 121379 130989
rect 121407 130961 121441 130989
rect 121469 130961 121504 130989
rect 121344 130944 121504 130961
rect 136704 131175 136864 131192
rect 136704 131147 136739 131175
rect 136767 131147 136801 131175
rect 136829 131147 136864 131175
rect 136704 131113 136864 131147
rect 136704 131085 136739 131113
rect 136767 131085 136801 131113
rect 136829 131085 136864 131113
rect 136704 131051 136864 131085
rect 136704 131023 136739 131051
rect 136767 131023 136801 131051
rect 136829 131023 136864 131051
rect 136704 130989 136864 131023
rect 136704 130961 136739 130989
rect 136767 130961 136801 130989
rect 136829 130961 136864 130989
rect 136704 130944 136864 130961
rect 52224 128175 52384 128192
rect 52224 128147 52259 128175
rect 52287 128147 52321 128175
rect 52349 128147 52384 128175
rect 52224 128113 52384 128147
rect 52224 128085 52259 128113
rect 52287 128085 52321 128113
rect 52349 128085 52384 128113
rect 52224 128051 52384 128085
rect 52224 128023 52259 128051
rect 52287 128023 52321 128051
rect 52349 128023 52384 128051
rect 52224 127989 52384 128023
rect 52224 127961 52259 127989
rect 52287 127961 52321 127989
rect 52349 127961 52384 127989
rect 52224 127944 52384 127961
rect 67584 128175 67744 128192
rect 67584 128147 67619 128175
rect 67647 128147 67681 128175
rect 67709 128147 67744 128175
rect 67584 128113 67744 128147
rect 67584 128085 67619 128113
rect 67647 128085 67681 128113
rect 67709 128085 67744 128113
rect 67584 128051 67744 128085
rect 67584 128023 67619 128051
rect 67647 128023 67681 128051
rect 67709 128023 67744 128051
rect 67584 127989 67744 128023
rect 67584 127961 67619 127989
rect 67647 127961 67681 127989
rect 67709 127961 67744 127989
rect 67584 127944 67744 127961
rect 82944 128175 83104 128192
rect 82944 128147 82979 128175
rect 83007 128147 83041 128175
rect 83069 128147 83104 128175
rect 82944 128113 83104 128147
rect 82944 128085 82979 128113
rect 83007 128085 83041 128113
rect 83069 128085 83104 128113
rect 82944 128051 83104 128085
rect 82944 128023 82979 128051
rect 83007 128023 83041 128051
rect 83069 128023 83104 128051
rect 82944 127989 83104 128023
rect 82944 127961 82979 127989
rect 83007 127961 83041 127989
rect 83069 127961 83104 127989
rect 82944 127944 83104 127961
rect 98304 128175 98464 128192
rect 98304 128147 98339 128175
rect 98367 128147 98401 128175
rect 98429 128147 98464 128175
rect 98304 128113 98464 128147
rect 98304 128085 98339 128113
rect 98367 128085 98401 128113
rect 98429 128085 98464 128113
rect 98304 128051 98464 128085
rect 98304 128023 98339 128051
rect 98367 128023 98401 128051
rect 98429 128023 98464 128051
rect 98304 127989 98464 128023
rect 98304 127961 98339 127989
rect 98367 127961 98401 127989
rect 98429 127961 98464 127989
rect 98304 127944 98464 127961
rect 113664 128175 113824 128192
rect 113664 128147 113699 128175
rect 113727 128147 113761 128175
rect 113789 128147 113824 128175
rect 113664 128113 113824 128147
rect 113664 128085 113699 128113
rect 113727 128085 113761 128113
rect 113789 128085 113824 128113
rect 113664 128051 113824 128085
rect 113664 128023 113699 128051
rect 113727 128023 113761 128051
rect 113789 128023 113824 128051
rect 113664 127989 113824 128023
rect 113664 127961 113699 127989
rect 113727 127961 113761 127989
rect 113789 127961 113824 127989
rect 113664 127944 113824 127961
rect 129024 128175 129184 128192
rect 129024 128147 129059 128175
rect 129087 128147 129121 128175
rect 129149 128147 129184 128175
rect 129024 128113 129184 128147
rect 129024 128085 129059 128113
rect 129087 128085 129121 128113
rect 129149 128085 129184 128113
rect 129024 128051 129184 128085
rect 129024 128023 129059 128051
rect 129087 128023 129121 128051
rect 129149 128023 129184 128051
rect 129024 127989 129184 128023
rect 129024 127961 129059 127989
rect 129087 127961 129121 127989
rect 129149 127961 129184 127989
rect 129024 127944 129184 127961
rect 144384 128175 144544 128192
rect 144384 128147 144419 128175
rect 144447 128147 144481 128175
rect 144509 128147 144544 128175
rect 144384 128113 144544 128147
rect 144384 128085 144419 128113
rect 144447 128085 144481 128113
rect 144509 128085 144544 128113
rect 144384 128051 144544 128085
rect 144384 128023 144419 128051
rect 144447 128023 144481 128051
rect 144509 128023 144544 128051
rect 144384 127989 144544 128023
rect 144384 127961 144419 127989
rect 144447 127961 144481 127989
rect 144509 127961 144544 127989
rect 144384 127944 144544 127961
rect 154577 128175 154887 136961
rect 154577 128147 154625 128175
rect 154653 128147 154687 128175
rect 154715 128147 154749 128175
rect 154777 128147 154811 128175
rect 154839 128147 154887 128175
rect 154577 128113 154887 128147
rect 154577 128085 154625 128113
rect 154653 128085 154687 128113
rect 154715 128085 154749 128113
rect 154777 128085 154811 128113
rect 154839 128085 154887 128113
rect 154577 128051 154887 128085
rect 154577 128023 154625 128051
rect 154653 128023 154687 128051
rect 154715 128023 154749 128051
rect 154777 128023 154811 128051
rect 154839 128023 154887 128051
rect 154577 127989 154887 128023
rect 154577 127961 154625 127989
rect 154653 127961 154687 127989
rect 154715 127961 154749 127989
rect 154777 127961 154811 127989
rect 154839 127961 154887 127989
rect 48437 122147 48485 122175
rect 48513 122147 48547 122175
rect 48575 122147 48609 122175
rect 48637 122147 48671 122175
rect 48699 122147 48747 122175
rect 48437 122113 48747 122147
rect 48437 122085 48485 122113
rect 48513 122085 48547 122113
rect 48575 122085 48609 122113
rect 48637 122085 48671 122113
rect 48699 122085 48747 122113
rect 48437 122051 48747 122085
rect 48437 122023 48485 122051
rect 48513 122023 48547 122051
rect 48575 122023 48609 122051
rect 48637 122023 48671 122051
rect 48699 122023 48747 122051
rect 48437 121989 48747 122023
rect 48437 121961 48485 121989
rect 48513 121961 48547 121989
rect 48575 121961 48609 121989
rect 48637 121961 48671 121989
rect 48699 121961 48747 121989
rect 48437 113175 48747 121961
rect 48437 113147 48485 113175
rect 48513 113147 48547 113175
rect 48575 113147 48609 113175
rect 48637 113147 48671 113175
rect 48699 113147 48747 113175
rect 48437 113113 48747 113147
rect 48437 113085 48485 113113
rect 48513 113085 48547 113113
rect 48575 113085 48609 113113
rect 48637 113085 48671 113113
rect 48699 113085 48747 113113
rect 48437 113051 48747 113085
rect 48437 113023 48485 113051
rect 48513 113023 48547 113051
rect 48575 113023 48609 113051
rect 48637 113023 48671 113051
rect 48699 113023 48747 113051
rect 48437 112989 48747 113023
rect 48437 112961 48485 112989
rect 48513 112961 48547 112989
rect 48575 112961 48609 112989
rect 48637 112961 48671 112989
rect 48699 112961 48747 112989
rect 48437 104175 48747 112961
rect 55577 119175 55887 124261
rect 55577 119147 55625 119175
rect 55653 119147 55687 119175
rect 55715 119147 55749 119175
rect 55777 119147 55811 119175
rect 55839 119147 55887 119175
rect 55577 119113 55887 119147
rect 55577 119085 55625 119113
rect 55653 119085 55687 119113
rect 55715 119085 55749 119113
rect 55777 119085 55811 119113
rect 55839 119085 55887 119113
rect 55577 119051 55887 119085
rect 55577 119023 55625 119051
rect 55653 119023 55687 119051
rect 55715 119023 55749 119051
rect 55777 119023 55811 119051
rect 55839 119023 55887 119051
rect 55577 118989 55887 119023
rect 55577 118961 55625 118989
rect 55653 118961 55687 118989
rect 55715 118961 55749 118989
rect 55777 118961 55811 118989
rect 55839 118961 55887 118989
rect 55577 110175 55887 118961
rect 55577 110147 55625 110175
rect 55653 110147 55687 110175
rect 55715 110147 55749 110175
rect 55777 110147 55811 110175
rect 55839 110147 55887 110175
rect 55577 110113 55887 110147
rect 55577 110085 55625 110113
rect 55653 110085 55687 110113
rect 55715 110085 55749 110113
rect 55777 110085 55811 110113
rect 55839 110085 55887 110113
rect 55577 110051 55887 110085
rect 55577 110023 55625 110051
rect 55653 110023 55687 110051
rect 55715 110023 55749 110051
rect 55777 110023 55811 110051
rect 55839 110023 55887 110051
rect 55577 109989 55887 110023
rect 55577 109961 55625 109989
rect 55653 109961 55687 109989
rect 55715 109961 55749 109989
rect 55777 109961 55811 109989
rect 55839 109961 55887 109989
rect 48437 104147 48485 104175
rect 48513 104147 48547 104175
rect 48575 104147 48609 104175
rect 48637 104147 48671 104175
rect 48699 104147 48747 104175
rect 48437 104113 48747 104147
rect 48437 104085 48485 104113
rect 48513 104085 48547 104113
rect 48575 104085 48609 104113
rect 48637 104085 48671 104113
rect 48699 104085 48747 104113
rect 48437 104051 48747 104085
rect 48437 104023 48485 104051
rect 48513 104023 48547 104051
rect 48575 104023 48609 104051
rect 48637 104023 48671 104051
rect 48699 104023 48747 104051
rect 48437 103989 48747 104023
rect 48437 103961 48485 103989
rect 48513 103961 48547 103989
rect 48575 103961 48609 103989
rect 48637 103961 48671 103989
rect 48699 103961 48747 103989
rect 48437 95175 48747 103961
rect 54474 104175 54634 104192
rect 54474 104147 54509 104175
rect 54537 104147 54571 104175
rect 54599 104147 54634 104175
rect 54474 104113 54634 104147
rect 54474 104085 54509 104113
rect 54537 104085 54571 104113
rect 54599 104085 54634 104113
rect 54474 104051 54634 104085
rect 54474 104023 54509 104051
rect 54537 104023 54571 104051
rect 54599 104023 54634 104051
rect 54474 103989 54634 104023
rect 54474 103961 54509 103989
rect 54537 103961 54571 103989
rect 54599 103961 54634 103989
rect 54474 103944 54634 103961
rect 52224 101175 52384 101192
rect 52224 101147 52259 101175
rect 52287 101147 52321 101175
rect 52349 101147 52384 101175
rect 52224 101113 52384 101147
rect 52224 101085 52259 101113
rect 52287 101085 52321 101113
rect 52349 101085 52384 101113
rect 52224 101051 52384 101085
rect 52224 101023 52259 101051
rect 52287 101023 52321 101051
rect 52349 101023 52384 101051
rect 52224 100989 52384 101023
rect 52224 100961 52259 100989
rect 52287 100961 52321 100989
rect 52349 100961 52384 100989
rect 52224 100944 52384 100961
rect 55577 101175 55887 109961
rect 57437 122175 57747 124261
rect 57437 122147 57485 122175
rect 57513 122147 57547 122175
rect 57575 122147 57609 122175
rect 57637 122147 57671 122175
rect 57699 122147 57747 122175
rect 57437 122113 57747 122147
rect 57437 122085 57485 122113
rect 57513 122085 57547 122113
rect 57575 122085 57609 122113
rect 57637 122085 57671 122113
rect 57699 122085 57747 122113
rect 57437 122051 57747 122085
rect 57437 122023 57485 122051
rect 57513 122023 57547 122051
rect 57575 122023 57609 122051
rect 57637 122023 57671 122051
rect 57699 122023 57747 122051
rect 57437 121989 57747 122023
rect 57437 121961 57485 121989
rect 57513 121961 57547 121989
rect 57575 121961 57609 121989
rect 57637 121961 57671 121989
rect 57699 121961 57747 121989
rect 57437 113175 57747 121961
rect 57437 113147 57485 113175
rect 57513 113147 57547 113175
rect 57575 113147 57609 113175
rect 57637 113147 57671 113175
rect 57699 113147 57747 113175
rect 57437 113113 57747 113147
rect 57437 113085 57485 113113
rect 57513 113085 57547 113113
rect 57575 113085 57609 113113
rect 57637 113085 57671 113113
rect 57699 113085 57747 113113
rect 57437 113051 57747 113085
rect 57437 113023 57485 113051
rect 57513 113023 57547 113051
rect 57575 113023 57609 113051
rect 57637 113023 57671 113051
rect 57699 113023 57747 113051
rect 57437 112989 57747 113023
rect 57437 112961 57485 112989
rect 57513 112961 57547 112989
rect 57575 112961 57609 112989
rect 57637 112961 57671 112989
rect 57699 112961 57747 112989
rect 57437 104175 57747 112961
rect 64577 119175 64887 124261
rect 64577 119147 64625 119175
rect 64653 119147 64687 119175
rect 64715 119147 64749 119175
rect 64777 119147 64811 119175
rect 64839 119147 64887 119175
rect 64577 119113 64887 119147
rect 64577 119085 64625 119113
rect 64653 119085 64687 119113
rect 64715 119085 64749 119113
rect 64777 119085 64811 119113
rect 64839 119085 64887 119113
rect 64577 119051 64887 119085
rect 64577 119023 64625 119051
rect 64653 119023 64687 119051
rect 64715 119023 64749 119051
rect 64777 119023 64811 119051
rect 64839 119023 64887 119051
rect 64577 118989 64887 119023
rect 64577 118961 64625 118989
rect 64653 118961 64687 118989
rect 64715 118961 64749 118989
rect 64777 118961 64811 118989
rect 64839 118961 64887 118989
rect 64577 110175 64887 118961
rect 64577 110147 64625 110175
rect 64653 110147 64687 110175
rect 64715 110147 64749 110175
rect 64777 110147 64811 110175
rect 64839 110147 64887 110175
rect 64577 110113 64887 110147
rect 64577 110085 64625 110113
rect 64653 110085 64687 110113
rect 64715 110085 64749 110113
rect 64777 110085 64811 110113
rect 64839 110085 64887 110113
rect 64577 110051 64887 110085
rect 64577 110023 64625 110051
rect 64653 110023 64687 110051
rect 64715 110023 64749 110051
rect 64777 110023 64811 110051
rect 64839 110023 64887 110051
rect 64577 109989 64887 110023
rect 64577 109961 64625 109989
rect 64653 109961 64687 109989
rect 64715 109961 64749 109989
rect 64777 109961 64811 109989
rect 64839 109961 64887 109989
rect 57437 104147 57485 104175
rect 57513 104147 57547 104175
rect 57575 104147 57609 104175
rect 57637 104147 57671 104175
rect 57699 104147 57747 104175
rect 57437 104113 57747 104147
rect 57437 104085 57485 104113
rect 57513 104085 57547 104113
rect 57575 104085 57609 104113
rect 57637 104085 57671 104113
rect 57699 104085 57747 104113
rect 57437 104051 57747 104085
rect 57437 104023 57485 104051
rect 57513 104023 57547 104051
rect 57575 104023 57609 104051
rect 57637 104023 57671 104051
rect 57699 104023 57747 104051
rect 57437 103989 57747 104023
rect 57437 103961 57485 103989
rect 57513 103961 57547 103989
rect 57575 103961 57609 103989
rect 57637 103961 57671 103989
rect 57699 103961 57747 103989
rect 55577 101147 55625 101175
rect 55653 101147 55687 101175
rect 55715 101147 55749 101175
rect 55777 101147 55811 101175
rect 55839 101147 55887 101175
rect 55577 101113 55887 101147
rect 55577 101085 55625 101113
rect 55653 101085 55687 101113
rect 55715 101085 55749 101113
rect 55777 101085 55811 101113
rect 55839 101085 55887 101113
rect 55577 101051 55887 101085
rect 55577 101023 55625 101051
rect 55653 101023 55687 101051
rect 55715 101023 55749 101051
rect 55777 101023 55811 101051
rect 55839 101023 55887 101051
rect 55577 100989 55887 101023
rect 55577 100961 55625 100989
rect 55653 100961 55687 100989
rect 55715 100961 55749 100989
rect 55777 100961 55811 100989
rect 55839 100961 55887 100989
rect 48437 95147 48485 95175
rect 48513 95147 48547 95175
rect 48575 95147 48609 95175
rect 48637 95147 48671 95175
rect 48699 95147 48747 95175
rect 48437 95113 48747 95147
rect 48437 95085 48485 95113
rect 48513 95085 48547 95113
rect 48575 95085 48609 95113
rect 48637 95085 48671 95113
rect 48699 95085 48747 95113
rect 48437 95051 48747 95085
rect 48437 95023 48485 95051
rect 48513 95023 48547 95051
rect 48575 95023 48609 95051
rect 48637 95023 48671 95051
rect 48699 95023 48747 95051
rect 48437 94989 48747 95023
rect 48437 94961 48485 94989
rect 48513 94961 48547 94989
rect 48575 94961 48609 94989
rect 48637 94961 48671 94989
rect 48699 94961 48747 94989
rect 48437 86175 48747 94961
rect 54474 95175 54634 95192
rect 54474 95147 54509 95175
rect 54537 95147 54571 95175
rect 54599 95147 54634 95175
rect 54474 95113 54634 95147
rect 54474 95085 54509 95113
rect 54537 95085 54571 95113
rect 54599 95085 54634 95113
rect 54474 95051 54634 95085
rect 54474 95023 54509 95051
rect 54537 95023 54571 95051
rect 54599 95023 54634 95051
rect 54474 94989 54634 95023
rect 54474 94961 54509 94989
rect 54537 94961 54571 94989
rect 54599 94961 54634 94989
rect 54474 94944 54634 94961
rect 52224 92175 52384 92192
rect 52224 92147 52259 92175
rect 52287 92147 52321 92175
rect 52349 92147 52384 92175
rect 52224 92113 52384 92147
rect 52224 92085 52259 92113
rect 52287 92085 52321 92113
rect 52349 92085 52384 92113
rect 52224 92051 52384 92085
rect 52224 92023 52259 92051
rect 52287 92023 52321 92051
rect 52349 92023 52384 92051
rect 52224 91989 52384 92023
rect 52224 91961 52259 91989
rect 52287 91961 52321 91989
rect 52349 91961 52384 91989
rect 52224 91944 52384 91961
rect 55577 92175 55887 100961
rect 56724 101175 56884 101192
rect 56724 101147 56759 101175
rect 56787 101147 56821 101175
rect 56849 101147 56884 101175
rect 56724 101113 56884 101147
rect 56724 101085 56759 101113
rect 56787 101085 56821 101113
rect 56849 101085 56884 101113
rect 56724 101051 56884 101085
rect 56724 101023 56759 101051
rect 56787 101023 56821 101051
rect 56849 101023 56884 101051
rect 56724 100989 56884 101023
rect 56724 100961 56759 100989
rect 56787 100961 56821 100989
rect 56849 100961 56884 100989
rect 56724 100944 56884 100961
rect 57437 95175 57747 103961
rect 58974 104175 59134 104192
rect 58974 104147 59009 104175
rect 59037 104147 59071 104175
rect 59099 104147 59134 104175
rect 58974 104113 59134 104147
rect 58974 104085 59009 104113
rect 59037 104085 59071 104113
rect 59099 104085 59134 104113
rect 58974 104051 59134 104085
rect 58974 104023 59009 104051
rect 59037 104023 59071 104051
rect 59099 104023 59134 104051
rect 58974 103989 59134 104023
rect 58974 103961 59009 103989
rect 59037 103961 59071 103989
rect 59099 103961 59134 103989
rect 58974 103944 59134 103961
rect 63474 104175 63634 104192
rect 63474 104147 63509 104175
rect 63537 104147 63571 104175
rect 63599 104147 63634 104175
rect 63474 104113 63634 104147
rect 63474 104085 63509 104113
rect 63537 104085 63571 104113
rect 63599 104085 63634 104113
rect 63474 104051 63634 104085
rect 63474 104023 63509 104051
rect 63537 104023 63571 104051
rect 63599 104023 63634 104051
rect 63474 103989 63634 104023
rect 63474 103961 63509 103989
rect 63537 103961 63571 103989
rect 63599 103961 63634 103989
rect 63474 103944 63634 103961
rect 61224 101175 61384 101192
rect 61224 101147 61259 101175
rect 61287 101147 61321 101175
rect 61349 101147 61384 101175
rect 61224 101113 61384 101147
rect 61224 101085 61259 101113
rect 61287 101085 61321 101113
rect 61349 101085 61384 101113
rect 61224 101051 61384 101085
rect 61224 101023 61259 101051
rect 61287 101023 61321 101051
rect 61349 101023 61384 101051
rect 61224 100989 61384 101023
rect 61224 100961 61259 100989
rect 61287 100961 61321 100989
rect 61349 100961 61384 100989
rect 61224 100944 61384 100961
rect 64577 101175 64887 109961
rect 66437 122175 66747 124261
rect 66437 122147 66485 122175
rect 66513 122147 66547 122175
rect 66575 122147 66609 122175
rect 66637 122147 66671 122175
rect 66699 122147 66747 122175
rect 66437 122113 66747 122147
rect 66437 122085 66485 122113
rect 66513 122085 66547 122113
rect 66575 122085 66609 122113
rect 66637 122085 66671 122113
rect 66699 122085 66747 122113
rect 66437 122051 66747 122085
rect 66437 122023 66485 122051
rect 66513 122023 66547 122051
rect 66575 122023 66609 122051
rect 66637 122023 66671 122051
rect 66699 122023 66747 122051
rect 66437 121989 66747 122023
rect 66437 121961 66485 121989
rect 66513 121961 66547 121989
rect 66575 121961 66609 121989
rect 66637 121961 66671 121989
rect 66699 121961 66747 121989
rect 66437 113175 66747 121961
rect 66437 113147 66485 113175
rect 66513 113147 66547 113175
rect 66575 113147 66609 113175
rect 66637 113147 66671 113175
rect 66699 113147 66747 113175
rect 66437 113113 66747 113147
rect 66437 113085 66485 113113
rect 66513 113085 66547 113113
rect 66575 113085 66609 113113
rect 66637 113085 66671 113113
rect 66699 113085 66747 113113
rect 66437 113051 66747 113085
rect 66437 113023 66485 113051
rect 66513 113023 66547 113051
rect 66575 113023 66609 113051
rect 66637 113023 66671 113051
rect 66699 113023 66747 113051
rect 66437 112989 66747 113023
rect 66437 112961 66485 112989
rect 66513 112961 66547 112989
rect 66575 112961 66609 112989
rect 66637 112961 66671 112989
rect 66699 112961 66747 112989
rect 66437 104175 66747 112961
rect 73577 119175 73887 124261
rect 73577 119147 73625 119175
rect 73653 119147 73687 119175
rect 73715 119147 73749 119175
rect 73777 119147 73811 119175
rect 73839 119147 73887 119175
rect 73577 119113 73887 119147
rect 73577 119085 73625 119113
rect 73653 119085 73687 119113
rect 73715 119085 73749 119113
rect 73777 119085 73811 119113
rect 73839 119085 73887 119113
rect 73577 119051 73887 119085
rect 73577 119023 73625 119051
rect 73653 119023 73687 119051
rect 73715 119023 73749 119051
rect 73777 119023 73811 119051
rect 73839 119023 73887 119051
rect 73577 118989 73887 119023
rect 73577 118961 73625 118989
rect 73653 118961 73687 118989
rect 73715 118961 73749 118989
rect 73777 118961 73811 118989
rect 73839 118961 73887 118989
rect 73577 110175 73887 118961
rect 73577 110147 73625 110175
rect 73653 110147 73687 110175
rect 73715 110147 73749 110175
rect 73777 110147 73811 110175
rect 73839 110147 73887 110175
rect 73577 110113 73887 110147
rect 73577 110085 73625 110113
rect 73653 110085 73687 110113
rect 73715 110085 73749 110113
rect 73777 110085 73811 110113
rect 73839 110085 73887 110113
rect 73577 110051 73887 110085
rect 73577 110023 73625 110051
rect 73653 110023 73687 110051
rect 73715 110023 73749 110051
rect 73777 110023 73811 110051
rect 73839 110023 73887 110051
rect 73577 109989 73887 110023
rect 73577 109961 73625 109989
rect 73653 109961 73687 109989
rect 73715 109961 73749 109989
rect 73777 109961 73811 109989
rect 73839 109961 73887 109989
rect 66437 104147 66485 104175
rect 66513 104147 66547 104175
rect 66575 104147 66609 104175
rect 66637 104147 66671 104175
rect 66699 104147 66747 104175
rect 66437 104113 66747 104147
rect 66437 104085 66485 104113
rect 66513 104085 66547 104113
rect 66575 104085 66609 104113
rect 66637 104085 66671 104113
rect 66699 104085 66747 104113
rect 66437 104051 66747 104085
rect 66437 104023 66485 104051
rect 66513 104023 66547 104051
rect 66575 104023 66609 104051
rect 66637 104023 66671 104051
rect 66699 104023 66747 104051
rect 66437 103989 66747 104023
rect 66437 103961 66485 103989
rect 66513 103961 66547 103989
rect 66575 103961 66609 103989
rect 66637 103961 66671 103989
rect 66699 103961 66747 103989
rect 64577 101147 64625 101175
rect 64653 101147 64687 101175
rect 64715 101147 64749 101175
rect 64777 101147 64811 101175
rect 64839 101147 64887 101175
rect 64577 101113 64887 101147
rect 64577 101085 64625 101113
rect 64653 101085 64687 101113
rect 64715 101085 64749 101113
rect 64777 101085 64811 101113
rect 64839 101085 64887 101113
rect 64577 101051 64887 101085
rect 64577 101023 64625 101051
rect 64653 101023 64687 101051
rect 64715 101023 64749 101051
rect 64777 101023 64811 101051
rect 64839 101023 64887 101051
rect 64577 100989 64887 101023
rect 64577 100961 64625 100989
rect 64653 100961 64687 100989
rect 64715 100961 64749 100989
rect 64777 100961 64811 100989
rect 64839 100961 64887 100989
rect 57437 95147 57485 95175
rect 57513 95147 57547 95175
rect 57575 95147 57609 95175
rect 57637 95147 57671 95175
rect 57699 95147 57747 95175
rect 57437 95113 57747 95147
rect 57437 95085 57485 95113
rect 57513 95085 57547 95113
rect 57575 95085 57609 95113
rect 57637 95085 57671 95113
rect 57699 95085 57747 95113
rect 57437 95051 57747 95085
rect 57437 95023 57485 95051
rect 57513 95023 57547 95051
rect 57575 95023 57609 95051
rect 57637 95023 57671 95051
rect 57699 95023 57747 95051
rect 57437 94989 57747 95023
rect 57437 94961 57485 94989
rect 57513 94961 57547 94989
rect 57575 94961 57609 94989
rect 57637 94961 57671 94989
rect 57699 94961 57747 94989
rect 55577 92147 55625 92175
rect 55653 92147 55687 92175
rect 55715 92147 55749 92175
rect 55777 92147 55811 92175
rect 55839 92147 55887 92175
rect 55577 92113 55887 92147
rect 55577 92085 55625 92113
rect 55653 92085 55687 92113
rect 55715 92085 55749 92113
rect 55777 92085 55811 92113
rect 55839 92085 55887 92113
rect 55577 92051 55887 92085
rect 55577 92023 55625 92051
rect 55653 92023 55687 92051
rect 55715 92023 55749 92051
rect 55777 92023 55811 92051
rect 55839 92023 55887 92051
rect 55577 91989 55887 92023
rect 55577 91961 55625 91989
rect 55653 91961 55687 91989
rect 55715 91961 55749 91989
rect 55777 91961 55811 91989
rect 55839 91961 55887 91989
rect 48437 86147 48485 86175
rect 48513 86147 48547 86175
rect 48575 86147 48609 86175
rect 48637 86147 48671 86175
rect 48699 86147 48747 86175
rect 48437 86113 48747 86147
rect 48437 86085 48485 86113
rect 48513 86085 48547 86113
rect 48575 86085 48609 86113
rect 48637 86085 48671 86113
rect 48699 86085 48747 86113
rect 48437 86051 48747 86085
rect 48437 86023 48485 86051
rect 48513 86023 48547 86051
rect 48575 86023 48609 86051
rect 48637 86023 48671 86051
rect 48699 86023 48747 86051
rect 48437 85989 48747 86023
rect 48437 85961 48485 85989
rect 48513 85961 48547 85989
rect 48575 85961 48609 85989
rect 48637 85961 48671 85989
rect 48699 85961 48747 85989
rect 48437 77175 48747 85961
rect 54474 86175 54634 86192
rect 54474 86147 54509 86175
rect 54537 86147 54571 86175
rect 54599 86147 54634 86175
rect 54474 86113 54634 86147
rect 54474 86085 54509 86113
rect 54537 86085 54571 86113
rect 54599 86085 54634 86113
rect 54474 86051 54634 86085
rect 54474 86023 54509 86051
rect 54537 86023 54571 86051
rect 54599 86023 54634 86051
rect 54474 85989 54634 86023
rect 54474 85961 54509 85989
rect 54537 85961 54571 85989
rect 54599 85961 54634 85989
rect 54474 85944 54634 85961
rect 52224 83175 52384 83192
rect 52224 83147 52259 83175
rect 52287 83147 52321 83175
rect 52349 83147 52384 83175
rect 52224 83113 52384 83147
rect 52224 83085 52259 83113
rect 52287 83085 52321 83113
rect 52349 83085 52384 83113
rect 52224 83051 52384 83085
rect 52224 83023 52259 83051
rect 52287 83023 52321 83051
rect 52349 83023 52384 83051
rect 52224 82989 52384 83023
rect 52224 82961 52259 82989
rect 52287 82961 52321 82989
rect 52349 82961 52384 82989
rect 52224 82944 52384 82961
rect 55577 83175 55887 91961
rect 56724 92175 56884 92192
rect 56724 92147 56759 92175
rect 56787 92147 56821 92175
rect 56849 92147 56884 92175
rect 56724 92113 56884 92147
rect 56724 92085 56759 92113
rect 56787 92085 56821 92113
rect 56849 92085 56884 92113
rect 56724 92051 56884 92085
rect 56724 92023 56759 92051
rect 56787 92023 56821 92051
rect 56849 92023 56884 92051
rect 56724 91989 56884 92023
rect 56724 91961 56759 91989
rect 56787 91961 56821 91989
rect 56849 91961 56884 91989
rect 56724 91944 56884 91961
rect 57437 86175 57747 94961
rect 58974 95175 59134 95192
rect 58974 95147 59009 95175
rect 59037 95147 59071 95175
rect 59099 95147 59134 95175
rect 58974 95113 59134 95147
rect 58974 95085 59009 95113
rect 59037 95085 59071 95113
rect 59099 95085 59134 95113
rect 58974 95051 59134 95085
rect 58974 95023 59009 95051
rect 59037 95023 59071 95051
rect 59099 95023 59134 95051
rect 58974 94989 59134 95023
rect 58974 94961 59009 94989
rect 59037 94961 59071 94989
rect 59099 94961 59134 94989
rect 58974 94944 59134 94961
rect 63474 95175 63634 95192
rect 63474 95147 63509 95175
rect 63537 95147 63571 95175
rect 63599 95147 63634 95175
rect 63474 95113 63634 95147
rect 63474 95085 63509 95113
rect 63537 95085 63571 95113
rect 63599 95085 63634 95113
rect 63474 95051 63634 95085
rect 63474 95023 63509 95051
rect 63537 95023 63571 95051
rect 63599 95023 63634 95051
rect 63474 94989 63634 95023
rect 63474 94961 63509 94989
rect 63537 94961 63571 94989
rect 63599 94961 63634 94989
rect 63474 94944 63634 94961
rect 61224 92175 61384 92192
rect 61224 92147 61259 92175
rect 61287 92147 61321 92175
rect 61349 92147 61384 92175
rect 61224 92113 61384 92147
rect 61224 92085 61259 92113
rect 61287 92085 61321 92113
rect 61349 92085 61384 92113
rect 61224 92051 61384 92085
rect 61224 92023 61259 92051
rect 61287 92023 61321 92051
rect 61349 92023 61384 92051
rect 61224 91989 61384 92023
rect 61224 91961 61259 91989
rect 61287 91961 61321 91989
rect 61349 91961 61384 91989
rect 61224 91944 61384 91961
rect 64577 92175 64887 100961
rect 65724 101175 65884 101192
rect 65724 101147 65759 101175
rect 65787 101147 65821 101175
rect 65849 101147 65884 101175
rect 65724 101113 65884 101147
rect 65724 101085 65759 101113
rect 65787 101085 65821 101113
rect 65849 101085 65884 101113
rect 65724 101051 65884 101085
rect 65724 101023 65759 101051
rect 65787 101023 65821 101051
rect 65849 101023 65884 101051
rect 65724 100989 65884 101023
rect 65724 100961 65759 100989
rect 65787 100961 65821 100989
rect 65849 100961 65884 100989
rect 65724 100944 65884 100961
rect 66437 95175 66747 103961
rect 67974 104175 68134 104192
rect 67974 104147 68009 104175
rect 68037 104147 68071 104175
rect 68099 104147 68134 104175
rect 67974 104113 68134 104147
rect 67974 104085 68009 104113
rect 68037 104085 68071 104113
rect 68099 104085 68134 104113
rect 67974 104051 68134 104085
rect 67974 104023 68009 104051
rect 68037 104023 68071 104051
rect 68099 104023 68134 104051
rect 67974 103989 68134 104023
rect 67974 103961 68009 103989
rect 68037 103961 68071 103989
rect 68099 103961 68134 103989
rect 67974 103944 68134 103961
rect 72474 104175 72634 104192
rect 72474 104147 72509 104175
rect 72537 104147 72571 104175
rect 72599 104147 72634 104175
rect 72474 104113 72634 104147
rect 72474 104085 72509 104113
rect 72537 104085 72571 104113
rect 72599 104085 72634 104113
rect 72474 104051 72634 104085
rect 72474 104023 72509 104051
rect 72537 104023 72571 104051
rect 72599 104023 72634 104051
rect 72474 103989 72634 104023
rect 72474 103961 72509 103989
rect 72537 103961 72571 103989
rect 72599 103961 72634 103989
rect 72474 103944 72634 103961
rect 70224 101175 70384 101192
rect 70224 101147 70259 101175
rect 70287 101147 70321 101175
rect 70349 101147 70384 101175
rect 70224 101113 70384 101147
rect 70224 101085 70259 101113
rect 70287 101085 70321 101113
rect 70349 101085 70384 101113
rect 70224 101051 70384 101085
rect 70224 101023 70259 101051
rect 70287 101023 70321 101051
rect 70349 101023 70384 101051
rect 70224 100989 70384 101023
rect 70224 100961 70259 100989
rect 70287 100961 70321 100989
rect 70349 100961 70384 100989
rect 70224 100944 70384 100961
rect 73577 101175 73887 109961
rect 75437 122175 75747 124261
rect 75437 122147 75485 122175
rect 75513 122147 75547 122175
rect 75575 122147 75609 122175
rect 75637 122147 75671 122175
rect 75699 122147 75747 122175
rect 75437 122113 75747 122147
rect 75437 122085 75485 122113
rect 75513 122085 75547 122113
rect 75575 122085 75609 122113
rect 75637 122085 75671 122113
rect 75699 122085 75747 122113
rect 75437 122051 75747 122085
rect 75437 122023 75485 122051
rect 75513 122023 75547 122051
rect 75575 122023 75609 122051
rect 75637 122023 75671 122051
rect 75699 122023 75747 122051
rect 75437 121989 75747 122023
rect 75437 121961 75485 121989
rect 75513 121961 75547 121989
rect 75575 121961 75609 121989
rect 75637 121961 75671 121989
rect 75699 121961 75747 121989
rect 75437 113175 75747 121961
rect 75437 113147 75485 113175
rect 75513 113147 75547 113175
rect 75575 113147 75609 113175
rect 75637 113147 75671 113175
rect 75699 113147 75747 113175
rect 75437 113113 75747 113147
rect 75437 113085 75485 113113
rect 75513 113085 75547 113113
rect 75575 113085 75609 113113
rect 75637 113085 75671 113113
rect 75699 113085 75747 113113
rect 75437 113051 75747 113085
rect 75437 113023 75485 113051
rect 75513 113023 75547 113051
rect 75575 113023 75609 113051
rect 75637 113023 75671 113051
rect 75699 113023 75747 113051
rect 75437 112989 75747 113023
rect 75437 112961 75485 112989
rect 75513 112961 75547 112989
rect 75575 112961 75609 112989
rect 75637 112961 75671 112989
rect 75699 112961 75747 112989
rect 75437 104175 75747 112961
rect 82577 119175 82887 124261
rect 82577 119147 82625 119175
rect 82653 119147 82687 119175
rect 82715 119147 82749 119175
rect 82777 119147 82811 119175
rect 82839 119147 82887 119175
rect 82577 119113 82887 119147
rect 82577 119085 82625 119113
rect 82653 119085 82687 119113
rect 82715 119085 82749 119113
rect 82777 119085 82811 119113
rect 82839 119085 82887 119113
rect 82577 119051 82887 119085
rect 82577 119023 82625 119051
rect 82653 119023 82687 119051
rect 82715 119023 82749 119051
rect 82777 119023 82811 119051
rect 82839 119023 82887 119051
rect 82577 118989 82887 119023
rect 82577 118961 82625 118989
rect 82653 118961 82687 118989
rect 82715 118961 82749 118989
rect 82777 118961 82811 118989
rect 82839 118961 82887 118989
rect 82577 110175 82887 118961
rect 82577 110147 82625 110175
rect 82653 110147 82687 110175
rect 82715 110147 82749 110175
rect 82777 110147 82811 110175
rect 82839 110147 82887 110175
rect 82577 110113 82887 110147
rect 82577 110085 82625 110113
rect 82653 110085 82687 110113
rect 82715 110085 82749 110113
rect 82777 110085 82811 110113
rect 82839 110085 82887 110113
rect 82577 110051 82887 110085
rect 82577 110023 82625 110051
rect 82653 110023 82687 110051
rect 82715 110023 82749 110051
rect 82777 110023 82811 110051
rect 82839 110023 82887 110051
rect 82577 109989 82887 110023
rect 82577 109961 82625 109989
rect 82653 109961 82687 109989
rect 82715 109961 82749 109989
rect 82777 109961 82811 109989
rect 82839 109961 82887 109989
rect 75437 104147 75485 104175
rect 75513 104147 75547 104175
rect 75575 104147 75609 104175
rect 75637 104147 75671 104175
rect 75699 104147 75747 104175
rect 75437 104113 75747 104147
rect 75437 104085 75485 104113
rect 75513 104085 75547 104113
rect 75575 104085 75609 104113
rect 75637 104085 75671 104113
rect 75699 104085 75747 104113
rect 75437 104051 75747 104085
rect 75437 104023 75485 104051
rect 75513 104023 75547 104051
rect 75575 104023 75609 104051
rect 75637 104023 75671 104051
rect 75699 104023 75747 104051
rect 75437 103989 75747 104023
rect 75437 103961 75485 103989
rect 75513 103961 75547 103989
rect 75575 103961 75609 103989
rect 75637 103961 75671 103989
rect 75699 103961 75747 103989
rect 73577 101147 73625 101175
rect 73653 101147 73687 101175
rect 73715 101147 73749 101175
rect 73777 101147 73811 101175
rect 73839 101147 73887 101175
rect 73577 101113 73887 101147
rect 73577 101085 73625 101113
rect 73653 101085 73687 101113
rect 73715 101085 73749 101113
rect 73777 101085 73811 101113
rect 73839 101085 73887 101113
rect 73577 101051 73887 101085
rect 73577 101023 73625 101051
rect 73653 101023 73687 101051
rect 73715 101023 73749 101051
rect 73777 101023 73811 101051
rect 73839 101023 73887 101051
rect 73577 100989 73887 101023
rect 73577 100961 73625 100989
rect 73653 100961 73687 100989
rect 73715 100961 73749 100989
rect 73777 100961 73811 100989
rect 73839 100961 73887 100989
rect 66437 95147 66485 95175
rect 66513 95147 66547 95175
rect 66575 95147 66609 95175
rect 66637 95147 66671 95175
rect 66699 95147 66747 95175
rect 66437 95113 66747 95147
rect 66437 95085 66485 95113
rect 66513 95085 66547 95113
rect 66575 95085 66609 95113
rect 66637 95085 66671 95113
rect 66699 95085 66747 95113
rect 66437 95051 66747 95085
rect 66437 95023 66485 95051
rect 66513 95023 66547 95051
rect 66575 95023 66609 95051
rect 66637 95023 66671 95051
rect 66699 95023 66747 95051
rect 66437 94989 66747 95023
rect 66437 94961 66485 94989
rect 66513 94961 66547 94989
rect 66575 94961 66609 94989
rect 66637 94961 66671 94989
rect 66699 94961 66747 94989
rect 64577 92147 64625 92175
rect 64653 92147 64687 92175
rect 64715 92147 64749 92175
rect 64777 92147 64811 92175
rect 64839 92147 64887 92175
rect 64577 92113 64887 92147
rect 64577 92085 64625 92113
rect 64653 92085 64687 92113
rect 64715 92085 64749 92113
rect 64777 92085 64811 92113
rect 64839 92085 64887 92113
rect 64577 92051 64887 92085
rect 64577 92023 64625 92051
rect 64653 92023 64687 92051
rect 64715 92023 64749 92051
rect 64777 92023 64811 92051
rect 64839 92023 64887 92051
rect 64577 91989 64887 92023
rect 64577 91961 64625 91989
rect 64653 91961 64687 91989
rect 64715 91961 64749 91989
rect 64777 91961 64811 91989
rect 64839 91961 64887 91989
rect 57437 86147 57485 86175
rect 57513 86147 57547 86175
rect 57575 86147 57609 86175
rect 57637 86147 57671 86175
rect 57699 86147 57747 86175
rect 57437 86113 57747 86147
rect 57437 86085 57485 86113
rect 57513 86085 57547 86113
rect 57575 86085 57609 86113
rect 57637 86085 57671 86113
rect 57699 86085 57747 86113
rect 57437 86051 57747 86085
rect 57437 86023 57485 86051
rect 57513 86023 57547 86051
rect 57575 86023 57609 86051
rect 57637 86023 57671 86051
rect 57699 86023 57747 86051
rect 57437 85989 57747 86023
rect 57437 85961 57485 85989
rect 57513 85961 57547 85989
rect 57575 85961 57609 85989
rect 57637 85961 57671 85989
rect 57699 85961 57747 85989
rect 55577 83147 55625 83175
rect 55653 83147 55687 83175
rect 55715 83147 55749 83175
rect 55777 83147 55811 83175
rect 55839 83147 55887 83175
rect 55577 83113 55887 83147
rect 55577 83085 55625 83113
rect 55653 83085 55687 83113
rect 55715 83085 55749 83113
rect 55777 83085 55811 83113
rect 55839 83085 55887 83113
rect 55577 83051 55887 83085
rect 55577 83023 55625 83051
rect 55653 83023 55687 83051
rect 55715 83023 55749 83051
rect 55777 83023 55811 83051
rect 55839 83023 55887 83051
rect 55577 82989 55887 83023
rect 55577 82961 55625 82989
rect 55653 82961 55687 82989
rect 55715 82961 55749 82989
rect 55777 82961 55811 82989
rect 55839 82961 55887 82989
rect 48437 77147 48485 77175
rect 48513 77147 48547 77175
rect 48575 77147 48609 77175
rect 48637 77147 48671 77175
rect 48699 77147 48747 77175
rect 48437 77113 48747 77147
rect 48437 77085 48485 77113
rect 48513 77085 48547 77113
rect 48575 77085 48609 77113
rect 48637 77085 48671 77113
rect 48699 77085 48747 77113
rect 48437 77051 48747 77085
rect 48437 77023 48485 77051
rect 48513 77023 48547 77051
rect 48575 77023 48609 77051
rect 48637 77023 48671 77051
rect 48699 77023 48747 77051
rect 48437 76989 48747 77023
rect 48437 76961 48485 76989
rect 48513 76961 48547 76989
rect 48575 76961 48609 76989
rect 48637 76961 48671 76989
rect 48699 76961 48747 76989
rect 48437 68175 48747 76961
rect 54474 77175 54634 77192
rect 54474 77147 54509 77175
rect 54537 77147 54571 77175
rect 54599 77147 54634 77175
rect 54474 77113 54634 77147
rect 54474 77085 54509 77113
rect 54537 77085 54571 77113
rect 54599 77085 54634 77113
rect 54474 77051 54634 77085
rect 54474 77023 54509 77051
rect 54537 77023 54571 77051
rect 54599 77023 54634 77051
rect 54474 76989 54634 77023
rect 54474 76961 54509 76989
rect 54537 76961 54571 76989
rect 54599 76961 54634 76989
rect 54474 76944 54634 76961
rect 52224 74175 52384 74192
rect 52224 74147 52259 74175
rect 52287 74147 52321 74175
rect 52349 74147 52384 74175
rect 52224 74113 52384 74147
rect 52224 74085 52259 74113
rect 52287 74085 52321 74113
rect 52349 74085 52384 74113
rect 52224 74051 52384 74085
rect 52224 74023 52259 74051
rect 52287 74023 52321 74051
rect 52349 74023 52384 74051
rect 52224 73989 52384 74023
rect 52224 73961 52259 73989
rect 52287 73961 52321 73989
rect 52349 73961 52384 73989
rect 52224 73944 52384 73961
rect 55577 74175 55887 82961
rect 56724 83175 56884 83192
rect 56724 83147 56759 83175
rect 56787 83147 56821 83175
rect 56849 83147 56884 83175
rect 56724 83113 56884 83147
rect 56724 83085 56759 83113
rect 56787 83085 56821 83113
rect 56849 83085 56884 83113
rect 56724 83051 56884 83085
rect 56724 83023 56759 83051
rect 56787 83023 56821 83051
rect 56849 83023 56884 83051
rect 56724 82989 56884 83023
rect 56724 82961 56759 82989
rect 56787 82961 56821 82989
rect 56849 82961 56884 82989
rect 56724 82944 56884 82961
rect 57437 77175 57747 85961
rect 58974 86175 59134 86192
rect 58974 86147 59009 86175
rect 59037 86147 59071 86175
rect 59099 86147 59134 86175
rect 58974 86113 59134 86147
rect 58974 86085 59009 86113
rect 59037 86085 59071 86113
rect 59099 86085 59134 86113
rect 58974 86051 59134 86085
rect 58974 86023 59009 86051
rect 59037 86023 59071 86051
rect 59099 86023 59134 86051
rect 58974 85989 59134 86023
rect 58974 85961 59009 85989
rect 59037 85961 59071 85989
rect 59099 85961 59134 85989
rect 58974 85944 59134 85961
rect 63474 86175 63634 86192
rect 63474 86147 63509 86175
rect 63537 86147 63571 86175
rect 63599 86147 63634 86175
rect 63474 86113 63634 86147
rect 63474 86085 63509 86113
rect 63537 86085 63571 86113
rect 63599 86085 63634 86113
rect 63474 86051 63634 86085
rect 63474 86023 63509 86051
rect 63537 86023 63571 86051
rect 63599 86023 63634 86051
rect 63474 85989 63634 86023
rect 63474 85961 63509 85989
rect 63537 85961 63571 85989
rect 63599 85961 63634 85989
rect 63474 85944 63634 85961
rect 61224 83175 61384 83192
rect 61224 83147 61259 83175
rect 61287 83147 61321 83175
rect 61349 83147 61384 83175
rect 61224 83113 61384 83147
rect 61224 83085 61259 83113
rect 61287 83085 61321 83113
rect 61349 83085 61384 83113
rect 61224 83051 61384 83085
rect 61224 83023 61259 83051
rect 61287 83023 61321 83051
rect 61349 83023 61384 83051
rect 61224 82989 61384 83023
rect 61224 82961 61259 82989
rect 61287 82961 61321 82989
rect 61349 82961 61384 82989
rect 61224 82944 61384 82961
rect 64577 83175 64887 91961
rect 65724 92175 65884 92192
rect 65724 92147 65759 92175
rect 65787 92147 65821 92175
rect 65849 92147 65884 92175
rect 65724 92113 65884 92147
rect 65724 92085 65759 92113
rect 65787 92085 65821 92113
rect 65849 92085 65884 92113
rect 65724 92051 65884 92085
rect 65724 92023 65759 92051
rect 65787 92023 65821 92051
rect 65849 92023 65884 92051
rect 65724 91989 65884 92023
rect 65724 91961 65759 91989
rect 65787 91961 65821 91989
rect 65849 91961 65884 91989
rect 65724 91944 65884 91961
rect 66437 86175 66747 94961
rect 67974 95175 68134 95192
rect 67974 95147 68009 95175
rect 68037 95147 68071 95175
rect 68099 95147 68134 95175
rect 67974 95113 68134 95147
rect 67974 95085 68009 95113
rect 68037 95085 68071 95113
rect 68099 95085 68134 95113
rect 67974 95051 68134 95085
rect 67974 95023 68009 95051
rect 68037 95023 68071 95051
rect 68099 95023 68134 95051
rect 67974 94989 68134 95023
rect 67974 94961 68009 94989
rect 68037 94961 68071 94989
rect 68099 94961 68134 94989
rect 67974 94944 68134 94961
rect 72474 95175 72634 95192
rect 72474 95147 72509 95175
rect 72537 95147 72571 95175
rect 72599 95147 72634 95175
rect 72474 95113 72634 95147
rect 72474 95085 72509 95113
rect 72537 95085 72571 95113
rect 72599 95085 72634 95113
rect 72474 95051 72634 95085
rect 72474 95023 72509 95051
rect 72537 95023 72571 95051
rect 72599 95023 72634 95051
rect 72474 94989 72634 95023
rect 72474 94961 72509 94989
rect 72537 94961 72571 94989
rect 72599 94961 72634 94989
rect 72474 94944 72634 94961
rect 70224 92175 70384 92192
rect 70224 92147 70259 92175
rect 70287 92147 70321 92175
rect 70349 92147 70384 92175
rect 70224 92113 70384 92147
rect 70224 92085 70259 92113
rect 70287 92085 70321 92113
rect 70349 92085 70384 92113
rect 70224 92051 70384 92085
rect 70224 92023 70259 92051
rect 70287 92023 70321 92051
rect 70349 92023 70384 92051
rect 70224 91989 70384 92023
rect 70224 91961 70259 91989
rect 70287 91961 70321 91989
rect 70349 91961 70384 91989
rect 70224 91944 70384 91961
rect 73577 92175 73887 100961
rect 74724 101175 74884 101192
rect 74724 101147 74759 101175
rect 74787 101147 74821 101175
rect 74849 101147 74884 101175
rect 74724 101113 74884 101147
rect 74724 101085 74759 101113
rect 74787 101085 74821 101113
rect 74849 101085 74884 101113
rect 74724 101051 74884 101085
rect 74724 101023 74759 101051
rect 74787 101023 74821 101051
rect 74849 101023 74884 101051
rect 74724 100989 74884 101023
rect 74724 100961 74759 100989
rect 74787 100961 74821 100989
rect 74849 100961 74884 100989
rect 74724 100944 74884 100961
rect 75437 95175 75747 103961
rect 76974 104175 77134 104192
rect 76974 104147 77009 104175
rect 77037 104147 77071 104175
rect 77099 104147 77134 104175
rect 76974 104113 77134 104147
rect 76974 104085 77009 104113
rect 77037 104085 77071 104113
rect 77099 104085 77134 104113
rect 76974 104051 77134 104085
rect 76974 104023 77009 104051
rect 77037 104023 77071 104051
rect 77099 104023 77134 104051
rect 76974 103989 77134 104023
rect 76974 103961 77009 103989
rect 77037 103961 77071 103989
rect 77099 103961 77134 103989
rect 76974 103944 77134 103961
rect 81474 104175 81634 104192
rect 81474 104147 81509 104175
rect 81537 104147 81571 104175
rect 81599 104147 81634 104175
rect 81474 104113 81634 104147
rect 81474 104085 81509 104113
rect 81537 104085 81571 104113
rect 81599 104085 81634 104113
rect 81474 104051 81634 104085
rect 81474 104023 81509 104051
rect 81537 104023 81571 104051
rect 81599 104023 81634 104051
rect 81474 103989 81634 104023
rect 81474 103961 81509 103989
rect 81537 103961 81571 103989
rect 81599 103961 81634 103989
rect 81474 103944 81634 103961
rect 79224 101175 79384 101192
rect 79224 101147 79259 101175
rect 79287 101147 79321 101175
rect 79349 101147 79384 101175
rect 79224 101113 79384 101147
rect 79224 101085 79259 101113
rect 79287 101085 79321 101113
rect 79349 101085 79384 101113
rect 79224 101051 79384 101085
rect 79224 101023 79259 101051
rect 79287 101023 79321 101051
rect 79349 101023 79384 101051
rect 79224 100989 79384 101023
rect 79224 100961 79259 100989
rect 79287 100961 79321 100989
rect 79349 100961 79384 100989
rect 79224 100944 79384 100961
rect 82577 101175 82887 109961
rect 84437 122175 84747 124261
rect 84437 122147 84485 122175
rect 84513 122147 84547 122175
rect 84575 122147 84609 122175
rect 84637 122147 84671 122175
rect 84699 122147 84747 122175
rect 84437 122113 84747 122147
rect 84437 122085 84485 122113
rect 84513 122085 84547 122113
rect 84575 122085 84609 122113
rect 84637 122085 84671 122113
rect 84699 122085 84747 122113
rect 84437 122051 84747 122085
rect 84437 122023 84485 122051
rect 84513 122023 84547 122051
rect 84575 122023 84609 122051
rect 84637 122023 84671 122051
rect 84699 122023 84747 122051
rect 84437 121989 84747 122023
rect 84437 121961 84485 121989
rect 84513 121961 84547 121989
rect 84575 121961 84609 121989
rect 84637 121961 84671 121989
rect 84699 121961 84747 121989
rect 84437 113175 84747 121961
rect 84437 113147 84485 113175
rect 84513 113147 84547 113175
rect 84575 113147 84609 113175
rect 84637 113147 84671 113175
rect 84699 113147 84747 113175
rect 84437 113113 84747 113147
rect 84437 113085 84485 113113
rect 84513 113085 84547 113113
rect 84575 113085 84609 113113
rect 84637 113085 84671 113113
rect 84699 113085 84747 113113
rect 84437 113051 84747 113085
rect 84437 113023 84485 113051
rect 84513 113023 84547 113051
rect 84575 113023 84609 113051
rect 84637 113023 84671 113051
rect 84699 113023 84747 113051
rect 84437 112989 84747 113023
rect 84437 112961 84485 112989
rect 84513 112961 84547 112989
rect 84575 112961 84609 112989
rect 84637 112961 84671 112989
rect 84699 112961 84747 112989
rect 84437 104175 84747 112961
rect 91577 119175 91887 124261
rect 91577 119147 91625 119175
rect 91653 119147 91687 119175
rect 91715 119147 91749 119175
rect 91777 119147 91811 119175
rect 91839 119147 91887 119175
rect 91577 119113 91887 119147
rect 91577 119085 91625 119113
rect 91653 119085 91687 119113
rect 91715 119085 91749 119113
rect 91777 119085 91811 119113
rect 91839 119085 91887 119113
rect 91577 119051 91887 119085
rect 91577 119023 91625 119051
rect 91653 119023 91687 119051
rect 91715 119023 91749 119051
rect 91777 119023 91811 119051
rect 91839 119023 91887 119051
rect 91577 118989 91887 119023
rect 91577 118961 91625 118989
rect 91653 118961 91687 118989
rect 91715 118961 91749 118989
rect 91777 118961 91811 118989
rect 91839 118961 91887 118989
rect 91577 110175 91887 118961
rect 91577 110147 91625 110175
rect 91653 110147 91687 110175
rect 91715 110147 91749 110175
rect 91777 110147 91811 110175
rect 91839 110147 91887 110175
rect 91577 110113 91887 110147
rect 91577 110085 91625 110113
rect 91653 110085 91687 110113
rect 91715 110085 91749 110113
rect 91777 110085 91811 110113
rect 91839 110085 91887 110113
rect 91577 110051 91887 110085
rect 91577 110023 91625 110051
rect 91653 110023 91687 110051
rect 91715 110023 91749 110051
rect 91777 110023 91811 110051
rect 91839 110023 91887 110051
rect 91577 109989 91887 110023
rect 91577 109961 91625 109989
rect 91653 109961 91687 109989
rect 91715 109961 91749 109989
rect 91777 109961 91811 109989
rect 91839 109961 91887 109989
rect 84437 104147 84485 104175
rect 84513 104147 84547 104175
rect 84575 104147 84609 104175
rect 84637 104147 84671 104175
rect 84699 104147 84747 104175
rect 84437 104113 84747 104147
rect 84437 104085 84485 104113
rect 84513 104085 84547 104113
rect 84575 104085 84609 104113
rect 84637 104085 84671 104113
rect 84699 104085 84747 104113
rect 84437 104051 84747 104085
rect 84437 104023 84485 104051
rect 84513 104023 84547 104051
rect 84575 104023 84609 104051
rect 84637 104023 84671 104051
rect 84699 104023 84747 104051
rect 84437 103989 84747 104023
rect 84437 103961 84485 103989
rect 84513 103961 84547 103989
rect 84575 103961 84609 103989
rect 84637 103961 84671 103989
rect 84699 103961 84747 103989
rect 82577 101147 82625 101175
rect 82653 101147 82687 101175
rect 82715 101147 82749 101175
rect 82777 101147 82811 101175
rect 82839 101147 82887 101175
rect 82577 101113 82887 101147
rect 82577 101085 82625 101113
rect 82653 101085 82687 101113
rect 82715 101085 82749 101113
rect 82777 101085 82811 101113
rect 82839 101085 82887 101113
rect 82577 101051 82887 101085
rect 82577 101023 82625 101051
rect 82653 101023 82687 101051
rect 82715 101023 82749 101051
rect 82777 101023 82811 101051
rect 82839 101023 82887 101051
rect 82577 100989 82887 101023
rect 82577 100961 82625 100989
rect 82653 100961 82687 100989
rect 82715 100961 82749 100989
rect 82777 100961 82811 100989
rect 82839 100961 82887 100989
rect 75437 95147 75485 95175
rect 75513 95147 75547 95175
rect 75575 95147 75609 95175
rect 75637 95147 75671 95175
rect 75699 95147 75747 95175
rect 75437 95113 75747 95147
rect 75437 95085 75485 95113
rect 75513 95085 75547 95113
rect 75575 95085 75609 95113
rect 75637 95085 75671 95113
rect 75699 95085 75747 95113
rect 75437 95051 75747 95085
rect 75437 95023 75485 95051
rect 75513 95023 75547 95051
rect 75575 95023 75609 95051
rect 75637 95023 75671 95051
rect 75699 95023 75747 95051
rect 75437 94989 75747 95023
rect 75437 94961 75485 94989
rect 75513 94961 75547 94989
rect 75575 94961 75609 94989
rect 75637 94961 75671 94989
rect 75699 94961 75747 94989
rect 73577 92147 73625 92175
rect 73653 92147 73687 92175
rect 73715 92147 73749 92175
rect 73777 92147 73811 92175
rect 73839 92147 73887 92175
rect 73577 92113 73887 92147
rect 73577 92085 73625 92113
rect 73653 92085 73687 92113
rect 73715 92085 73749 92113
rect 73777 92085 73811 92113
rect 73839 92085 73887 92113
rect 73577 92051 73887 92085
rect 73577 92023 73625 92051
rect 73653 92023 73687 92051
rect 73715 92023 73749 92051
rect 73777 92023 73811 92051
rect 73839 92023 73887 92051
rect 73577 91989 73887 92023
rect 73577 91961 73625 91989
rect 73653 91961 73687 91989
rect 73715 91961 73749 91989
rect 73777 91961 73811 91989
rect 73839 91961 73887 91989
rect 66437 86147 66485 86175
rect 66513 86147 66547 86175
rect 66575 86147 66609 86175
rect 66637 86147 66671 86175
rect 66699 86147 66747 86175
rect 66437 86113 66747 86147
rect 66437 86085 66485 86113
rect 66513 86085 66547 86113
rect 66575 86085 66609 86113
rect 66637 86085 66671 86113
rect 66699 86085 66747 86113
rect 66437 86051 66747 86085
rect 66437 86023 66485 86051
rect 66513 86023 66547 86051
rect 66575 86023 66609 86051
rect 66637 86023 66671 86051
rect 66699 86023 66747 86051
rect 66437 85989 66747 86023
rect 66437 85961 66485 85989
rect 66513 85961 66547 85989
rect 66575 85961 66609 85989
rect 66637 85961 66671 85989
rect 66699 85961 66747 85989
rect 64577 83147 64625 83175
rect 64653 83147 64687 83175
rect 64715 83147 64749 83175
rect 64777 83147 64811 83175
rect 64839 83147 64887 83175
rect 64577 83113 64887 83147
rect 64577 83085 64625 83113
rect 64653 83085 64687 83113
rect 64715 83085 64749 83113
rect 64777 83085 64811 83113
rect 64839 83085 64887 83113
rect 64577 83051 64887 83085
rect 64577 83023 64625 83051
rect 64653 83023 64687 83051
rect 64715 83023 64749 83051
rect 64777 83023 64811 83051
rect 64839 83023 64887 83051
rect 64577 82989 64887 83023
rect 64577 82961 64625 82989
rect 64653 82961 64687 82989
rect 64715 82961 64749 82989
rect 64777 82961 64811 82989
rect 64839 82961 64887 82989
rect 57437 77147 57485 77175
rect 57513 77147 57547 77175
rect 57575 77147 57609 77175
rect 57637 77147 57671 77175
rect 57699 77147 57747 77175
rect 57437 77113 57747 77147
rect 57437 77085 57485 77113
rect 57513 77085 57547 77113
rect 57575 77085 57609 77113
rect 57637 77085 57671 77113
rect 57699 77085 57747 77113
rect 57437 77051 57747 77085
rect 57437 77023 57485 77051
rect 57513 77023 57547 77051
rect 57575 77023 57609 77051
rect 57637 77023 57671 77051
rect 57699 77023 57747 77051
rect 57437 76989 57747 77023
rect 57437 76961 57485 76989
rect 57513 76961 57547 76989
rect 57575 76961 57609 76989
rect 57637 76961 57671 76989
rect 57699 76961 57747 76989
rect 55577 74147 55625 74175
rect 55653 74147 55687 74175
rect 55715 74147 55749 74175
rect 55777 74147 55811 74175
rect 55839 74147 55887 74175
rect 55577 74113 55887 74147
rect 55577 74085 55625 74113
rect 55653 74085 55687 74113
rect 55715 74085 55749 74113
rect 55777 74085 55811 74113
rect 55839 74085 55887 74113
rect 55577 74051 55887 74085
rect 55577 74023 55625 74051
rect 55653 74023 55687 74051
rect 55715 74023 55749 74051
rect 55777 74023 55811 74051
rect 55839 74023 55887 74051
rect 55577 73989 55887 74023
rect 55577 73961 55625 73989
rect 55653 73961 55687 73989
rect 55715 73961 55749 73989
rect 55777 73961 55811 73989
rect 55839 73961 55887 73989
rect 48437 68147 48485 68175
rect 48513 68147 48547 68175
rect 48575 68147 48609 68175
rect 48637 68147 48671 68175
rect 48699 68147 48747 68175
rect 48437 68113 48747 68147
rect 48437 68085 48485 68113
rect 48513 68085 48547 68113
rect 48575 68085 48609 68113
rect 48637 68085 48671 68113
rect 48699 68085 48747 68113
rect 48437 68051 48747 68085
rect 48437 68023 48485 68051
rect 48513 68023 48547 68051
rect 48575 68023 48609 68051
rect 48637 68023 48671 68051
rect 48699 68023 48747 68051
rect 48437 67989 48747 68023
rect 48437 67961 48485 67989
rect 48513 67961 48547 67989
rect 48575 67961 48609 67989
rect 48637 67961 48671 67989
rect 48699 67961 48747 67989
rect 48437 59175 48747 67961
rect 54474 68175 54634 68192
rect 54474 68147 54509 68175
rect 54537 68147 54571 68175
rect 54599 68147 54634 68175
rect 54474 68113 54634 68147
rect 54474 68085 54509 68113
rect 54537 68085 54571 68113
rect 54599 68085 54634 68113
rect 54474 68051 54634 68085
rect 54474 68023 54509 68051
rect 54537 68023 54571 68051
rect 54599 68023 54634 68051
rect 54474 67989 54634 68023
rect 54474 67961 54509 67989
rect 54537 67961 54571 67989
rect 54599 67961 54634 67989
rect 54474 67944 54634 67961
rect 52224 65175 52384 65192
rect 52224 65147 52259 65175
rect 52287 65147 52321 65175
rect 52349 65147 52384 65175
rect 52224 65113 52384 65147
rect 52224 65085 52259 65113
rect 52287 65085 52321 65113
rect 52349 65085 52384 65113
rect 52224 65051 52384 65085
rect 52224 65023 52259 65051
rect 52287 65023 52321 65051
rect 52349 65023 52384 65051
rect 52224 64989 52384 65023
rect 52224 64961 52259 64989
rect 52287 64961 52321 64989
rect 52349 64961 52384 64989
rect 52224 64944 52384 64961
rect 55577 65175 55887 73961
rect 56724 74175 56884 74192
rect 56724 74147 56759 74175
rect 56787 74147 56821 74175
rect 56849 74147 56884 74175
rect 56724 74113 56884 74147
rect 56724 74085 56759 74113
rect 56787 74085 56821 74113
rect 56849 74085 56884 74113
rect 56724 74051 56884 74085
rect 56724 74023 56759 74051
rect 56787 74023 56821 74051
rect 56849 74023 56884 74051
rect 56724 73989 56884 74023
rect 56724 73961 56759 73989
rect 56787 73961 56821 73989
rect 56849 73961 56884 73989
rect 56724 73944 56884 73961
rect 57437 68175 57747 76961
rect 58974 77175 59134 77192
rect 58974 77147 59009 77175
rect 59037 77147 59071 77175
rect 59099 77147 59134 77175
rect 58974 77113 59134 77147
rect 58974 77085 59009 77113
rect 59037 77085 59071 77113
rect 59099 77085 59134 77113
rect 58974 77051 59134 77085
rect 58974 77023 59009 77051
rect 59037 77023 59071 77051
rect 59099 77023 59134 77051
rect 58974 76989 59134 77023
rect 58974 76961 59009 76989
rect 59037 76961 59071 76989
rect 59099 76961 59134 76989
rect 58974 76944 59134 76961
rect 63474 77175 63634 77192
rect 63474 77147 63509 77175
rect 63537 77147 63571 77175
rect 63599 77147 63634 77175
rect 63474 77113 63634 77147
rect 63474 77085 63509 77113
rect 63537 77085 63571 77113
rect 63599 77085 63634 77113
rect 63474 77051 63634 77085
rect 63474 77023 63509 77051
rect 63537 77023 63571 77051
rect 63599 77023 63634 77051
rect 63474 76989 63634 77023
rect 63474 76961 63509 76989
rect 63537 76961 63571 76989
rect 63599 76961 63634 76989
rect 63474 76944 63634 76961
rect 61224 74175 61384 74192
rect 61224 74147 61259 74175
rect 61287 74147 61321 74175
rect 61349 74147 61384 74175
rect 61224 74113 61384 74147
rect 61224 74085 61259 74113
rect 61287 74085 61321 74113
rect 61349 74085 61384 74113
rect 61224 74051 61384 74085
rect 61224 74023 61259 74051
rect 61287 74023 61321 74051
rect 61349 74023 61384 74051
rect 61224 73989 61384 74023
rect 61224 73961 61259 73989
rect 61287 73961 61321 73989
rect 61349 73961 61384 73989
rect 61224 73944 61384 73961
rect 64577 74175 64887 82961
rect 65724 83175 65884 83192
rect 65724 83147 65759 83175
rect 65787 83147 65821 83175
rect 65849 83147 65884 83175
rect 65724 83113 65884 83147
rect 65724 83085 65759 83113
rect 65787 83085 65821 83113
rect 65849 83085 65884 83113
rect 65724 83051 65884 83085
rect 65724 83023 65759 83051
rect 65787 83023 65821 83051
rect 65849 83023 65884 83051
rect 65724 82989 65884 83023
rect 65724 82961 65759 82989
rect 65787 82961 65821 82989
rect 65849 82961 65884 82989
rect 65724 82944 65884 82961
rect 66437 77175 66747 85961
rect 67974 86175 68134 86192
rect 67974 86147 68009 86175
rect 68037 86147 68071 86175
rect 68099 86147 68134 86175
rect 67974 86113 68134 86147
rect 67974 86085 68009 86113
rect 68037 86085 68071 86113
rect 68099 86085 68134 86113
rect 67974 86051 68134 86085
rect 67974 86023 68009 86051
rect 68037 86023 68071 86051
rect 68099 86023 68134 86051
rect 67974 85989 68134 86023
rect 67974 85961 68009 85989
rect 68037 85961 68071 85989
rect 68099 85961 68134 85989
rect 67974 85944 68134 85961
rect 72474 86175 72634 86192
rect 72474 86147 72509 86175
rect 72537 86147 72571 86175
rect 72599 86147 72634 86175
rect 72474 86113 72634 86147
rect 72474 86085 72509 86113
rect 72537 86085 72571 86113
rect 72599 86085 72634 86113
rect 72474 86051 72634 86085
rect 72474 86023 72509 86051
rect 72537 86023 72571 86051
rect 72599 86023 72634 86051
rect 72474 85989 72634 86023
rect 72474 85961 72509 85989
rect 72537 85961 72571 85989
rect 72599 85961 72634 85989
rect 72474 85944 72634 85961
rect 70224 83175 70384 83192
rect 70224 83147 70259 83175
rect 70287 83147 70321 83175
rect 70349 83147 70384 83175
rect 70224 83113 70384 83147
rect 70224 83085 70259 83113
rect 70287 83085 70321 83113
rect 70349 83085 70384 83113
rect 70224 83051 70384 83085
rect 70224 83023 70259 83051
rect 70287 83023 70321 83051
rect 70349 83023 70384 83051
rect 70224 82989 70384 83023
rect 70224 82961 70259 82989
rect 70287 82961 70321 82989
rect 70349 82961 70384 82989
rect 70224 82944 70384 82961
rect 73577 83175 73887 91961
rect 74724 92175 74884 92192
rect 74724 92147 74759 92175
rect 74787 92147 74821 92175
rect 74849 92147 74884 92175
rect 74724 92113 74884 92147
rect 74724 92085 74759 92113
rect 74787 92085 74821 92113
rect 74849 92085 74884 92113
rect 74724 92051 74884 92085
rect 74724 92023 74759 92051
rect 74787 92023 74821 92051
rect 74849 92023 74884 92051
rect 74724 91989 74884 92023
rect 74724 91961 74759 91989
rect 74787 91961 74821 91989
rect 74849 91961 74884 91989
rect 74724 91944 74884 91961
rect 75437 86175 75747 94961
rect 76974 95175 77134 95192
rect 76974 95147 77009 95175
rect 77037 95147 77071 95175
rect 77099 95147 77134 95175
rect 76974 95113 77134 95147
rect 76974 95085 77009 95113
rect 77037 95085 77071 95113
rect 77099 95085 77134 95113
rect 76974 95051 77134 95085
rect 76974 95023 77009 95051
rect 77037 95023 77071 95051
rect 77099 95023 77134 95051
rect 76974 94989 77134 95023
rect 76974 94961 77009 94989
rect 77037 94961 77071 94989
rect 77099 94961 77134 94989
rect 76974 94944 77134 94961
rect 81474 95175 81634 95192
rect 81474 95147 81509 95175
rect 81537 95147 81571 95175
rect 81599 95147 81634 95175
rect 81474 95113 81634 95147
rect 81474 95085 81509 95113
rect 81537 95085 81571 95113
rect 81599 95085 81634 95113
rect 81474 95051 81634 95085
rect 81474 95023 81509 95051
rect 81537 95023 81571 95051
rect 81599 95023 81634 95051
rect 81474 94989 81634 95023
rect 81474 94961 81509 94989
rect 81537 94961 81571 94989
rect 81599 94961 81634 94989
rect 81474 94944 81634 94961
rect 79224 92175 79384 92192
rect 79224 92147 79259 92175
rect 79287 92147 79321 92175
rect 79349 92147 79384 92175
rect 79224 92113 79384 92147
rect 79224 92085 79259 92113
rect 79287 92085 79321 92113
rect 79349 92085 79384 92113
rect 79224 92051 79384 92085
rect 79224 92023 79259 92051
rect 79287 92023 79321 92051
rect 79349 92023 79384 92051
rect 79224 91989 79384 92023
rect 79224 91961 79259 91989
rect 79287 91961 79321 91989
rect 79349 91961 79384 91989
rect 79224 91944 79384 91961
rect 82577 92175 82887 100961
rect 83724 101175 83884 101192
rect 83724 101147 83759 101175
rect 83787 101147 83821 101175
rect 83849 101147 83884 101175
rect 83724 101113 83884 101147
rect 83724 101085 83759 101113
rect 83787 101085 83821 101113
rect 83849 101085 83884 101113
rect 83724 101051 83884 101085
rect 83724 101023 83759 101051
rect 83787 101023 83821 101051
rect 83849 101023 83884 101051
rect 83724 100989 83884 101023
rect 83724 100961 83759 100989
rect 83787 100961 83821 100989
rect 83849 100961 83884 100989
rect 83724 100944 83884 100961
rect 84437 95175 84747 103961
rect 85974 104175 86134 104192
rect 85974 104147 86009 104175
rect 86037 104147 86071 104175
rect 86099 104147 86134 104175
rect 85974 104113 86134 104147
rect 85974 104085 86009 104113
rect 86037 104085 86071 104113
rect 86099 104085 86134 104113
rect 85974 104051 86134 104085
rect 85974 104023 86009 104051
rect 86037 104023 86071 104051
rect 86099 104023 86134 104051
rect 85974 103989 86134 104023
rect 85974 103961 86009 103989
rect 86037 103961 86071 103989
rect 86099 103961 86134 103989
rect 85974 103944 86134 103961
rect 90474 104175 90634 104192
rect 90474 104147 90509 104175
rect 90537 104147 90571 104175
rect 90599 104147 90634 104175
rect 90474 104113 90634 104147
rect 90474 104085 90509 104113
rect 90537 104085 90571 104113
rect 90599 104085 90634 104113
rect 90474 104051 90634 104085
rect 90474 104023 90509 104051
rect 90537 104023 90571 104051
rect 90599 104023 90634 104051
rect 90474 103989 90634 104023
rect 90474 103961 90509 103989
rect 90537 103961 90571 103989
rect 90599 103961 90634 103989
rect 90474 103944 90634 103961
rect 88224 101175 88384 101192
rect 88224 101147 88259 101175
rect 88287 101147 88321 101175
rect 88349 101147 88384 101175
rect 88224 101113 88384 101147
rect 88224 101085 88259 101113
rect 88287 101085 88321 101113
rect 88349 101085 88384 101113
rect 88224 101051 88384 101085
rect 88224 101023 88259 101051
rect 88287 101023 88321 101051
rect 88349 101023 88384 101051
rect 88224 100989 88384 101023
rect 88224 100961 88259 100989
rect 88287 100961 88321 100989
rect 88349 100961 88384 100989
rect 88224 100944 88384 100961
rect 91577 101175 91887 109961
rect 93437 122175 93747 124261
rect 93437 122147 93485 122175
rect 93513 122147 93547 122175
rect 93575 122147 93609 122175
rect 93637 122147 93671 122175
rect 93699 122147 93747 122175
rect 93437 122113 93747 122147
rect 93437 122085 93485 122113
rect 93513 122085 93547 122113
rect 93575 122085 93609 122113
rect 93637 122085 93671 122113
rect 93699 122085 93747 122113
rect 93437 122051 93747 122085
rect 93437 122023 93485 122051
rect 93513 122023 93547 122051
rect 93575 122023 93609 122051
rect 93637 122023 93671 122051
rect 93699 122023 93747 122051
rect 93437 121989 93747 122023
rect 93437 121961 93485 121989
rect 93513 121961 93547 121989
rect 93575 121961 93609 121989
rect 93637 121961 93671 121989
rect 93699 121961 93747 121989
rect 93437 113175 93747 121961
rect 93437 113147 93485 113175
rect 93513 113147 93547 113175
rect 93575 113147 93609 113175
rect 93637 113147 93671 113175
rect 93699 113147 93747 113175
rect 93437 113113 93747 113147
rect 93437 113085 93485 113113
rect 93513 113085 93547 113113
rect 93575 113085 93609 113113
rect 93637 113085 93671 113113
rect 93699 113085 93747 113113
rect 93437 113051 93747 113085
rect 93437 113023 93485 113051
rect 93513 113023 93547 113051
rect 93575 113023 93609 113051
rect 93637 113023 93671 113051
rect 93699 113023 93747 113051
rect 93437 112989 93747 113023
rect 93437 112961 93485 112989
rect 93513 112961 93547 112989
rect 93575 112961 93609 112989
rect 93637 112961 93671 112989
rect 93699 112961 93747 112989
rect 93437 104175 93747 112961
rect 100577 119175 100887 124261
rect 100577 119147 100625 119175
rect 100653 119147 100687 119175
rect 100715 119147 100749 119175
rect 100777 119147 100811 119175
rect 100839 119147 100887 119175
rect 100577 119113 100887 119147
rect 100577 119085 100625 119113
rect 100653 119085 100687 119113
rect 100715 119085 100749 119113
rect 100777 119085 100811 119113
rect 100839 119085 100887 119113
rect 100577 119051 100887 119085
rect 100577 119023 100625 119051
rect 100653 119023 100687 119051
rect 100715 119023 100749 119051
rect 100777 119023 100811 119051
rect 100839 119023 100887 119051
rect 100577 118989 100887 119023
rect 100577 118961 100625 118989
rect 100653 118961 100687 118989
rect 100715 118961 100749 118989
rect 100777 118961 100811 118989
rect 100839 118961 100887 118989
rect 100577 110175 100887 118961
rect 100577 110147 100625 110175
rect 100653 110147 100687 110175
rect 100715 110147 100749 110175
rect 100777 110147 100811 110175
rect 100839 110147 100887 110175
rect 100577 110113 100887 110147
rect 100577 110085 100625 110113
rect 100653 110085 100687 110113
rect 100715 110085 100749 110113
rect 100777 110085 100811 110113
rect 100839 110085 100887 110113
rect 100577 110051 100887 110085
rect 100577 110023 100625 110051
rect 100653 110023 100687 110051
rect 100715 110023 100749 110051
rect 100777 110023 100811 110051
rect 100839 110023 100887 110051
rect 100577 109989 100887 110023
rect 100577 109961 100625 109989
rect 100653 109961 100687 109989
rect 100715 109961 100749 109989
rect 100777 109961 100811 109989
rect 100839 109961 100887 109989
rect 93437 104147 93485 104175
rect 93513 104147 93547 104175
rect 93575 104147 93609 104175
rect 93637 104147 93671 104175
rect 93699 104147 93747 104175
rect 93437 104113 93747 104147
rect 93437 104085 93485 104113
rect 93513 104085 93547 104113
rect 93575 104085 93609 104113
rect 93637 104085 93671 104113
rect 93699 104085 93747 104113
rect 93437 104051 93747 104085
rect 93437 104023 93485 104051
rect 93513 104023 93547 104051
rect 93575 104023 93609 104051
rect 93637 104023 93671 104051
rect 93699 104023 93747 104051
rect 93437 103989 93747 104023
rect 93437 103961 93485 103989
rect 93513 103961 93547 103989
rect 93575 103961 93609 103989
rect 93637 103961 93671 103989
rect 93699 103961 93747 103989
rect 91577 101147 91625 101175
rect 91653 101147 91687 101175
rect 91715 101147 91749 101175
rect 91777 101147 91811 101175
rect 91839 101147 91887 101175
rect 91577 101113 91887 101147
rect 91577 101085 91625 101113
rect 91653 101085 91687 101113
rect 91715 101085 91749 101113
rect 91777 101085 91811 101113
rect 91839 101085 91887 101113
rect 91577 101051 91887 101085
rect 91577 101023 91625 101051
rect 91653 101023 91687 101051
rect 91715 101023 91749 101051
rect 91777 101023 91811 101051
rect 91839 101023 91887 101051
rect 91577 100989 91887 101023
rect 91577 100961 91625 100989
rect 91653 100961 91687 100989
rect 91715 100961 91749 100989
rect 91777 100961 91811 100989
rect 91839 100961 91887 100989
rect 84437 95147 84485 95175
rect 84513 95147 84547 95175
rect 84575 95147 84609 95175
rect 84637 95147 84671 95175
rect 84699 95147 84747 95175
rect 84437 95113 84747 95147
rect 84437 95085 84485 95113
rect 84513 95085 84547 95113
rect 84575 95085 84609 95113
rect 84637 95085 84671 95113
rect 84699 95085 84747 95113
rect 84437 95051 84747 95085
rect 84437 95023 84485 95051
rect 84513 95023 84547 95051
rect 84575 95023 84609 95051
rect 84637 95023 84671 95051
rect 84699 95023 84747 95051
rect 84437 94989 84747 95023
rect 84437 94961 84485 94989
rect 84513 94961 84547 94989
rect 84575 94961 84609 94989
rect 84637 94961 84671 94989
rect 84699 94961 84747 94989
rect 82577 92147 82625 92175
rect 82653 92147 82687 92175
rect 82715 92147 82749 92175
rect 82777 92147 82811 92175
rect 82839 92147 82887 92175
rect 82577 92113 82887 92147
rect 82577 92085 82625 92113
rect 82653 92085 82687 92113
rect 82715 92085 82749 92113
rect 82777 92085 82811 92113
rect 82839 92085 82887 92113
rect 82577 92051 82887 92085
rect 82577 92023 82625 92051
rect 82653 92023 82687 92051
rect 82715 92023 82749 92051
rect 82777 92023 82811 92051
rect 82839 92023 82887 92051
rect 82577 91989 82887 92023
rect 82577 91961 82625 91989
rect 82653 91961 82687 91989
rect 82715 91961 82749 91989
rect 82777 91961 82811 91989
rect 82839 91961 82887 91989
rect 75437 86147 75485 86175
rect 75513 86147 75547 86175
rect 75575 86147 75609 86175
rect 75637 86147 75671 86175
rect 75699 86147 75747 86175
rect 75437 86113 75747 86147
rect 75437 86085 75485 86113
rect 75513 86085 75547 86113
rect 75575 86085 75609 86113
rect 75637 86085 75671 86113
rect 75699 86085 75747 86113
rect 75437 86051 75747 86085
rect 75437 86023 75485 86051
rect 75513 86023 75547 86051
rect 75575 86023 75609 86051
rect 75637 86023 75671 86051
rect 75699 86023 75747 86051
rect 75437 85989 75747 86023
rect 75437 85961 75485 85989
rect 75513 85961 75547 85989
rect 75575 85961 75609 85989
rect 75637 85961 75671 85989
rect 75699 85961 75747 85989
rect 73577 83147 73625 83175
rect 73653 83147 73687 83175
rect 73715 83147 73749 83175
rect 73777 83147 73811 83175
rect 73839 83147 73887 83175
rect 73577 83113 73887 83147
rect 73577 83085 73625 83113
rect 73653 83085 73687 83113
rect 73715 83085 73749 83113
rect 73777 83085 73811 83113
rect 73839 83085 73887 83113
rect 73577 83051 73887 83085
rect 73577 83023 73625 83051
rect 73653 83023 73687 83051
rect 73715 83023 73749 83051
rect 73777 83023 73811 83051
rect 73839 83023 73887 83051
rect 73577 82989 73887 83023
rect 73577 82961 73625 82989
rect 73653 82961 73687 82989
rect 73715 82961 73749 82989
rect 73777 82961 73811 82989
rect 73839 82961 73887 82989
rect 66437 77147 66485 77175
rect 66513 77147 66547 77175
rect 66575 77147 66609 77175
rect 66637 77147 66671 77175
rect 66699 77147 66747 77175
rect 66437 77113 66747 77147
rect 66437 77085 66485 77113
rect 66513 77085 66547 77113
rect 66575 77085 66609 77113
rect 66637 77085 66671 77113
rect 66699 77085 66747 77113
rect 66437 77051 66747 77085
rect 66437 77023 66485 77051
rect 66513 77023 66547 77051
rect 66575 77023 66609 77051
rect 66637 77023 66671 77051
rect 66699 77023 66747 77051
rect 66437 76989 66747 77023
rect 66437 76961 66485 76989
rect 66513 76961 66547 76989
rect 66575 76961 66609 76989
rect 66637 76961 66671 76989
rect 66699 76961 66747 76989
rect 64577 74147 64625 74175
rect 64653 74147 64687 74175
rect 64715 74147 64749 74175
rect 64777 74147 64811 74175
rect 64839 74147 64887 74175
rect 64577 74113 64887 74147
rect 64577 74085 64625 74113
rect 64653 74085 64687 74113
rect 64715 74085 64749 74113
rect 64777 74085 64811 74113
rect 64839 74085 64887 74113
rect 64577 74051 64887 74085
rect 64577 74023 64625 74051
rect 64653 74023 64687 74051
rect 64715 74023 64749 74051
rect 64777 74023 64811 74051
rect 64839 74023 64887 74051
rect 64577 73989 64887 74023
rect 64577 73961 64625 73989
rect 64653 73961 64687 73989
rect 64715 73961 64749 73989
rect 64777 73961 64811 73989
rect 64839 73961 64887 73989
rect 57437 68147 57485 68175
rect 57513 68147 57547 68175
rect 57575 68147 57609 68175
rect 57637 68147 57671 68175
rect 57699 68147 57747 68175
rect 57437 68113 57747 68147
rect 57437 68085 57485 68113
rect 57513 68085 57547 68113
rect 57575 68085 57609 68113
rect 57637 68085 57671 68113
rect 57699 68085 57747 68113
rect 57437 68051 57747 68085
rect 57437 68023 57485 68051
rect 57513 68023 57547 68051
rect 57575 68023 57609 68051
rect 57637 68023 57671 68051
rect 57699 68023 57747 68051
rect 57437 67989 57747 68023
rect 57437 67961 57485 67989
rect 57513 67961 57547 67989
rect 57575 67961 57609 67989
rect 57637 67961 57671 67989
rect 57699 67961 57747 67989
rect 55577 65147 55625 65175
rect 55653 65147 55687 65175
rect 55715 65147 55749 65175
rect 55777 65147 55811 65175
rect 55839 65147 55887 65175
rect 55577 65113 55887 65147
rect 55577 65085 55625 65113
rect 55653 65085 55687 65113
rect 55715 65085 55749 65113
rect 55777 65085 55811 65113
rect 55839 65085 55887 65113
rect 55577 65051 55887 65085
rect 55577 65023 55625 65051
rect 55653 65023 55687 65051
rect 55715 65023 55749 65051
rect 55777 65023 55811 65051
rect 55839 65023 55887 65051
rect 55577 64989 55887 65023
rect 55577 64961 55625 64989
rect 55653 64961 55687 64989
rect 55715 64961 55749 64989
rect 55777 64961 55811 64989
rect 55839 64961 55887 64989
rect 48437 59147 48485 59175
rect 48513 59147 48547 59175
rect 48575 59147 48609 59175
rect 48637 59147 48671 59175
rect 48699 59147 48747 59175
rect 48437 59113 48747 59147
rect 48437 59085 48485 59113
rect 48513 59085 48547 59113
rect 48575 59085 48609 59113
rect 48637 59085 48671 59113
rect 48699 59085 48747 59113
rect 48437 59051 48747 59085
rect 48437 59023 48485 59051
rect 48513 59023 48547 59051
rect 48575 59023 48609 59051
rect 48637 59023 48671 59051
rect 48699 59023 48747 59051
rect 48437 58989 48747 59023
rect 48437 58961 48485 58989
rect 48513 58961 48547 58989
rect 48575 58961 48609 58989
rect 48637 58961 48671 58989
rect 48699 58961 48747 58989
rect 48437 50175 48747 58961
rect 54474 59175 54634 59192
rect 54474 59147 54509 59175
rect 54537 59147 54571 59175
rect 54599 59147 54634 59175
rect 54474 59113 54634 59147
rect 54474 59085 54509 59113
rect 54537 59085 54571 59113
rect 54599 59085 54634 59113
rect 54474 59051 54634 59085
rect 54474 59023 54509 59051
rect 54537 59023 54571 59051
rect 54599 59023 54634 59051
rect 54474 58989 54634 59023
rect 54474 58961 54509 58989
rect 54537 58961 54571 58989
rect 54599 58961 54634 58989
rect 54474 58944 54634 58961
rect 52224 56175 52384 56192
rect 52224 56147 52259 56175
rect 52287 56147 52321 56175
rect 52349 56147 52384 56175
rect 52224 56113 52384 56147
rect 52224 56085 52259 56113
rect 52287 56085 52321 56113
rect 52349 56085 52384 56113
rect 52224 56051 52384 56085
rect 52224 56023 52259 56051
rect 52287 56023 52321 56051
rect 52349 56023 52384 56051
rect 52224 55989 52384 56023
rect 52224 55961 52259 55989
rect 52287 55961 52321 55989
rect 52349 55961 52384 55989
rect 52224 55944 52384 55961
rect 55577 56175 55887 64961
rect 56724 65175 56884 65192
rect 56724 65147 56759 65175
rect 56787 65147 56821 65175
rect 56849 65147 56884 65175
rect 56724 65113 56884 65147
rect 56724 65085 56759 65113
rect 56787 65085 56821 65113
rect 56849 65085 56884 65113
rect 56724 65051 56884 65085
rect 56724 65023 56759 65051
rect 56787 65023 56821 65051
rect 56849 65023 56884 65051
rect 56724 64989 56884 65023
rect 56724 64961 56759 64989
rect 56787 64961 56821 64989
rect 56849 64961 56884 64989
rect 56724 64944 56884 64961
rect 57437 59175 57747 67961
rect 58974 68175 59134 68192
rect 58974 68147 59009 68175
rect 59037 68147 59071 68175
rect 59099 68147 59134 68175
rect 58974 68113 59134 68147
rect 58974 68085 59009 68113
rect 59037 68085 59071 68113
rect 59099 68085 59134 68113
rect 58974 68051 59134 68085
rect 58974 68023 59009 68051
rect 59037 68023 59071 68051
rect 59099 68023 59134 68051
rect 58974 67989 59134 68023
rect 58974 67961 59009 67989
rect 59037 67961 59071 67989
rect 59099 67961 59134 67989
rect 58974 67944 59134 67961
rect 63474 68175 63634 68192
rect 63474 68147 63509 68175
rect 63537 68147 63571 68175
rect 63599 68147 63634 68175
rect 63474 68113 63634 68147
rect 63474 68085 63509 68113
rect 63537 68085 63571 68113
rect 63599 68085 63634 68113
rect 63474 68051 63634 68085
rect 63474 68023 63509 68051
rect 63537 68023 63571 68051
rect 63599 68023 63634 68051
rect 63474 67989 63634 68023
rect 63474 67961 63509 67989
rect 63537 67961 63571 67989
rect 63599 67961 63634 67989
rect 63474 67944 63634 67961
rect 61224 65175 61384 65192
rect 61224 65147 61259 65175
rect 61287 65147 61321 65175
rect 61349 65147 61384 65175
rect 61224 65113 61384 65147
rect 61224 65085 61259 65113
rect 61287 65085 61321 65113
rect 61349 65085 61384 65113
rect 61224 65051 61384 65085
rect 61224 65023 61259 65051
rect 61287 65023 61321 65051
rect 61349 65023 61384 65051
rect 61224 64989 61384 65023
rect 61224 64961 61259 64989
rect 61287 64961 61321 64989
rect 61349 64961 61384 64989
rect 61224 64944 61384 64961
rect 64577 65175 64887 73961
rect 65724 74175 65884 74192
rect 65724 74147 65759 74175
rect 65787 74147 65821 74175
rect 65849 74147 65884 74175
rect 65724 74113 65884 74147
rect 65724 74085 65759 74113
rect 65787 74085 65821 74113
rect 65849 74085 65884 74113
rect 65724 74051 65884 74085
rect 65724 74023 65759 74051
rect 65787 74023 65821 74051
rect 65849 74023 65884 74051
rect 65724 73989 65884 74023
rect 65724 73961 65759 73989
rect 65787 73961 65821 73989
rect 65849 73961 65884 73989
rect 65724 73944 65884 73961
rect 66437 68175 66747 76961
rect 67974 77175 68134 77192
rect 67974 77147 68009 77175
rect 68037 77147 68071 77175
rect 68099 77147 68134 77175
rect 67974 77113 68134 77147
rect 67974 77085 68009 77113
rect 68037 77085 68071 77113
rect 68099 77085 68134 77113
rect 67974 77051 68134 77085
rect 67974 77023 68009 77051
rect 68037 77023 68071 77051
rect 68099 77023 68134 77051
rect 67974 76989 68134 77023
rect 67974 76961 68009 76989
rect 68037 76961 68071 76989
rect 68099 76961 68134 76989
rect 67974 76944 68134 76961
rect 72474 77175 72634 77192
rect 72474 77147 72509 77175
rect 72537 77147 72571 77175
rect 72599 77147 72634 77175
rect 72474 77113 72634 77147
rect 72474 77085 72509 77113
rect 72537 77085 72571 77113
rect 72599 77085 72634 77113
rect 72474 77051 72634 77085
rect 72474 77023 72509 77051
rect 72537 77023 72571 77051
rect 72599 77023 72634 77051
rect 72474 76989 72634 77023
rect 72474 76961 72509 76989
rect 72537 76961 72571 76989
rect 72599 76961 72634 76989
rect 72474 76944 72634 76961
rect 70224 74175 70384 74192
rect 70224 74147 70259 74175
rect 70287 74147 70321 74175
rect 70349 74147 70384 74175
rect 70224 74113 70384 74147
rect 70224 74085 70259 74113
rect 70287 74085 70321 74113
rect 70349 74085 70384 74113
rect 70224 74051 70384 74085
rect 70224 74023 70259 74051
rect 70287 74023 70321 74051
rect 70349 74023 70384 74051
rect 70224 73989 70384 74023
rect 70224 73961 70259 73989
rect 70287 73961 70321 73989
rect 70349 73961 70384 73989
rect 70224 73944 70384 73961
rect 73577 74175 73887 82961
rect 74724 83175 74884 83192
rect 74724 83147 74759 83175
rect 74787 83147 74821 83175
rect 74849 83147 74884 83175
rect 74724 83113 74884 83147
rect 74724 83085 74759 83113
rect 74787 83085 74821 83113
rect 74849 83085 74884 83113
rect 74724 83051 74884 83085
rect 74724 83023 74759 83051
rect 74787 83023 74821 83051
rect 74849 83023 74884 83051
rect 74724 82989 74884 83023
rect 74724 82961 74759 82989
rect 74787 82961 74821 82989
rect 74849 82961 74884 82989
rect 74724 82944 74884 82961
rect 75437 77175 75747 85961
rect 76974 86175 77134 86192
rect 76974 86147 77009 86175
rect 77037 86147 77071 86175
rect 77099 86147 77134 86175
rect 76974 86113 77134 86147
rect 76974 86085 77009 86113
rect 77037 86085 77071 86113
rect 77099 86085 77134 86113
rect 76974 86051 77134 86085
rect 76974 86023 77009 86051
rect 77037 86023 77071 86051
rect 77099 86023 77134 86051
rect 76974 85989 77134 86023
rect 76974 85961 77009 85989
rect 77037 85961 77071 85989
rect 77099 85961 77134 85989
rect 76974 85944 77134 85961
rect 81474 86175 81634 86192
rect 81474 86147 81509 86175
rect 81537 86147 81571 86175
rect 81599 86147 81634 86175
rect 81474 86113 81634 86147
rect 81474 86085 81509 86113
rect 81537 86085 81571 86113
rect 81599 86085 81634 86113
rect 81474 86051 81634 86085
rect 81474 86023 81509 86051
rect 81537 86023 81571 86051
rect 81599 86023 81634 86051
rect 81474 85989 81634 86023
rect 81474 85961 81509 85989
rect 81537 85961 81571 85989
rect 81599 85961 81634 85989
rect 81474 85944 81634 85961
rect 79224 83175 79384 83192
rect 79224 83147 79259 83175
rect 79287 83147 79321 83175
rect 79349 83147 79384 83175
rect 79224 83113 79384 83147
rect 79224 83085 79259 83113
rect 79287 83085 79321 83113
rect 79349 83085 79384 83113
rect 79224 83051 79384 83085
rect 79224 83023 79259 83051
rect 79287 83023 79321 83051
rect 79349 83023 79384 83051
rect 79224 82989 79384 83023
rect 79224 82961 79259 82989
rect 79287 82961 79321 82989
rect 79349 82961 79384 82989
rect 79224 82944 79384 82961
rect 82577 83175 82887 91961
rect 83724 92175 83884 92192
rect 83724 92147 83759 92175
rect 83787 92147 83821 92175
rect 83849 92147 83884 92175
rect 83724 92113 83884 92147
rect 83724 92085 83759 92113
rect 83787 92085 83821 92113
rect 83849 92085 83884 92113
rect 83724 92051 83884 92085
rect 83724 92023 83759 92051
rect 83787 92023 83821 92051
rect 83849 92023 83884 92051
rect 83724 91989 83884 92023
rect 83724 91961 83759 91989
rect 83787 91961 83821 91989
rect 83849 91961 83884 91989
rect 83724 91944 83884 91961
rect 84437 86175 84747 94961
rect 85974 95175 86134 95192
rect 85974 95147 86009 95175
rect 86037 95147 86071 95175
rect 86099 95147 86134 95175
rect 85974 95113 86134 95147
rect 85974 95085 86009 95113
rect 86037 95085 86071 95113
rect 86099 95085 86134 95113
rect 85974 95051 86134 95085
rect 85974 95023 86009 95051
rect 86037 95023 86071 95051
rect 86099 95023 86134 95051
rect 85974 94989 86134 95023
rect 85974 94961 86009 94989
rect 86037 94961 86071 94989
rect 86099 94961 86134 94989
rect 85974 94944 86134 94961
rect 90474 95175 90634 95192
rect 90474 95147 90509 95175
rect 90537 95147 90571 95175
rect 90599 95147 90634 95175
rect 90474 95113 90634 95147
rect 90474 95085 90509 95113
rect 90537 95085 90571 95113
rect 90599 95085 90634 95113
rect 90474 95051 90634 95085
rect 90474 95023 90509 95051
rect 90537 95023 90571 95051
rect 90599 95023 90634 95051
rect 90474 94989 90634 95023
rect 90474 94961 90509 94989
rect 90537 94961 90571 94989
rect 90599 94961 90634 94989
rect 90474 94944 90634 94961
rect 88224 92175 88384 92192
rect 88224 92147 88259 92175
rect 88287 92147 88321 92175
rect 88349 92147 88384 92175
rect 88224 92113 88384 92147
rect 88224 92085 88259 92113
rect 88287 92085 88321 92113
rect 88349 92085 88384 92113
rect 88224 92051 88384 92085
rect 88224 92023 88259 92051
rect 88287 92023 88321 92051
rect 88349 92023 88384 92051
rect 88224 91989 88384 92023
rect 88224 91961 88259 91989
rect 88287 91961 88321 91989
rect 88349 91961 88384 91989
rect 88224 91944 88384 91961
rect 91577 92175 91887 100961
rect 92724 101175 92884 101192
rect 92724 101147 92759 101175
rect 92787 101147 92821 101175
rect 92849 101147 92884 101175
rect 92724 101113 92884 101147
rect 92724 101085 92759 101113
rect 92787 101085 92821 101113
rect 92849 101085 92884 101113
rect 92724 101051 92884 101085
rect 92724 101023 92759 101051
rect 92787 101023 92821 101051
rect 92849 101023 92884 101051
rect 92724 100989 92884 101023
rect 92724 100961 92759 100989
rect 92787 100961 92821 100989
rect 92849 100961 92884 100989
rect 92724 100944 92884 100961
rect 93437 100635 93747 103961
rect 94974 104175 95134 104192
rect 94974 104147 95009 104175
rect 95037 104147 95071 104175
rect 95099 104147 95134 104175
rect 94974 104113 95134 104147
rect 94974 104085 95009 104113
rect 95037 104085 95071 104113
rect 95099 104085 95134 104113
rect 94974 104051 95134 104085
rect 94974 104023 95009 104051
rect 95037 104023 95071 104051
rect 95099 104023 95134 104051
rect 94974 103989 95134 104023
rect 94974 103961 95009 103989
rect 95037 103961 95071 103989
rect 95099 103961 95134 103989
rect 94974 103944 95134 103961
rect 99474 104175 99634 104192
rect 99474 104147 99509 104175
rect 99537 104147 99571 104175
rect 99599 104147 99634 104175
rect 99474 104113 99634 104147
rect 99474 104085 99509 104113
rect 99537 104085 99571 104113
rect 99599 104085 99634 104113
rect 99474 104051 99634 104085
rect 99474 104023 99509 104051
rect 99537 104023 99571 104051
rect 99599 104023 99634 104051
rect 99474 103989 99634 104023
rect 99474 103961 99509 103989
rect 99537 103961 99571 103989
rect 99599 103961 99634 103989
rect 99474 103944 99634 103961
rect 97224 101175 97384 101192
rect 97224 101147 97259 101175
rect 97287 101147 97321 101175
rect 97349 101147 97384 101175
rect 97224 101113 97384 101147
rect 97224 101085 97259 101113
rect 97287 101085 97321 101113
rect 97349 101085 97384 101113
rect 97224 101051 97384 101085
rect 97224 101023 97259 101051
rect 97287 101023 97321 101051
rect 97349 101023 97384 101051
rect 97224 100989 97384 101023
rect 97224 100961 97259 100989
rect 97287 100961 97321 100989
rect 97349 100961 97384 100989
rect 97224 100944 97384 100961
rect 100577 101175 100887 109961
rect 102437 122175 102747 124261
rect 102437 122147 102485 122175
rect 102513 122147 102547 122175
rect 102575 122147 102609 122175
rect 102637 122147 102671 122175
rect 102699 122147 102747 122175
rect 102437 122113 102747 122147
rect 102437 122085 102485 122113
rect 102513 122085 102547 122113
rect 102575 122085 102609 122113
rect 102637 122085 102671 122113
rect 102699 122085 102747 122113
rect 102437 122051 102747 122085
rect 102437 122023 102485 122051
rect 102513 122023 102547 122051
rect 102575 122023 102609 122051
rect 102637 122023 102671 122051
rect 102699 122023 102747 122051
rect 102437 121989 102747 122023
rect 102437 121961 102485 121989
rect 102513 121961 102547 121989
rect 102575 121961 102609 121989
rect 102637 121961 102671 121989
rect 102699 121961 102747 121989
rect 102437 113175 102747 121961
rect 102437 113147 102485 113175
rect 102513 113147 102547 113175
rect 102575 113147 102609 113175
rect 102637 113147 102671 113175
rect 102699 113147 102747 113175
rect 102437 113113 102747 113147
rect 102437 113085 102485 113113
rect 102513 113085 102547 113113
rect 102575 113085 102609 113113
rect 102637 113085 102671 113113
rect 102699 113085 102747 113113
rect 102437 113051 102747 113085
rect 102437 113023 102485 113051
rect 102513 113023 102547 113051
rect 102575 113023 102609 113051
rect 102637 113023 102671 113051
rect 102699 113023 102747 113051
rect 102437 112989 102747 113023
rect 102437 112961 102485 112989
rect 102513 112961 102547 112989
rect 102575 112961 102609 112989
rect 102637 112961 102671 112989
rect 102699 112961 102747 112989
rect 102437 104175 102747 112961
rect 109577 119175 109887 124261
rect 109577 119147 109625 119175
rect 109653 119147 109687 119175
rect 109715 119147 109749 119175
rect 109777 119147 109811 119175
rect 109839 119147 109887 119175
rect 109577 119113 109887 119147
rect 109577 119085 109625 119113
rect 109653 119085 109687 119113
rect 109715 119085 109749 119113
rect 109777 119085 109811 119113
rect 109839 119085 109887 119113
rect 109577 119051 109887 119085
rect 109577 119023 109625 119051
rect 109653 119023 109687 119051
rect 109715 119023 109749 119051
rect 109777 119023 109811 119051
rect 109839 119023 109887 119051
rect 109577 118989 109887 119023
rect 109577 118961 109625 118989
rect 109653 118961 109687 118989
rect 109715 118961 109749 118989
rect 109777 118961 109811 118989
rect 109839 118961 109887 118989
rect 109577 110175 109887 118961
rect 109577 110147 109625 110175
rect 109653 110147 109687 110175
rect 109715 110147 109749 110175
rect 109777 110147 109811 110175
rect 109839 110147 109887 110175
rect 109577 110113 109887 110147
rect 109577 110085 109625 110113
rect 109653 110085 109687 110113
rect 109715 110085 109749 110113
rect 109777 110085 109811 110113
rect 109839 110085 109887 110113
rect 109577 110051 109887 110085
rect 109577 110023 109625 110051
rect 109653 110023 109687 110051
rect 109715 110023 109749 110051
rect 109777 110023 109811 110051
rect 109839 110023 109887 110051
rect 109577 109989 109887 110023
rect 109577 109961 109625 109989
rect 109653 109961 109687 109989
rect 109715 109961 109749 109989
rect 109777 109961 109811 109989
rect 109839 109961 109887 109989
rect 102437 104147 102485 104175
rect 102513 104147 102547 104175
rect 102575 104147 102609 104175
rect 102637 104147 102671 104175
rect 102699 104147 102747 104175
rect 102437 104113 102747 104147
rect 102437 104085 102485 104113
rect 102513 104085 102547 104113
rect 102575 104085 102609 104113
rect 102637 104085 102671 104113
rect 102699 104085 102747 104113
rect 102437 104051 102747 104085
rect 102437 104023 102485 104051
rect 102513 104023 102547 104051
rect 102575 104023 102609 104051
rect 102637 104023 102671 104051
rect 102699 104023 102747 104051
rect 102437 103989 102747 104023
rect 102437 103961 102485 103989
rect 102513 103961 102547 103989
rect 102575 103961 102609 103989
rect 102637 103961 102671 103989
rect 102699 103961 102747 103989
rect 100577 101147 100625 101175
rect 100653 101147 100687 101175
rect 100715 101147 100749 101175
rect 100777 101147 100811 101175
rect 100839 101147 100887 101175
rect 100577 101113 100887 101147
rect 100577 101085 100625 101113
rect 100653 101085 100687 101113
rect 100715 101085 100749 101113
rect 100777 101085 100811 101113
rect 100839 101085 100887 101113
rect 100577 101051 100887 101085
rect 100577 101023 100625 101051
rect 100653 101023 100687 101051
rect 100715 101023 100749 101051
rect 100777 101023 100811 101051
rect 100839 101023 100887 101051
rect 100577 100989 100887 101023
rect 100577 100961 100625 100989
rect 100653 100961 100687 100989
rect 100715 100961 100749 100989
rect 100777 100961 100811 100989
rect 100839 100961 100887 100989
rect 100577 100635 100887 100961
rect 101724 101175 101884 101192
rect 101724 101147 101759 101175
rect 101787 101147 101821 101175
rect 101849 101147 101884 101175
rect 101724 101113 101884 101147
rect 101724 101085 101759 101113
rect 101787 101085 101821 101113
rect 101849 101085 101884 101113
rect 101724 101051 101884 101085
rect 101724 101023 101759 101051
rect 101787 101023 101821 101051
rect 101849 101023 101884 101051
rect 101724 100989 101884 101023
rect 101724 100961 101759 100989
rect 101787 100961 101821 100989
rect 101849 100961 101884 100989
rect 101724 100944 101884 100961
rect 102437 100635 102747 103961
rect 103974 104175 104134 104192
rect 103974 104147 104009 104175
rect 104037 104147 104071 104175
rect 104099 104147 104134 104175
rect 103974 104113 104134 104147
rect 103974 104085 104009 104113
rect 104037 104085 104071 104113
rect 104099 104085 104134 104113
rect 103974 104051 104134 104085
rect 103974 104023 104009 104051
rect 104037 104023 104071 104051
rect 104099 104023 104134 104051
rect 103974 103989 104134 104023
rect 103974 103961 104009 103989
rect 104037 103961 104071 103989
rect 104099 103961 104134 103989
rect 103974 103944 104134 103961
rect 108474 104175 108634 104192
rect 108474 104147 108509 104175
rect 108537 104147 108571 104175
rect 108599 104147 108634 104175
rect 108474 104113 108634 104147
rect 108474 104085 108509 104113
rect 108537 104085 108571 104113
rect 108599 104085 108634 104113
rect 108474 104051 108634 104085
rect 108474 104023 108509 104051
rect 108537 104023 108571 104051
rect 108599 104023 108634 104051
rect 108474 103989 108634 104023
rect 108474 103961 108509 103989
rect 108537 103961 108571 103989
rect 108599 103961 108634 103989
rect 108474 103944 108634 103961
rect 106224 101175 106384 101192
rect 106224 101147 106259 101175
rect 106287 101147 106321 101175
rect 106349 101147 106384 101175
rect 106224 101113 106384 101147
rect 106224 101085 106259 101113
rect 106287 101085 106321 101113
rect 106349 101085 106384 101113
rect 106224 101051 106384 101085
rect 106224 101023 106259 101051
rect 106287 101023 106321 101051
rect 106349 101023 106384 101051
rect 106224 100989 106384 101023
rect 106224 100961 106259 100989
rect 106287 100961 106321 100989
rect 106349 100961 106384 100989
rect 106224 100944 106384 100961
rect 109577 101175 109887 109961
rect 111437 122175 111747 124261
rect 111437 122147 111485 122175
rect 111513 122147 111547 122175
rect 111575 122147 111609 122175
rect 111637 122147 111671 122175
rect 111699 122147 111747 122175
rect 111437 122113 111747 122147
rect 111437 122085 111485 122113
rect 111513 122085 111547 122113
rect 111575 122085 111609 122113
rect 111637 122085 111671 122113
rect 111699 122085 111747 122113
rect 111437 122051 111747 122085
rect 111437 122023 111485 122051
rect 111513 122023 111547 122051
rect 111575 122023 111609 122051
rect 111637 122023 111671 122051
rect 111699 122023 111747 122051
rect 111437 121989 111747 122023
rect 111437 121961 111485 121989
rect 111513 121961 111547 121989
rect 111575 121961 111609 121989
rect 111637 121961 111671 121989
rect 111699 121961 111747 121989
rect 111437 113175 111747 121961
rect 111437 113147 111485 113175
rect 111513 113147 111547 113175
rect 111575 113147 111609 113175
rect 111637 113147 111671 113175
rect 111699 113147 111747 113175
rect 111437 113113 111747 113147
rect 111437 113085 111485 113113
rect 111513 113085 111547 113113
rect 111575 113085 111609 113113
rect 111637 113085 111671 113113
rect 111699 113085 111747 113113
rect 111437 113051 111747 113085
rect 111437 113023 111485 113051
rect 111513 113023 111547 113051
rect 111575 113023 111609 113051
rect 111637 113023 111671 113051
rect 111699 113023 111747 113051
rect 111437 112989 111747 113023
rect 111437 112961 111485 112989
rect 111513 112961 111547 112989
rect 111575 112961 111609 112989
rect 111637 112961 111671 112989
rect 111699 112961 111747 112989
rect 111437 104175 111747 112961
rect 118577 119175 118887 124261
rect 118577 119147 118625 119175
rect 118653 119147 118687 119175
rect 118715 119147 118749 119175
rect 118777 119147 118811 119175
rect 118839 119147 118887 119175
rect 118577 119113 118887 119147
rect 118577 119085 118625 119113
rect 118653 119085 118687 119113
rect 118715 119085 118749 119113
rect 118777 119085 118811 119113
rect 118839 119085 118887 119113
rect 118577 119051 118887 119085
rect 118577 119023 118625 119051
rect 118653 119023 118687 119051
rect 118715 119023 118749 119051
rect 118777 119023 118811 119051
rect 118839 119023 118887 119051
rect 118577 118989 118887 119023
rect 118577 118961 118625 118989
rect 118653 118961 118687 118989
rect 118715 118961 118749 118989
rect 118777 118961 118811 118989
rect 118839 118961 118887 118989
rect 118577 110175 118887 118961
rect 118577 110147 118625 110175
rect 118653 110147 118687 110175
rect 118715 110147 118749 110175
rect 118777 110147 118811 110175
rect 118839 110147 118887 110175
rect 118577 110113 118887 110147
rect 118577 110085 118625 110113
rect 118653 110085 118687 110113
rect 118715 110085 118749 110113
rect 118777 110085 118811 110113
rect 118839 110085 118887 110113
rect 118577 110051 118887 110085
rect 118577 110023 118625 110051
rect 118653 110023 118687 110051
rect 118715 110023 118749 110051
rect 118777 110023 118811 110051
rect 118839 110023 118887 110051
rect 118577 109989 118887 110023
rect 118577 109961 118625 109989
rect 118653 109961 118687 109989
rect 118715 109961 118749 109989
rect 118777 109961 118811 109989
rect 118839 109961 118887 109989
rect 111437 104147 111485 104175
rect 111513 104147 111547 104175
rect 111575 104147 111609 104175
rect 111637 104147 111671 104175
rect 111699 104147 111747 104175
rect 111437 104113 111747 104147
rect 111437 104085 111485 104113
rect 111513 104085 111547 104113
rect 111575 104085 111609 104113
rect 111637 104085 111671 104113
rect 111699 104085 111747 104113
rect 111437 104051 111747 104085
rect 111437 104023 111485 104051
rect 111513 104023 111547 104051
rect 111575 104023 111609 104051
rect 111637 104023 111671 104051
rect 111699 104023 111747 104051
rect 111437 103989 111747 104023
rect 111437 103961 111485 103989
rect 111513 103961 111547 103989
rect 111575 103961 111609 103989
rect 111637 103961 111671 103989
rect 111699 103961 111747 103989
rect 109577 101147 109625 101175
rect 109653 101147 109687 101175
rect 109715 101147 109749 101175
rect 109777 101147 109811 101175
rect 109839 101147 109887 101175
rect 109577 101113 109887 101147
rect 109577 101085 109625 101113
rect 109653 101085 109687 101113
rect 109715 101085 109749 101113
rect 109777 101085 109811 101113
rect 109839 101085 109887 101113
rect 109577 101051 109887 101085
rect 109577 101023 109625 101051
rect 109653 101023 109687 101051
rect 109715 101023 109749 101051
rect 109777 101023 109811 101051
rect 109839 101023 109887 101051
rect 109577 100989 109887 101023
rect 109577 100961 109625 100989
rect 109653 100961 109687 100989
rect 109715 100961 109749 100989
rect 109777 100961 109811 100989
rect 109839 100961 109887 100989
rect 109577 100635 109887 100961
rect 110724 101175 110884 101192
rect 110724 101147 110759 101175
rect 110787 101147 110821 101175
rect 110849 101147 110884 101175
rect 110724 101113 110884 101147
rect 110724 101085 110759 101113
rect 110787 101085 110821 101113
rect 110849 101085 110884 101113
rect 110724 101051 110884 101085
rect 110724 101023 110759 101051
rect 110787 101023 110821 101051
rect 110849 101023 110884 101051
rect 110724 100989 110884 101023
rect 110724 100961 110759 100989
rect 110787 100961 110821 100989
rect 110849 100961 110884 100989
rect 110724 100944 110884 100961
rect 111437 100635 111747 103961
rect 112974 104175 113134 104192
rect 112974 104147 113009 104175
rect 113037 104147 113071 104175
rect 113099 104147 113134 104175
rect 112974 104113 113134 104147
rect 112974 104085 113009 104113
rect 113037 104085 113071 104113
rect 113099 104085 113134 104113
rect 112974 104051 113134 104085
rect 112974 104023 113009 104051
rect 113037 104023 113071 104051
rect 113099 104023 113134 104051
rect 112974 103989 113134 104023
rect 112974 103961 113009 103989
rect 113037 103961 113071 103989
rect 113099 103961 113134 103989
rect 112974 103944 113134 103961
rect 117474 104175 117634 104192
rect 117474 104147 117509 104175
rect 117537 104147 117571 104175
rect 117599 104147 117634 104175
rect 117474 104113 117634 104147
rect 117474 104085 117509 104113
rect 117537 104085 117571 104113
rect 117599 104085 117634 104113
rect 117474 104051 117634 104085
rect 117474 104023 117509 104051
rect 117537 104023 117571 104051
rect 117599 104023 117634 104051
rect 117474 103989 117634 104023
rect 117474 103961 117509 103989
rect 117537 103961 117571 103989
rect 117599 103961 117634 103989
rect 117474 103944 117634 103961
rect 115224 101175 115384 101192
rect 115224 101147 115259 101175
rect 115287 101147 115321 101175
rect 115349 101147 115384 101175
rect 115224 101113 115384 101147
rect 115224 101085 115259 101113
rect 115287 101085 115321 101113
rect 115349 101085 115384 101113
rect 115224 101051 115384 101085
rect 115224 101023 115259 101051
rect 115287 101023 115321 101051
rect 115349 101023 115384 101051
rect 115224 100989 115384 101023
rect 115224 100961 115259 100989
rect 115287 100961 115321 100989
rect 115349 100961 115384 100989
rect 115224 100944 115384 100961
rect 118577 101175 118887 109961
rect 118577 101147 118625 101175
rect 118653 101147 118687 101175
rect 118715 101147 118749 101175
rect 118777 101147 118811 101175
rect 118839 101147 118887 101175
rect 118577 101113 118887 101147
rect 118577 101085 118625 101113
rect 118653 101085 118687 101113
rect 118715 101085 118749 101113
rect 118777 101085 118811 101113
rect 118839 101085 118887 101113
rect 118577 101051 118887 101085
rect 118577 101023 118625 101051
rect 118653 101023 118687 101051
rect 118715 101023 118749 101051
rect 118777 101023 118811 101051
rect 118839 101023 118887 101051
rect 118577 100989 118887 101023
rect 118577 100961 118625 100989
rect 118653 100961 118687 100989
rect 118715 100961 118749 100989
rect 118777 100961 118811 100989
rect 118839 100961 118887 100989
rect 118577 100635 118887 100961
rect 120437 122175 120747 124261
rect 120437 122147 120485 122175
rect 120513 122147 120547 122175
rect 120575 122147 120609 122175
rect 120637 122147 120671 122175
rect 120699 122147 120747 122175
rect 120437 122113 120747 122147
rect 120437 122085 120485 122113
rect 120513 122085 120547 122113
rect 120575 122085 120609 122113
rect 120637 122085 120671 122113
rect 120699 122085 120747 122113
rect 120437 122051 120747 122085
rect 120437 122023 120485 122051
rect 120513 122023 120547 122051
rect 120575 122023 120609 122051
rect 120637 122023 120671 122051
rect 120699 122023 120747 122051
rect 120437 121989 120747 122023
rect 120437 121961 120485 121989
rect 120513 121961 120547 121989
rect 120575 121961 120609 121989
rect 120637 121961 120671 121989
rect 120699 121961 120747 121989
rect 120437 113175 120747 121961
rect 120437 113147 120485 113175
rect 120513 113147 120547 113175
rect 120575 113147 120609 113175
rect 120637 113147 120671 113175
rect 120699 113147 120747 113175
rect 120437 113113 120747 113147
rect 120437 113085 120485 113113
rect 120513 113085 120547 113113
rect 120575 113085 120609 113113
rect 120637 113085 120671 113113
rect 120699 113085 120747 113113
rect 120437 113051 120747 113085
rect 120437 113023 120485 113051
rect 120513 113023 120547 113051
rect 120575 113023 120609 113051
rect 120637 113023 120671 113051
rect 120699 113023 120747 113051
rect 120437 112989 120747 113023
rect 120437 112961 120485 112989
rect 120513 112961 120547 112989
rect 120575 112961 120609 112989
rect 120637 112961 120671 112989
rect 120699 112961 120747 112989
rect 120437 104175 120747 112961
rect 120437 104147 120485 104175
rect 120513 104147 120547 104175
rect 120575 104147 120609 104175
rect 120637 104147 120671 104175
rect 120699 104147 120747 104175
rect 120437 104113 120747 104147
rect 120437 104085 120485 104113
rect 120513 104085 120547 104113
rect 120575 104085 120609 104113
rect 120637 104085 120671 104113
rect 120699 104085 120747 104113
rect 120437 104051 120747 104085
rect 120437 104023 120485 104051
rect 120513 104023 120547 104051
rect 120575 104023 120609 104051
rect 120637 104023 120671 104051
rect 120699 104023 120747 104051
rect 120437 103989 120747 104023
rect 120437 103961 120485 103989
rect 120513 103961 120547 103989
rect 120575 103961 120609 103989
rect 120637 103961 120671 103989
rect 120699 103961 120747 103989
rect 94974 95175 95134 95192
rect 94974 95147 95009 95175
rect 95037 95147 95071 95175
rect 95099 95147 95134 95175
rect 94974 95113 95134 95147
rect 94974 95085 95009 95113
rect 95037 95085 95071 95113
rect 95099 95085 95134 95113
rect 94974 95051 95134 95085
rect 94974 95023 95009 95051
rect 95037 95023 95071 95051
rect 95099 95023 95134 95051
rect 94974 94989 95134 95023
rect 94974 94961 95009 94989
rect 95037 94961 95071 94989
rect 95099 94961 95134 94989
rect 94974 94944 95134 94961
rect 99474 95175 99634 95192
rect 99474 95147 99509 95175
rect 99537 95147 99571 95175
rect 99599 95147 99634 95175
rect 99474 95113 99634 95147
rect 99474 95085 99509 95113
rect 99537 95085 99571 95113
rect 99599 95085 99634 95113
rect 99474 95051 99634 95085
rect 99474 95023 99509 95051
rect 99537 95023 99571 95051
rect 99599 95023 99634 95051
rect 99474 94989 99634 95023
rect 99474 94961 99509 94989
rect 99537 94961 99571 94989
rect 99599 94961 99634 94989
rect 99474 94944 99634 94961
rect 103974 95175 104134 95192
rect 103974 95147 104009 95175
rect 104037 95147 104071 95175
rect 104099 95147 104134 95175
rect 103974 95113 104134 95147
rect 103974 95085 104009 95113
rect 104037 95085 104071 95113
rect 104099 95085 104134 95113
rect 103974 95051 104134 95085
rect 103974 95023 104009 95051
rect 104037 95023 104071 95051
rect 104099 95023 104134 95051
rect 103974 94989 104134 95023
rect 103974 94961 104009 94989
rect 104037 94961 104071 94989
rect 104099 94961 104134 94989
rect 103974 94944 104134 94961
rect 108474 95175 108634 95192
rect 108474 95147 108509 95175
rect 108537 95147 108571 95175
rect 108599 95147 108634 95175
rect 108474 95113 108634 95147
rect 108474 95085 108509 95113
rect 108537 95085 108571 95113
rect 108599 95085 108634 95113
rect 108474 95051 108634 95085
rect 108474 95023 108509 95051
rect 108537 95023 108571 95051
rect 108599 95023 108634 95051
rect 108474 94989 108634 95023
rect 108474 94961 108509 94989
rect 108537 94961 108571 94989
rect 108599 94961 108634 94989
rect 108474 94944 108634 94961
rect 112974 95175 113134 95192
rect 112974 95147 113009 95175
rect 113037 95147 113071 95175
rect 113099 95147 113134 95175
rect 112974 95113 113134 95147
rect 112974 95085 113009 95113
rect 113037 95085 113071 95113
rect 113099 95085 113134 95113
rect 112974 95051 113134 95085
rect 112974 95023 113009 95051
rect 113037 95023 113071 95051
rect 113099 95023 113134 95051
rect 112974 94989 113134 95023
rect 112974 94961 113009 94989
rect 113037 94961 113071 94989
rect 113099 94961 113134 94989
rect 112974 94944 113134 94961
rect 117474 95175 117634 95192
rect 117474 95147 117509 95175
rect 117537 95147 117571 95175
rect 117599 95147 117634 95175
rect 117474 95113 117634 95147
rect 117474 95085 117509 95113
rect 117537 95085 117571 95113
rect 117599 95085 117634 95113
rect 117474 95051 117634 95085
rect 117474 95023 117509 95051
rect 117537 95023 117571 95051
rect 117599 95023 117634 95051
rect 117474 94989 117634 95023
rect 117474 94961 117509 94989
rect 117537 94961 117571 94989
rect 117599 94961 117634 94989
rect 117474 94944 117634 94961
rect 120437 95175 120747 103961
rect 120437 95147 120485 95175
rect 120513 95147 120547 95175
rect 120575 95147 120609 95175
rect 120637 95147 120671 95175
rect 120699 95147 120747 95175
rect 120437 95113 120747 95147
rect 120437 95085 120485 95113
rect 120513 95085 120547 95113
rect 120575 95085 120609 95113
rect 120637 95085 120671 95113
rect 120699 95085 120747 95113
rect 120437 95051 120747 95085
rect 120437 95023 120485 95051
rect 120513 95023 120547 95051
rect 120575 95023 120609 95051
rect 120637 95023 120671 95051
rect 120699 95023 120747 95051
rect 120437 94989 120747 95023
rect 120437 94961 120485 94989
rect 120513 94961 120547 94989
rect 120575 94961 120609 94989
rect 120637 94961 120671 94989
rect 120699 94961 120747 94989
rect 91577 92147 91625 92175
rect 91653 92147 91687 92175
rect 91715 92147 91749 92175
rect 91777 92147 91811 92175
rect 91839 92147 91887 92175
rect 91577 92113 91887 92147
rect 91577 92085 91625 92113
rect 91653 92085 91687 92113
rect 91715 92085 91749 92113
rect 91777 92085 91811 92113
rect 91839 92085 91887 92113
rect 91577 92051 91887 92085
rect 91577 92023 91625 92051
rect 91653 92023 91687 92051
rect 91715 92023 91749 92051
rect 91777 92023 91811 92051
rect 91839 92023 91887 92051
rect 91577 91989 91887 92023
rect 91577 91961 91625 91989
rect 91653 91961 91687 91989
rect 91715 91961 91749 91989
rect 91777 91961 91811 91989
rect 91839 91961 91887 91989
rect 84437 86147 84485 86175
rect 84513 86147 84547 86175
rect 84575 86147 84609 86175
rect 84637 86147 84671 86175
rect 84699 86147 84747 86175
rect 84437 86113 84747 86147
rect 84437 86085 84485 86113
rect 84513 86085 84547 86113
rect 84575 86085 84609 86113
rect 84637 86085 84671 86113
rect 84699 86085 84747 86113
rect 84437 86051 84747 86085
rect 84437 86023 84485 86051
rect 84513 86023 84547 86051
rect 84575 86023 84609 86051
rect 84637 86023 84671 86051
rect 84699 86023 84747 86051
rect 84437 85989 84747 86023
rect 84437 85961 84485 85989
rect 84513 85961 84547 85989
rect 84575 85961 84609 85989
rect 84637 85961 84671 85989
rect 84699 85961 84747 85989
rect 82577 83147 82625 83175
rect 82653 83147 82687 83175
rect 82715 83147 82749 83175
rect 82777 83147 82811 83175
rect 82839 83147 82887 83175
rect 82577 83113 82887 83147
rect 82577 83085 82625 83113
rect 82653 83085 82687 83113
rect 82715 83085 82749 83113
rect 82777 83085 82811 83113
rect 82839 83085 82887 83113
rect 82577 83051 82887 83085
rect 82577 83023 82625 83051
rect 82653 83023 82687 83051
rect 82715 83023 82749 83051
rect 82777 83023 82811 83051
rect 82839 83023 82887 83051
rect 82577 82989 82887 83023
rect 82577 82961 82625 82989
rect 82653 82961 82687 82989
rect 82715 82961 82749 82989
rect 82777 82961 82811 82989
rect 82839 82961 82887 82989
rect 75437 77147 75485 77175
rect 75513 77147 75547 77175
rect 75575 77147 75609 77175
rect 75637 77147 75671 77175
rect 75699 77147 75747 77175
rect 75437 77113 75747 77147
rect 75437 77085 75485 77113
rect 75513 77085 75547 77113
rect 75575 77085 75609 77113
rect 75637 77085 75671 77113
rect 75699 77085 75747 77113
rect 75437 77051 75747 77085
rect 75437 77023 75485 77051
rect 75513 77023 75547 77051
rect 75575 77023 75609 77051
rect 75637 77023 75671 77051
rect 75699 77023 75747 77051
rect 75437 76989 75747 77023
rect 75437 76961 75485 76989
rect 75513 76961 75547 76989
rect 75575 76961 75609 76989
rect 75637 76961 75671 76989
rect 75699 76961 75747 76989
rect 73577 74147 73625 74175
rect 73653 74147 73687 74175
rect 73715 74147 73749 74175
rect 73777 74147 73811 74175
rect 73839 74147 73887 74175
rect 73577 74113 73887 74147
rect 73577 74085 73625 74113
rect 73653 74085 73687 74113
rect 73715 74085 73749 74113
rect 73777 74085 73811 74113
rect 73839 74085 73887 74113
rect 73577 74051 73887 74085
rect 73577 74023 73625 74051
rect 73653 74023 73687 74051
rect 73715 74023 73749 74051
rect 73777 74023 73811 74051
rect 73839 74023 73887 74051
rect 73577 73989 73887 74023
rect 73577 73961 73625 73989
rect 73653 73961 73687 73989
rect 73715 73961 73749 73989
rect 73777 73961 73811 73989
rect 73839 73961 73887 73989
rect 66437 68147 66485 68175
rect 66513 68147 66547 68175
rect 66575 68147 66609 68175
rect 66637 68147 66671 68175
rect 66699 68147 66747 68175
rect 66437 68113 66747 68147
rect 66437 68085 66485 68113
rect 66513 68085 66547 68113
rect 66575 68085 66609 68113
rect 66637 68085 66671 68113
rect 66699 68085 66747 68113
rect 66437 68051 66747 68085
rect 66437 68023 66485 68051
rect 66513 68023 66547 68051
rect 66575 68023 66609 68051
rect 66637 68023 66671 68051
rect 66699 68023 66747 68051
rect 66437 67989 66747 68023
rect 66437 67961 66485 67989
rect 66513 67961 66547 67989
rect 66575 67961 66609 67989
rect 66637 67961 66671 67989
rect 66699 67961 66747 67989
rect 64577 65147 64625 65175
rect 64653 65147 64687 65175
rect 64715 65147 64749 65175
rect 64777 65147 64811 65175
rect 64839 65147 64887 65175
rect 64577 65113 64887 65147
rect 64577 65085 64625 65113
rect 64653 65085 64687 65113
rect 64715 65085 64749 65113
rect 64777 65085 64811 65113
rect 64839 65085 64887 65113
rect 64577 65051 64887 65085
rect 64577 65023 64625 65051
rect 64653 65023 64687 65051
rect 64715 65023 64749 65051
rect 64777 65023 64811 65051
rect 64839 65023 64887 65051
rect 64577 64989 64887 65023
rect 64577 64961 64625 64989
rect 64653 64961 64687 64989
rect 64715 64961 64749 64989
rect 64777 64961 64811 64989
rect 64839 64961 64887 64989
rect 57437 59147 57485 59175
rect 57513 59147 57547 59175
rect 57575 59147 57609 59175
rect 57637 59147 57671 59175
rect 57699 59147 57747 59175
rect 57437 59113 57747 59147
rect 57437 59085 57485 59113
rect 57513 59085 57547 59113
rect 57575 59085 57609 59113
rect 57637 59085 57671 59113
rect 57699 59085 57747 59113
rect 57437 59051 57747 59085
rect 57437 59023 57485 59051
rect 57513 59023 57547 59051
rect 57575 59023 57609 59051
rect 57637 59023 57671 59051
rect 57699 59023 57747 59051
rect 57437 58989 57747 59023
rect 57437 58961 57485 58989
rect 57513 58961 57547 58989
rect 57575 58961 57609 58989
rect 57637 58961 57671 58989
rect 57699 58961 57747 58989
rect 55577 56147 55625 56175
rect 55653 56147 55687 56175
rect 55715 56147 55749 56175
rect 55777 56147 55811 56175
rect 55839 56147 55887 56175
rect 55577 56113 55887 56147
rect 55577 56085 55625 56113
rect 55653 56085 55687 56113
rect 55715 56085 55749 56113
rect 55777 56085 55811 56113
rect 55839 56085 55887 56113
rect 55577 56051 55887 56085
rect 55577 56023 55625 56051
rect 55653 56023 55687 56051
rect 55715 56023 55749 56051
rect 55777 56023 55811 56051
rect 55839 56023 55887 56051
rect 55577 55989 55887 56023
rect 55577 55961 55625 55989
rect 55653 55961 55687 55989
rect 55715 55961 55749 55989
rect 55777 55961 55811 55989
rect 55839 55961 55887 55989
rect 48437 50147 48485 50175
rect 48513 50147 48547 50175
rect 48575 50147 48609 50175
rect 48637 50147 48671 50175
rect 48699 50147 48747 50175
rect 48437 50113 48747 50147
rect 48437 50085 48485 50113
rect 48513 50085 48547 50113
rect 48575 50085 48609 50113
rect 48637 50085 48671 50113
rect 48699 50085 48747 50113
rect 48437 50051 48747 50085
rect 48437 50023 48485 50051
rect 48513 50023 48547 50051
rect 48575 50023 48609 50051
rect 48637 50023 48671 50051
rect 48699 50023 48747 50051
rect 48437 49989 48747 50023
rect 48437 49961 48485 49989
rect 48513 49961 48547 49989
rect 48575 49961 48609 49989
rect 48637 49961 48671 49989
rect 48699 49961 48747 49989
rect 48437 41175 48747 49961
rect 48437 41147 48485 41175
rect 48513 41147 48547 41175
rect 48575 41147 48609 41175
rect 48637 41147 48671 41175
rect 48699 41147 48747 41175
rect 48437 41113 48747 41147
rect 48437 41085 48485 41113
rect 48513 41085 48547 41113
rect 48575 41085 48609 41113
rect 48637 41085 48671 41113
rect 48699 41085 48747 41113
rect 48437 41051 48747 41085
rect 48437 41023 48485 41051
rect 48513 41023 48547 41051
rect 48575 41023 48609 41051
rect 48637 41023 48671 41051
rect 48699 41023 48747 41051
rect 48437 40989 48747 41023
rect 48437 40961 48485 40989
rect 48513 40961 48547 40989
rect 48575 40961 48609 40989
rect 48637 40961 48671 40989
rect 48699 40961 48747 40989
rect 48437 32175 48747 40961
rect 48437 32147 48485 32175
rect 48513 32147 48547 32175
rect 48575 32147 48609 32175
rect 48637 32147 48671 32175
rect 48699 32147 48747 32175
rect 48437 32113 48747 32147
rect 48437 32085 48485 32113
rect 48513 32085 48547 32113
rect 48575 32085 48609 32113
rect 48637 32085 48671 32113
rect 48699 32085 48747 32113
rect 48437 32051 48747 32085
rect 48437 32023 48485 32051
rect 48513 32023 48547 32051
rect 48575 32023 48609 32051
rect 48637 32023 48671 32051
rect 48699 32023 48747 32051
rect 48437 31989 48747 32023
rect 48437 31961 48485 31989
rect 48513 31961 48547 31989
rect 48575 31961 48609 31989
rect 48637 31961 48671 31989
rect 48699 31961 48747 31989
rect 48437 23175 48747 31961
rect 48437 23147 48485 23175
rect 48513 23147 48547 23175
rect 48575 23147 48609 23175
rect 48637 23147 48671 23175
rect 48699 23147 48747 23175
rect 48437 23113 48747 23147
rect 48437 23085 48485 23113
rect 48513 23085 48547 23113
rect 48575 23085 48609 23113
rect 48637 23085 48671 23113
rect 48699 23085 48747 23113
rect 48437 23051 48747 23085
rect 48437 23023 48485 23051
rect 48513 23023 48547 23051
rect 48575 23023 48609 23051
rect 48637 23023 48671 23051
rect 48699 23023 48747 23051
rect 48437 22989 48747 23023
rect 48437 22961 48485 22989
rect 48513 22961 48547 22989
rect 48575 22961 48609 22989
rect 48637 22961 48671 22989
rect 48699 22961 48747 22989
rect 48437 14175 48747 22961
rect 48437 14147 48485 14175
rect 48513 14147 48547 14175
rect 48575 14147 48609 14175
rect 48637 14147 48671 14175
rect 48699 14147 48747 14175
rect 48437 14113 48747 14147
rect 48437 14085 48485 14113
rect 48513 14085 48547 14113
rect 48575 14085 48609 14113
rect 48637 14085 48671 14113
rect 48699 14085 48747 14113
rect 48437 14051 48747 14085
rect 48437 14023 48485 14051
rect 48513 14023 48547 14051
rect 48575 14023 48609 14051
rect 48637 14023 48671 14051
rect 48699 14023 48747 14051
rect 48437 13989 48747 14023
rect 48437 13961 48485 13989
rect 48513 13961 48547 13989
rect 48575 13961 48609 13989
rect 48637 13961 48671 13989
rect 48699 13961 48747 13989
rect 48437 5175 48747 13961
rect 48437 5147 48485 5175
rect 48513 5147 48547 5175
rect 48575 5147 48609 5175
rect 48637 5147 48671 5175
rect 48699 5147 48747 5175
rect 48437 5113 48747 5147
rect 48437 5085 48485 5113
rect 48513 5085 48547 5113
rect 48575 5085 48609 5113
rect 48637 5085 48671 5113
rect 48699 5085 48747 5113
rect 48437 5051 48747 5085
rect 48437 5023 48485 5051
rect 48513 5023 48547 5051
rect 48575 5023 48609 5051
rect 48637 5023 48671 5051
rect 48699 5023 48747 5051
rect 48437 4989 48747 5023
rect 48437 4961 48485 4989
rect 48513 4961 48547 4989
rect 48575 4961 48609 4989
rect 48637 4961 48671 4989
rect 48699 4961 48747 4989
rect 48437 -560 48747 4961
rect 48437 -588 48485 -560
rect 48513 -588 48547 -560
rect 48575 -588 48609 -560
rect 48637 -588 48671 -560
rect 48699 -588 48747 -560
rect 48437 -622 48747 -588
rect 48437 -650 48485 -622
rect 48513 -650 48547 -622
rect 48575 -650 48609 -622
rect 48637 -650 48671 -622
rect 48699 -650 48747 -622
rect 48437 -684 48747 -650
rect 48437 -712 48485 -684
rect 48513 -712 48547 -684
rect 48575 -712 48609 -684
rect 48637 -712 48671 -684
rect 48699 -712 48747 -684
rect 48437 -746 48747 -712
rect 48437 -774 48485 -746
rect 48513 -774 48547 -746
rect 48575 -774 48609 -746
rect 48637 -774 48671 -746
rect 48699 -774 48747 -746
rect 48437 -822 48747 -774
rect 55577 47175 55887 55961
rect 56724 56175 56884 56192
rect 56724 56147 56759 56175
rect 56787 56147 56821 56175
rect 56849 56147 56884 56175
rect 56724 56113 56884 56147
rect 56724 56085 56759 56113
rect 56787 56085 56821 56113
rect 56849 56085 56884 56113
rect 56724 56051 56884 56085
rect 56724 56023 56759 56051
rect 56787 56023 56821 56051
rect 56849 56023 56884 56051
rect 56724 55989 56884 56023
rect 56724 55961 56759 55989
rect 56787 55961 56821 55989
rect 56849 55961 56884 55989
rect 56724 55944 56884 55961
rect 55577 47147 55625 47175
rect 55653 47147 55687 47175
rect 55715 47147 55749 47175
rect 55777 47147 55811 47175
rect 55839 47147 55887 47175
rect 55577 47113 55887 47147
rect 55577 47085 55625 47113
rect 55653 47085 55687 47113
rect 55715 47085 55749 47113
rect 55777 47085 55811 47113
rect 55839 47085 55887 47113
rect 55577 47051 55887 47085
rect 55577 47023 55625 47051
rect 55653 47023 55687 47051
rect 55715 47023 55749 47051
rect 55777 47023 55811 47051
rect 55839 47023 55887 47051
rect 55577 46989 55887 47023
rect 55577 46961 55625 46989
rect 55653 46961 55687 46989
rect 55715 46961 55749 46989
rect 55777 46961 55811 46989
rect 55839 46961 55887 46989
rect 55577 38175 55887 46961
rect 55577 38147 55625 38175
rect 55653 38147 55687 38175
rect 55715 38147 55749 38175
rect 55777 38147 55811 38175
rect 55839 38147 55887 38175
rect 55577 38113 55887 38147
rect 55577 38085 55625 38113
rect 55653 38085 55687 38113
rect 55715 38085 55749 38113
rect 55777 38085 55811 38113
rect 55839 38085 55887 38113
rect 55577 38051 55887 38085
rect 55577 38023 55625 38051
rect 55653 38023 55687 38051
rect 55715 38023 55749 38051
rect 55777 38023 55811 38051
rect 55839 38023 55887 38051
rect 55577 37989 55887 38023
rect 55577 37961 55625 37989
rect 55653 37961 55687 37989
rect 55715 37961 55749 37989
rect 55777 37961 55811 37989
rect 55839 37961 55887 37989
rect 55577 29175 55887 37961
rect 55577 29147 55625 29175
rect 55653 29147 55687 29175
rect 55715 29147 55749 29175
rect 55777 29147 55811 29175
rect 55839 29147 55887 29175
rect 55577 29113 55887 29147
rect 55577 29085 55625 29113
rect 55653 29085 55687 29113
rect 55715 29085 55749 29113
rect 55777 29085 55811 29113
rect 55839 29085 55887 29113
rect 55577 29051 55887 29085
rect 55577 29023 55625 29051
rect 55653 29023 55687 29051
rect 55715 29023 55749 29051
rect 55777 29023 55811 29051
rect 55839 29023 55887 29051
rect 55577 28989 55887 29023
rect 55577 28961 55625 28989
rect 55653 28961 55687 28989
rect 55715 28961 55749 28989
rect 55777 28961 55811 28989
rect 55839 28961 55887 28989
rect 55577 20175 55887 28961
rect 55577 20147 55625 20175
rect 55653 20147 55687 20175
rect 55715 20147 55749 20175
rect 55777 20147 55811 20175
rect 55839 20147 55887 20175
rect 55577 20113 55887 20147
rect 55577 20085 55625 20113
rect 55653 20085 55687 20113
rect 55715 20085 55749 20113
rect 55777 20085 55811 20113
rect 55839 20085 55887 20113
rect 55577 20051 55887 20085
rect 55577 20023 55625 20051
rect 55653 20023 55687 20051
rect 55715 20023 55749 20051
rect 55777 20023 55811 20051
rect 55839 20023 55887 20051
rect 55577 19989 55887 20023
rect 55577 19961 55625 19989
rect 55653 19961 55687 19989
rect 55715 19961 55749 19989
rect 55777 19961 55811 19989
rect 55839 19961 55887 19989
rect 55577 11175 55887 19961
rect 55577 11147 55625 11175
rect 55653 11147 55687 11175
rect 55715 11147 55749 11175
rect 55777 11147 55811 11175
rect 55839 11147 55887 11175
rect 55577 11113 55887 11147
rect 55577 11085 55625 11113
rect 55653 11085 55687 11113
rect 55715 11085 55749 11113
rect 55777 11085 55811 11113
rect 55839 11085 55887 11113
rect 55577 11051 55887 11085
rect 55577 11023 55625 11051
rect 55653 11023 55687 11051
rect 55715 11023 55749 11051
rect 55777 11023 55811 11051
rect 55839 11023 55887 11051
rect 55577 10989 55887 11023
rect 55577 10961 55625 10989
rect 55653 10961 55687 10989
rect 55715 10961 55749 10989
rect 55777 10961 55811 10989
rect 55839 10961 55887 10989
rect 55577 2175 55887 10961
rect 55577 2147 55625 2175
rect 55653 2147 55687 2175
rect 55715 2147 55749 2175
rect 55777 2147 55811 2175
rect 55839 2147 55887 2175
rect 55577 2113 55887 2147
rect 55577 2085 55625 2113
rect 55653 2085 55687 2113
rect 55715 2085 55749 2113
rect 55777 2085 55811 2113
rect 55839 2085 55887 2113
rect 55577 2051 55887 2085
rect 55577 2023 55625 2051
rect 55653 2023 55687 2051
rect 55715 2023 55749 2051
rect 55777 2023 55811 2051
rect 55839 2023 55887 2051
rect 55577 1989 55887 2023
rect 55577 1961 55625 1989
rect 55653 1961 55687 1989
rect 55715 1961 55749 1989
rect 55777 1961 55811 1989
rect 55839 1961 55887 1989
rect 55577 -80 55887 1961
rect 55577 -108 55625 -80
rect 55653 -108 55687 -80
rect 55715 -108 55749 -80
rect 55777 -108 55811 -80
rect 55839 -108 55887 -80
rect 55577 -142 55887 -108
rect 55577 -170 55625 -142
rect 55653 -170 55687 -142
rect 55715 -170 55749 -142
rect 55777 -170 55811 -142
rect 55839 -170 55887 -142
rect 55577 -204 55887 -170
rect 55577 -232 55625 -204
rect 55653 -232 55687 -204
rect 55715 -232 55749 -204
rect 55777 -232 55811 -204
rect 55839 -232 55887 -204
rect 55577 -266 55887 -232
rect 55577 -294 55625 -266
rect 55653 -294 55687 -266
rect 55715 -294 55749 -266
rect 55777 -294 55811 -266
rect 55839 -294 55887 -266
rect 55577 -822 55887 -294
rect 57437 50175 57747 58961
rect 58974 59175 59134 59192
rect 58974 59147 59009 59175
rect 59037 59147 59071 59175
rect 59099 59147 59134 59175
rect 58974 59113 59134 59147
rect 58974 59085 59009 59113
rect 59037 59085 59071 59113
rect 59099 59085 59134 59113
rect 58974 59051 59134 59085
rect 58974 59023 59009 59051
rect 59037 59023 59071 59051
rect 59099 59023 59134 59051
rect 58974 58989 59134 59023
rect 58974 58961 59009 58989
rect 59037 58961 59071 58989
rect 59099 58961 59134 58989
rect 58974 58944 59134 58961
rect 63474 59175 63634 59192
rect 63474 59147 63509 59175
rect 63537 59147 63571 59175
rect 63599 59147 63634 59175
rect 63474 59113 63634 59147
rect 63474 59085 63509 59113
rect 63537 59085 63571 59113
rect 63599 59085 63634 59113
rect 63474 59051 63634 59085
rect 63474 59023 63509 59051
rect 63537 59023 63571 59051
rect 63599 59023 63634 59051
rect 63474 58989 63634 59023
rect 63474 58961 63509 58989
rect 63537 58961 63571 58989
rect 63599 58961 63634 58989
rect 63474 58944 63634 58961
rect 61224 56175 61384 56192
rect 61224 56147 61259 56175
rect 61287 56147 61321 56175
rect 61349 56147 61384 56175
rect 61224 56113 61384 56147
rect 61224 56085 61259 56113
rect 61287 56085 61321 56113
rect 61349 56085 61384 56113
rect 61224 56051 61384 56085
rect 61224 56023 61259 56051
rect 61287 56023 61321 56051
rect 61349 56023 61384 56051
rect 61224 55989 61384 56023
rect 61224 55961 61259 55989
rect 61287 55961 61321 55989
rect 61349 55961 61384 55989
rect 61224 55944 61384 55961
rect 64577 56175 64887 64961
rect 65724 65175 65884 65192
rect 65724 65147 65759 65175
rect 65787 65147 65821 65175
rect 65849 65147 65884 65175
rect 65724 65113 65884 65147
rect 65724 65085 65759 65113
rect 65787 65085 65821 65113
rect 65849 65085 65884 65113
rect 65724 65051 65884 65085
rect 65724 65023 65759 65051
rect 65787 65023 65821 65051
rect 65849 65023 65884 65051
rect 65724 64989 65884 65023
rect 65724 64961 65759 64989
rect 65787 64961 65821 64989
rect 65849 64961 65884 64989
rect 65724 64944 65884 64961
rect 66437 59175 66747 67961
rect 67974 68175 68134 68192
rect 67974 68147 68009 68175
rect 68037 68147 68071 68175
rect 68099 68147 68134 68175
rect 67974 68113 68134 68147
rect 67974 68085 68009 68113
rect 68037 68085 68071 68113
rect 68099 68085 68134 68113
rect 67974 68051 68134 68085
rect 67974 68023 68009 68051
rect 68037 68023 68071 68051
rect 68099 68023 68134 68051
rect 67974 67989 68134 68023
rect 67974 67961 68009 67989
rect 68037 67961 68071 67989
rect 68099 67961 68134 67989
rect 67974 67944 68134 67961
rect 72474 68175 72634 68192
rect 72474 68147 72509 68175
rect 72537 68147 72571 68175
rect 72599 68147 72634 68175
rect 72474 68113 72634 68147
rect 72474 68085 72509 68113
rect 72537 68085 72571 68113
rect 72599 68085 72634 68113
rect 72474 68051 72634 68085
rect 72474 68023 72509 68051
rect 72537 68023 72571 68051
rect 72599 68023 72634 68051
rect 72474 67989 72634 68023
rect 72474 67961 72509 67989
rect 72537 67961 72571 67989
rect 72599 67961 72634 67989
rect 72474 67944 72634 67961
rect 70224 65175 70384 65192
rect 70224 65147 70259 65175
rect 70287 65147 70321 65175
rect 70349 65147 70384 65175
rect 70224 65113 70384 65147
rect 70224 65085 70259 65113
rect 70287 65085 70321 65113
rect 70349 65085 70384 65113
rect 70224 65051 70384 65085
rect 70224 65023 70259 65051
rect 70287 65023 70321 65051
rect 70349 65023 70384 65051
rect 70224 64989 70384 65023
rect 70224 64961 70259 64989
rect 70287 64961 70321 64989
rect 70349 64961 70384 64989
rect 70224 64944 70384 64961
rect 73577 65175 73887 73961
rect 74724 74175 74884 74192
rect 74724 74147 74759 74175
rect 74787 74147 74821 74175
rect 74849 74147 74884 74175
rect 74724 74113 74884 74147
rect 74724 74085 74759 74113
rect 74787 74085 74821 74113
rect 74849 74085 74884 74113
rect 74724 74051 74884 74085
rect 74724 74023 74759 74051
rect 74787 74023 74821 74051
rect 74849 74023 74884 74051
rect 74724 73989 74884 74023
rect 74724 73961 74759 73989
rect 74787 73961 74821 73989
rect 74849 73961 74884 73989
rect 74724 73944 74884 73961
rect 75437 68175 75747 76961
rect 76974 77175 77134 77192
rect 76974 77147 77009 77175
rect 77037 77147 77071 77175
rect 77099 77147 77134 77175
rect 76974 77113 77134 77147
rect 76974 77085 77009 77113
rect 77037 77085 77071 77113
rect 77099 77085 77134 77113
rect 76974 77051 77134 77085
rect 76974 77023 77009 77051
rect 77037 77023 77071 77051
rect 77099 77023 77134 77051
rect 76974 76989 77134 77023
rect 76974 76961 77009 76989
rect 77037 76961 77071 76989
rect 77099 76961 77134 76989
rect 76974 76944 77134 76961
rect 81474 77175 81634 77192
rect 81474 77147 81509 77175
rect 81537 77147 81571 77175
rect 81599 77147 81634 77175
rect 81474 77113 81634 77147
rect 81474 77085 81509 77113
rect 81537 77085 81571 77113
rect 81599 77085 81634 77113
rect 81474 77051 81634 77085
rect 81474 77023 81509 77051
rect 81537 77023 81571 77051
rect 81599 77023 81634 77051
rect 81474 76989 81634 77023
rect 81474 76961 81509 76989
rect 81537 76961 81571 76989
rect 81599 76961 81634 76989
rect 81474 76944 81634 76961
rect 79224 74175 79384 74192
rect 79224 74147 79259 74175
rect 79287 74147 79321 74175
rect 79349 74147 79384 74175
rect 79224 74113 79384 74147
rect 79224 74085 79259 74113
rect 79287 74085 79321 74113
rect 79349 74085 79384 74113
rect 79224 74051 79384 74085
rect 79224 74023 79259 74051
rect 79287 74023 79321 74051
rect 79349 74023 79384 74051
rect 79224 73989 79384 74023
rect 79224 73961 79259 73989
rect 79287 73961 79321 73989
rect 79349 73961 79384 73989
rect 79224 73944 79384 73961
rect 82577 74175 82887 82961
rect 83724 83175 83884 83192
rect 83724 83147 83759 83175
rect 83787 83147 83821 83175
rect 83849 83147 83884 83175
rect 83724 83113 83884 83147
rect 83724 83085 83759 83113
rect 83787 83085 83821 83113
rect 83849 83085 83884 83113
rect 83724 83051 83884 83085
rect 83724 83023 83759 83051
rect 83787 83023 83821 83051
rect 83849 83023 83884 83051
rect 83724 82989 83884 83023
rect 83724 82961 83759 82989
rect 83787 82961 83821 82989
rect 83849 82961 83884 82989
rect 83724 82944 83884 82961
rect 84437 77175 84747 85961
rect 85974 86175 86134 86192
rect 85974 86147 86009 86175
rect 86037 86147 86071 86175
rect 86099 86147 86134 86175
rect 85974 86113 86134 86147
rect 85974 86085 86009 86113
rect 86037 86085 86071 86113
rect 86099 86085 86134 86113
rect 85974 86051 86134 86085
rect 85974 86023 86009 86051
rect 86037 86023 86071 86051
rect 86099 86023 86134 86051
rect 85974 85989 86134 86023
rect 85974 85961 86009 85989
rect 86037 85961 86071 85989
rect 86099 85961 86134 85989
rect 85974 85944 86134 85961
rect 90474 86175 90634 86192
rect 90474 86147 90509 86175
rect 90537 86147 90571 86175
rect 90599 86147 90634 86175
rect 90474 86113 90634 86147
rect 90474 86085 90509 86113
rect 90537 86085 90571 86113
rect 90599 86085 90634 86113
rect 90474 86051 90634 86085
rect 90474 86023 90509 86051
rect 90537 86023 90571 86051
rect 90599 86023 90634 86051
rect 90474 85989 90634 86023
rect 90474 85961 90509 85989
rect 90537 85961 90571 85989
rect 90599 85961 90634 85989
rect 90474 85944 90634 85961
rect 88224 83175 88384 83192
rect 88224 83147 88259 83175
rect 88287 83147 88321 83175
rect 88349 83147 88384 83175
rect 88224 83113 88384 83147
rect 88224 83085 88259 83113
rect 88287 83085 88321 83113
rect 88349 83085 88384 83113
rect 88224 83051 88384 83085
rect 88224 83023 88259 83051
rect 88287 83023 88321 83051
rect 88349 83023 88384 83051
rect 88224 82989 88384 83023
rect 88224 82961 88259 82989
rect 88287 82961 88321 82989
rect 88349 82961 88384 82989
rect 88224 82944 88384 82961
rect 91577 83175 91887 91961
rect 92724 92175 92884 92192
rect 92724 92147 92759 92175
rect 92787 92147 92821 92175
rect 92849 92147 92884 92175
rect 92724 92113 92884 92147
rect 92724 92085 92759 92113
rect 92787 92085 92821 92113
rect 92849 92085 92884 92113
rect 92724 92051 92884 92085
rect 92724 92023 92759 92051
rect 92787 92023 92821 92051
rect 92849 92023 92884 92051
rect 92724 91989 92884 92023
rect 92724 91961 92759 91989
rect 92787 91961 92821 91989
rect 92849 91961 92884 91989
rect 92724 91944 92884 91961
rect 97224 92175 97384 92192
rect 97224 92147 97259 92175
rect 97287 92147 97321 92175
rect 97349 92147 97384 92175
rect 97224 92113 97384 92147
rect 97224 92085 97259 92113
rect 97287 92085 97321 92113
rect 97349 92085 97384 92113
rect 97224 92051 97384 92085
rect 97224 92023 97259 92051
rect 97287 92023 97321 92051
rect 97349 92023 97384 92051
rect 97224 91989 97384 92023
rect 97224 91961 97259 91989
rect 97287 91961 97321 91989
rect 97349 91961 97384 91989
rect 97224 91944 97384 91961
rect 101724 92175 101884 92192
rect 101724 92147 101759 92175
rect 101787 92147 101821 92175
rect 101849 92147 101884 92175
rect 101724 92113 101884 92147
rect 101724 92085 101759 92113
rect 101787 92085 101821 92113
rect 101849 92085 101884 92113
rect 101724 92051 101884 92085
rect 101724 92023 101759 92051
rect 101787 92023 101821 92051
rect 101849 92023 101884 92051
rect 101724 91989 101884 92023
rect 101724 91961 101759 91989
rect 101787 91961 101821 91989
rect 101849 91961 101884 91989
rect 101724 91944 101884 91961
rect 106224 92175 106384 92192
rect 106224 92147 106259 92175
rect 106287 92147 106321 92175
rect 106349 92147 106384 92175
rect 106224 92113 106384 92147
rect 106224 92085 106259 92113
rect 106287 92085 106321 92113
rect 106349 92085 106384 92113
rect 106224 92051 106384 92085
rect 106224 92023 106259 92051
rect 106287 92023 106321 92051
rect 106349 92023 106384 92051
rect 106224 91989 106384 92023
rect 106224 91961 106259 91989
rect 106287 91961 106321 91989
rect 106349 91961 106384 91989
rect 106224 91944 106384 91961
rect 110724 92175 110884 92192
rect 110724 92147 110759 92175
rect 110787 92147 110821 92175
rect 110849 92147 110884 92175
rect 110724 92113 110884 92147
rect 110724 92085 110759 92113
rect 110787 92085 110821 92113
rect 110849 92085 110884 92113
rect 110724 92051 110884 92085
rect 110724 92023 110759 92051
rect 110787 92023 110821 92051
rect 110849 92023 110884 92051
rect 110724 91989 110884 92023
rect 110724 91961 110759 91989
rect 110787 91961 110821 91989
rect 110849 91961 110884 91989
rect 110724 91944 110884 91961
rect 115224 92175 115384 92192
rect 115224 92147 115259 92175
rect 115287 92147 115321 92175
rect 115349 92147 115384 92175
rect 115224 92113 115384 92147
rect 115224 92085 115259 92113
rect 115287 92085 115321 92113
rect 115349 92085 115384 92113
rect 115224 92051 115384 92085
rect 115224 92023 115259 92051
rect 115287 92023 115321 92051
rect 115349 92023 115384 92051
rect 115224 91989 115384 92023
rect 115224 91961 115259 91989
rect 115287 91961 115321 91989
rect 115349 91961 115384 91989
rect 115224 91944 115384 91961
rect 94974 86175 95134 86192
rect 94974 86147 95009 86175
rect 95037 86147 95071 86175
rect 95099 86147 95134 86175
rect 94974 86113 95134 86147
rect 94974 86085 95009 86113
rect 95037 86085 95071 86113
rect 95099 86085 95134 86113
rect 94974 86051 95134 86085
rect 94974 86023 95009 86051
rect 95037 86023 95071 86051
rect 95099 86023 95134 86051
rect 94974 85989 95134 86023
rect 94974 85961 95009 85989
rect 95037 85961 95071 85989
rect 95099 85961 95134 85989
rect 94974 85944 95134 85961
rect 99474 86175 99634 86192
rect 99474 86147 99509 86175
rect 99537 86147 99571 86175
rect 99599 86147 99634 86175
rect 99474 86113 99634 86147
rect 99474 86085 99509 86113
rect 99537 86085 99571 86113
rect 99599 86085 99634 86113
rect 99474 86051 99634 86085
rect 99474 86023 99509 86051
rect 99537 86023 99571 86051
rect 99599 86023 99634 86051
rect 99474 85989 99634 86023
rect 99474 85961 99509 85989
rect 99537 85961 99571 85989
rect 99599 85961 99634 85989
rect 99474 85944 99634 85961
rect 103974 86175 104134 86192
rect 103974 86147 104009 86175
rect 104037 86147 104071 86175
rect 104099 86147 104134 86175
rect 103974 86113 104134 86147
rect 103974 86085 104009 86113
rect 104037 86085 104071 86113
rect 104099 86085 104134 86113
rect 103974 86051 104134 86085
rect 103974 86023 104009 86051
rect 104037 86023 104071 86051
rect 104099 86023 104134 86051
rect 103974 85989 104134 86023
rect 103974 85961 104009 85989
rect 104037 85961 104071 85989
rect 104099 85961 104134 85989
rect 103974 85944 104134 85961
rect 108474 86175 108634 86192
rect 108474 86147 108509 86175
rect 108537 86147 108571 86175
rect 108599 86147 108634 86175
rect 108474 86113 108634 86147
rect 108474 86085 108509 86113
rect 108537 86085 108571 86113
rect 108599 86085 108634 86113
rect 108474 86051 108634 86085
rect 108474 86023 108509 86051
rect 108537 86023 108571 86051
rect 108599 86023 108634 86051
rect 108474 85989 108634 86023
rect 108474 85961 108509 85989
rect 108537 85961 108571 85989
rect 108599 85961 108634 85989
rect 108474 85944 108634 85961
rect 112974 86175 113134 86192
rect 112974 86147 113009 86175
rect 113037 86147 113071 86175
rect 113099 86147 113134 86175
rect 112974 86113 113134 86147
rect 112974 86085 113009 86113
rect 113037 86085 113071 86113
rect 113099 86085 113134 86113
rect 112974 86051 113134 86085
rect 112974 86023 113009 86051
rect 113037 86023 113071 86051
rect 113099 86023 113134 86051
rect 112974 85989 113134 86023
rect 112974 85961 113009 85989
rect 113037 85961 113071 85989
rect 113099 85961 113134 85989
rect 112974 85944 113134 85961
rect 117474 86175 117634 86192
rect 117474 86147 117509 86175
rect 117537 86147 117571 86175
rect 117599 86147 117634 86175
rect 117474 86113 117634 86147
rect 117474 86085 117509 86113
rect 117537 86085 117571 86113
rect 117599 86085 117634 86113
rect 117474 86051 117634 86085
rect 117474 86023 117509 86051
rect 117537 86023 117571 86051
rect 117599 86023 117634 86051
rect 117474 85989 117634 86023
rect 117474 85961 117509 85989
rect 117537 85961 117571 85989
rect 117599 85961 117634 85989
rect 117474 85944 117634 85961
rect 120437 86175 120747 94961
rect 120437 86147 120485 86175
rect 120513 86147 120547 86175
rect 120575 86147 120609 86175
rect 120637 86147 120671 86175
rect 120699 86147 120747 86175
rect 120437 86113 120747 86147
rect 120437 86085 120485 86113
rect 120513 86085 120547 86113
rect 120575 86085 120609 86113
rect 120637 86085 120671 86113
rect 120699 86085 120747 86113
rect 120437 86051 120747 86085
rect 120437 86023 120485 86051
rect 120513 86023 120547 86051
rect 120575 86023 120609 86051
rect 120637 86023 120671 86051
rect 120699 86023 120747 86051
rect 120437 85989 120747 86023
rect 120437 85961 120485 85989
rect 120513 85961 120547 85989
rect 120575 85961 120609 85989
rect 120637 85961 120671 85989
rect 120699 85961 120747 85989
rect 91577 83147 91625 83175
rect 91653 83147 91687 83175
rect 91715 83147 91749 83175
rect 91777 83147 91811 83175
rect 91839 83147 91887 83175
rect 91577 83113 91887 83147
rect 91577 83085 91625 83113
rect 91653 83085 91687 83113
rect 91715 83085 91749 83113
rect 91777 83085 91811 83113
rect 91839 83085 91887 83113
rect 91577 83051 91887 83085
rect 91577 83023 91625 83051
rect 91653 83023 91687 83051
rect 91715 83023 91749 83051
rect 91777 83023 91811 83051
rect 91839 83023 91887 83051
rect 91577 82989 91887 83023
rect 91577 82961 91625 82989
rect 91653 82961 91687 82989
rect 91715 82961 91749 82989
rect 91777 82961 91811 82989
rect 91839 82961 91887 82989
rect 84437 77147 84485 77175
rect 84513 77147 84547 77175
rect 84575 77147 84609 77175
rect 84637 77147 84671 77175
rect 84699 77147 84747 77175
rect 84437 77113 84747 77147
rect 84437 77085 84485 77113
rect 84513 77085 84547 77113
rect 84575 77085 84609 77113
rect 84637 77085 84671 77113
rect 84699 77085 84747 77113
rect 84437 77051 84747 77085
rect 84437 77023 84485 77051
rect 84513 77023 84547 77051
rect 84575 77023 84609 77051
rect 84637 77023 84671 77051
rect 84699 77023 84747 77051
rect 84437 76989 84747 77023
rect 84437 76961 84485 76989
rect 84513 76961 84547 76989
rect 84575 76961 84609 76989
rect 84637 76961 84671 76989
rect 84699 76961 84747 76989
rect 82577 74147 82625 74175
rect 82653 74147 82687 74175
rect 82715 74147 82749 74175
rect 82777 74147 82811 74175
rect 82839 74147 82887 74175
rect 82577 74113 82887 74147
rect 82577 74085 82625 74113
rect 82653 74085 82687 74113
rect 82715 74085 82749 74113
rect 82777 74085 82811 74113
rect 82839 74085 82887 74113
rect 82577 74051 82887 74085
rect 82577 74023 82625 74051
rect 82653 74023 82687 74051
rect 82715 74023 82749 74051
rect 82777 74023 82811 74051
rect 82839 74023 82887 74051
rect 82577 73989 82887 74023
rect 82577 73961 82625 73989
rect 82653 73961 82687 73989
rect 82715 73961 82749 73989
rect 82777 73961 82811 73989
rect 82839 73961 82887 73989
rect 75437 68147 75485 68175
rect 75513 68147 75547 68175
rect 75575 68147 75609 68175
rect 75637 68147 75671 68175
rect 75699 68147 75747 68175
rect 75437 68113 75747 68147
rect 75437 68085 75485 68113
rect 75513 68085 75547 68113
rect 75575 68085 75609 68113
rect 75637 68085 75671 68113
rect 75699 68085 75747 68113
rect 75437 68051 75747 68085
rect 75437 68023 75485 68051
rect 75513 68023 75547 68051
rect 75575 68023 75609 68051
rect 75637 68023 75671 68051
rect 75699 68023 75747 68051
rect 75437 67989 75747 68023
rect 75437 67961 75485 67989
rect 75513 67961 75547 67989
rect 75575 67961 75609 67989
rect 75637 67961 75671 67989
rect 75699 67961 75747 67989
rect 73577 65147 73625 65175
rect 73653 65147 73687 65175
rect 73715 65147 73749 65175
rect 73777 65147 73811 65175
rect 73839 65147 73887 65175
rect 73577 65113 73887 65147
rect 73577 65085 73625 65113
rect 73653 65085 73687 65113
rect 73715 65085 73749 65113
rect 73777 65085 73811 65113
rect 73839 65085 73887 65113
rect 73577 65051 73887 65085
rect 73577 65023 73625 65051
rect 73653 65023 73687 65051
rect 73715 65023 73749 65051
rect 73777 65023 73811 65051
rect 73839 65023 73887 65051
rect 73577 64989 73887 65023
rect 73577 64961 73625 64989
rect 73653 64961 73687 64989
rect 73715 64961 73749 64989
rect 73777 64961 73811 64989
rect 73839 64961 73887 64989
rect 66437 59147 66485 59175
rect 66513 59147 66547 59175
rect 66575 59147 66609 59175
rect 66637 59147 66671 59175
rect 66699 59147 66747 59175
rect 66437 59113 66747 59147
rect 66437 59085 66485 59113
rect 66513 59085 66547 59113
rect 66575 59085 66609 59113
rect 66637 59085 66671 59113
rect 66699 59085 66747 59113
rect 66437 59051 66747 59085
rect 66437 59023 66485 59051
rect 66513 59023 66547 59051
rect 66575 59023 66609 59051
rect 66637 59023 66671 59051
rect 66699 59023 66747 59051
rect 66437 58989 66747 59023
rect 66437 58961 66485 58989
rect 66513 58961 66547 58989
rect 66575 58961 66609 58989
rect 66637 58961 66671 58989
rect 66699 58961 66747 58989
rect 64577 56147 64625 56175
rect 64653 56147 64687 56175
rect 64715 56147 64749 56175
rect 64777 56147 64811 56175
rect 64839 56147 64887 56175
rect 64577 56113 64887 56147
rect 64577 56085 64625 56113
rect 64653 56085 64687 56113
rect 64715 56085 64749 56113
rect 64777 56085 64811 56113
rect 64839 56085 64887 56113
rect 64577 56051 64887 56085
rect 64577 56023 64625 56051
rect 64653 56023 64687 56051
rect 64715 56023 64749 56051
rect 64777 56023 64811 56051
rect 64839 56023 64887 56051
rect 64577 55989 64887 56023
rect 64577 55961 64625 55989
rect 64653 55961 64687 55989
rect 64715 55961 64749 55989
rect 64777 55961 64811 55989
rect 64839 55961 64887 55989
rect 57437 50147 57485 50175
rect 57513 50147 57547 50175
rect 57575 50147 57609 50175
rect 57637 50147 57671 50175
rect 57699 50147 57747 50175
rect 57437 50113 57747 50147
rect 57437 50085 57485 50113
rect 57513 50085 57547 50113
rect 57575 50085 57609 50113
rect 57637 50085 57671 50113
rect 57699 50085 57747 50113
rect 57437 50051 57747 50085
rect 57437 50023 57485 50051
rect 57513 50023 57547 50051
rect 57575 50023 57609 50051
rect 57637 50023 57671 50051
rect 57699 50023 57747 50051
rect 57437 49989 57747 50023
rect 57437 49961 57485 49989
rect 57513 49961 57547 49989
rect 57575 49961 57609 49989
rect 57637 49961 57671 49989
rect 57699 49961 57747 49989
rect 57437 41175 57747 49961
rect 57437 41147 57485 41175
rect 57513 41147 57547 41175
rect 57575 41147 57609 41175
rect 57637 41147 57671 41175
rect 57699 41147 57747 41175
rect 57437 41113 57747 41147
rect 57437 41085 57485 41113
rect 57513 41085 57547 41113
rect 57575 41085 57609 41113
rect 57637 41085 57671 41113
rect 57699 41085 57747 41113
rect 57437 41051 57747 41085
rect 57437 41023 57485 41051
rect 57513 41023 57547 41051
rect 57575 41023 57609 41051
rect 57637 41023 57671 41051
rect 57699 41023 57747 41051
rect 57437 40989 57747 41023
rect 57437 40961 57485 40989
rect 57513 40961 57547 40989
rect 57575 40961 57609 40989
rect 57637 40961 57671 40989
rect 57699 40961 57747 40989
rect 57437 32175 57747 40961
rect 57437 32147 57485 32175
rect 57513 32147 57547 32175
rect 57575 32147 57609 32175
rect 57637 32147 57671 32175
rect 57699 32147 57747 32175
rect 57437 32113 57747 32147
rect 57437 32085 57485 32113
rect 57513 32085 57547 32113
rect 57575 32085 57609 32113
rect 57637 32085 57671 32113
rect 57699 32085 57747 32113
rect 57437 32051 57747 32085
rect 57437 32023 57485 32051
rect 57513 32023 57547 32051
rect 57575 32023 57609 32051
rect 57637 32023 57671 32051
rect 57699 32023 57747 32051
rect 57437 31989 57747 32023
rect 57437 31961 57485 31989
rect 57513 31961 57547 31989
rect 57575 31961 57609 31989
rect 57637 31961 57671 31989
rect 57699 31961 57747 31989
rect 57437 23175 57747 31961
rect 57437 23147 57485 23175
rect 57513 23147 57547 23175
rect 57575 23147 57609 23175
rect 57637 23147 57671 23175
rect 57699 23147 57747 23175
rect 57437 23113 57747 23147
rect 57437 23085 57485 23113
rect 57513 23085 57547 23113
rect 57575 23085 57609 23113
rect 57637 23085 57671 23113
rect 57699 23085 57747 23113
rect 57437 23051 57747 23085
rect 57437 23023 57485 23051
rect 57513 23023 57547 23051
rect 57575 23023 57609 23051
rect 57637 23023 57671 23051
rect 57699 23023 57747 23051
rect 57437 22989 57747 23023
rect 57437 22961 57485 22989
rect 57513 22961 57547 22989
rect 57575 22961 57609 22989
rect 57637 22961 57671 22989
rect 57699 22961 57747 22989
rect 57437 14175 57747 22961
rect 57437 14147 57485 14175
rect 57513 14147 57547 14175
rect 57575 14147 57609 14175
rect 57637 14147 57671 14175
rect 57699 14147 57747 14175
rect 57437 14113 57747 14147
rect 57437 14085 57485 14113
rect 57513 14085 57547 14113
rect 57575 14085 57609 14113
rect 57637 14085 57671 14113
rect 57699 14085 57747 14113
rect 57437 14051 57747 14085
rect 57437 14023 57485 14051
rect 57513 14023 57547 14051
rect 57575 14023 57609 14051
rect 57637 14023 57671 14051
rect 57699 14023 57747 14051
rect 57437 13989 57747 14023
rect 57437 13961 57485 13989
rect 57513 13961 57547 13989
rect 57575 13961 57609 13989
rect 57637 13961 57671 13989
rect 57699 13961 57747 13989
rect 57437 5175 57747 13961
rect 57437 5147 57485 5175
rect 57513 5147 57547 5175
rect 57575 5147 57609 5175
rect 57637 5147 57671 5175
rect 57699 5147 57747 5175
rect 57437 5113 57747 5147
rect 57437 5085 57485 5113
rect 57513 5085 57547 5113
rect 57575 5085 57609 5113
rect 57637 5085 57671 5113
rect 57699 5085 57747 5113
rect 57437 5051 57747 5085
rect 57437 5023 57485 5051
rect 57513 5023 57547 5051
rect 57575 5023 57609 5051
rect 57637 5023 57671 5051
rect 57699 5023 57747 5051
rect 57437 4989 57747 5023
rect 57437 4961 57485 4989
rect 57513 4961 57547 4989
rect 57575 4961 57609 4989
rect 57637 4961 57671 4989
rect 57699 4961 57747 4989
rect 57437 -560 57747 4961
rect 57437 -588 57485 -560
rect 57513 -588 57547 -560
rect 57575 -588 57609 -560
rect 57637 -588 57671 -560
rect 57699 -588 57747 -560
rect 57437 -622 57747 -588
rect 57437 -650 57485 -622
rect 57513 -650 57547 -622
rect 57575 -650 57609 -622
rect 57637 -650 57671 -622
rect 57699 -650 57747 -622
rect 57437 -684 57747 -650
rect 57437 -712 57485 -684
rect 57513 -712 57547 -684
rect 57575 -712 57609 -684
rect 57637 -712 57671 -684
rect 57699 -712 57747 -684
rect 57437 -746 57747 -712
rect 57437 -774 57485 -746
rect 57513 -774 57547 -746
rect 57575 -774 57609 -746
rect 57637 -774 57671 -746
rect 57699 -774 57747 -746
rect 57437 -822 57747 -774
rect 64577 47175 64887 55961
rect 65724 56175 65884 56192
rect 65724 56147 65759 56175
rect 65787 56147 65821 56175
rect 65849 56147 65884 56175
rect 65724 56113 65884 56147
rect 65724 56085 65759 56113
rect 65787 56085 65821 56113
rect 65849 56085 65884 56113
rect 65724 56051 65884 56085
rect 65724 56023 65759 56051
rect 65787 56023 65821 56051
rect 65849 56023 65884 56051
rect 65724 55989 65884 56023
rect 65724 55961 65759 55989
rect 65787 55961 65821 55989
rect 65849 55961 65884 55989
rect 65724 55944 65884 55961
rect 64577 47147 64625 47175
rect 64653 47147 64687 47175
rect 64715 47147 64749 47175
rect 64777 47147 64811 47175
rect 64839 47147 64887 47175
rect 64577 47113 64887 47147
rect 64577 47085 64625 47113
rect 64653 47085 64687 47113
rect 64715 47085 64749 47113
rect 64777 47085 64811 47113
rect 64839 47085 64887 47113
rect 64577 47051 64887 47085
rect 64577 47023 64625 47051
rect 64653 47023 64687 47051
rect 64715 47023 64749 47051
rect 64777 47023 64811 47051
rect 64839 47023 64887 47051
rect 64577 46989 64887 47023
rect 64577 46961 64625 46989
rect 64653 46961 64687 46989
rect 64715 46961 64749 46989
rect 64777 46961 64811 46989
rect 64839 46961 64887 46989
rect 64577 38175 64887 46961
rect 64577 38147 64625 38175
rect 64653 38147 64687 38175
rect 64715 38147 64749 38175
rect 64777 38147 64811 38175
rect 64839 38147 64887 38175
rect 64577 38113 64887 38147
rect 64577 38085 64625 38113
rect 64653 38085 64687 38113
rect 64715 38085 64749 38113
rect 64777 38085 64811 38113
rect 64839 38085 64887 38113
rect 64577 38051 64887 38085
rect 64577 38023 64625 38051
rect 64653 38023 64687 38051
rect 64715 38023 64749 38051
rect 64777 38023 64811 38051
rect 64839 38023 64887 38051
rect 64577 37989 64887 38023
rect 64577 37961 64625 37989
rect 64653 37961 64687 37989
rect 64715 37961 64749 37989
rect 64777 37961 64811 37989
rect 64839 37961 64887 37989
rect 64577 29175 64887 37961
rect 64577 29147 64625 29175
rect 64653 29147 64687 29175
rect 64715 29147 64749 29175
rect 64777 29147 64811 29175
rect 64839 29147 64887 29175
rect 64577 29113 64887 29147
rect 64577 29085 64625 29113
rect 64653 29085 64687 29113
rect 64715 29085 64749 29113
rect 64777 29085 64811 29113
rect 64839 29085 64887 29113
rect 64577 29051 64887 29085
rect 64577 29023 64625 29051
rect 64653 29023 64687 29051
rect 64715 29023 64749 29051
rect 64777 29023 64811 29051
rect 64839 29023 64887 29051
rect 64577 28989 64887 29023
rect 64577 28961 64625 28989
rect 64653 28961 64687 28989
rect 64715 28961 64749 28989
rect 64777 28961 64811 28989
rect 64839 28961 64887 28989
rect 64577 20175 64887 28961
rect 64577 20147 64625 20175
rect 64653 20147 64687 20175
rect 64715 20147 64749 20175
rect 64777 20147 64811 20175
rect 64839 20147 64887 20175
rect 64577 20113 64887 20147
rect 64577 20085 64625 20113
rect 64653 20085 64687 20113
rect 64715 20085 64749 20113
rect 64777 20085 64811 20113
rect 64839 20085 64887 20113
rect 64577 20051 64887 20085
rect 64577 20023 64625 20051
rect 64653 20023 64687 20051
rect 64715 20023 64749 20051
rect 64777 20023 64811 20051
rect 64839 20023 64887 20051
rect 64577 19989 64887 20023
rect 64577 19961 64625 19989
rect 64653 19961 64687 19989
rect 64715 19961 64749 19989
rect 64777 19961 64811 19989
rect 64839 19961 64887 19989
rect 64577 11175 64887 19961
rect 64577 11147 64625 11175
rect 64653 11147 64687 11175
rect 64715 11147 64749 11175
rect 64777 11147 64811 11175
rect 64839 11147 64887 11175
rect 64577 11113 64887 11147
rect 64577 11085 64625 11113
rect 64653 11085 64687 11113
rect 64715 11085 64749 11113
rect 64777 11085 64811 11113
rect 64839 11085 64887 11113
rect 64577 11051 64887 11085
rect 64577 11023 64625 11051
rect 64653 11023 64687 11051
rect 64715 11023 64749 11051
rect 64777 11023 64811 11051
rect 64839 11023 64887 11051
rect 64577 10989 64887 11023
rect 64577 10961 64625 10989
rect 64653 10961 64687 10989
rect 64715 10961 64749 10989
rect 64777 10961 64811 10989
rect 64839 10961 64887 10989
rect 64577 2175 64887 10961
rect 64577 2147 64625 2175
rect 64653 2147 64687 2175
rect 64715 2147 64749 2175
rect 64777 2147 64811 2175
rect 64839 2147 64887 2175
rect 64577 2113 64887 2147
rect 64577 2085 64625 2113
rect 64653 2085 64687 2113
rect 64715 2085 64749 2113
rect 64777 2085 64811 2113
rect 64839 2085 64887 2113
rect 64577 2051 64887 2085
rect 64577 2023 64625 2051
rect 64653 2023 64687 2051
rect 64715 2023 64749 2051
rect 64777 2023 64811 2051
rect 64839 2023 64887 2051
rect 64577 1989 64887 2023
rect 64577 1961 64625 1989
rect 64653 1961 64687 1989
rect 64715 1961 64749 1989
rect 64777 1961 64811 1989
rect 64839 1961 64887 1989
rect 64577 -80 64887 1961
rect 64577 -108 64625 -80
rect 64653 -108 64687 -80
rect 64715 -108 64749 -80
rect 64777 -108 64811 -80
rect 64839 -108 64887 -80
rect 64577 -142 64887 -108
rect 64577 -170 64625 -142
rect 64653 -170 64687 -142
rect 64715 -170 64749 -142
rect 64777 -170 64811 -142
rect 64839 -170 64887 -142
rect 64577 -204 64887 -170
rect 64577 -232 64625 -204
rect 64653 -232 64687 -204
rect 64715 -232 64749 -204
rect 64777 -232 64811 -204
rect 64839 -232 64887 -204
rect 64577 -266 64887 -232
rect 64577 -294 64625 -266
rect 64653 -294 64687 -266
rect 64715 -294 64749 -266
rect 64777 -294 64811 -266
rect 64839 -294 64887 -266
rect 64577 -822 64887 -294
rect 66437 50175 66747 58961
rect 67974 59175 68134 59192
rect 67974 59147 68009 59175
rect 68037 59147 68071 59175
rect 68099 59147 68134 59175
rect 67974 59113 68134 59147
rect 67974 59085 68009 59113
rect 68037 59085 68071 59113
rect 68099 59085 68134 59113
rect 67974 59051 68134 59085
rect 67974 59023 68009 59051
rect 68037 59023 68071 59051
rect 68099 59023 68134 59051
rect 67974 58989 68134 59023
rect 67974 58961 68009 58989
rect 68037 58961 68071 58989
rect 68099 58961 68134 58989
rect 67974 58944 68134 58961
rect 72474 59175 72634 59192
rect 72474 59147 72509 59175
rect 72537 59147 72571 59175
rect 72599 59147 72634 59175
rect 72474 59113 72634 59147
rect 72474 59085 72509 59113
rect 72537 59085 72571 59113
rect 72599 59085 72634 59113
rect 72474 59051 72634 59085
rect 72474 59023 72509 59051
rect 72537 59023 72571 59051
rect 72599 59023 72634 59051
rect 72474 58989 72634 59023
rect 72474 58961 72509 58989
rect 72537 58961 72571 58989
rect 72599 58961 72634 58989
rect 72474 58944 72634 58961
rect 70224 56175 70384 56192
rect 70224 56147 70259 56175
rect 70287 56147 70321 56175
rect 70349 56147 70384 56175
rect 70224 56113 70384 56147
rect 70224 56085 70259 56113
rect 70287 56085 70321 56113
rect 70349 56085 70384 56113
rect 70224 56051 70384 56085
rect 70224 56023 70259 56051
rect 70287 56023 70321 56051
rect 70349 56023 70384 56051
rect 70224 55989 70384 56023
rect 70224 55961 70259 55989
rect 70287 55961 70321 55989
rect 70349 55961 70384 55989
rect 70224 55944 70384 55961
rect 73577 56175 73887 64961
rect 74724 65175 74884 65192
rect 74724 65147 74759 65175
rect 74787 65147 74821 65175
rect 74849 65147 74884 65175
rect 74724 65113 74884 65147
rect 74724 65085 74759 65113
rect 74787 65085 74821 65113
rect 74849 65085 74884 65113
rect 74724 65051 74884 65085
rect 74724 65023 74759 65051
rect 74787 65023 74821 65051
rect 74849 65023 74884 65051
rect 74724 64989 74884 65023
rect 74724 64961 74759 64989
rect 74787 64961 74821 64989
rect 74849 64961 74884 64989
rect 74724 64944 74884 64961
rect 75437 59175 75747 67961
rect 76974 68175 77134 68192
rect 76974 68147 77009 68175
rect 77037 68147 77071 68175
rect 77099 68147 77134 68175
rect 76974 68113 77134 68147
rect 76974 68085 77009 68113
rect 77037 68085 77071 68113
rect 77099 68085 77134 68113
rect 76974 68051 77134 68085
rect 76974 68023 77009 68051
rect 77037 68023 77071 68051
rect 77099 68023 77134 68051
rect 76974 67989 77134 68023
rect 76974 67961 77009 67989
rect 77037 67961 77071 67989
rect 77099 67961 77134 67989
rect 76974 67944 77134 67961
rect 81474 68175 81634 68192
rect 81474 68147 81509 68175
rect 81537 68147 81571 68175
rect 81599 68147 81634 68175
rect 81474 68113 81634 68147
rect 81474 68085 81509 68113
rect 81537 68085 81571 68113
rect 81599 68085 81634 68113
rect 81474 68051 81634 68085
rect 81474 68023 81509 68051
rect 81537 68023 81571 68051
rect 81599 68023 81634 68051
rect 81474 67989 81634 68023
rect 81474 67961 81509 67989
rect 81537 67961 81571 67989
rect 81599 67961 81634 67989
rect 81474 67944 81634 67961
rect 79224 65175 79384 65192
rect 79224 65147 79259 65175
rect 79287 65147 79321 65175
rect 79349 65147 79384 65175
rect 79224 65113 79384 65147
rect 79224 65085 79259 65113
rect 79287 65085 79321 65113
rect 79349 65085 79384 65113
rect 79224 65051 79384 65085
rect 79224 65023 79259 65051
rect 79287 65023 79321 65051
rect 79349 65023 79384 65051
rect 79224 64989 79384 65023
rect 79224 64961 79259 64989
rect 79287 64961 79321 64989
rect 79349 64961 79384 64989
rect 79224 64944 79384 64961
rect 82577 65175 82887 73961
rect 83724 74175 83884 74192
rect 83724 74147 83759 74175
rect 83787 74147 83821 74175
rect 83849 74147 83884 74175
rect 83724 74113 83884 74147
rect 83724 74085 83759 74113
rect 83787 74085 83821 74113
rect 83849 74085 83884 74113
rect 83724 74051 83884 74085
rect 83724 74023 83759 74051
rect 83787 74023 83821 74051
rect 83849 74023 83884 74051
rect 83724 73989 83884 74023
rect 83724 73961 83759 73989
rect 83787 73961 83821 73989
rect 83849 73961 83884 73989
rect 83724 73944 83884 73961
rect 84437 68175 84747 76961
rect 85974 77175 86134 77192
rect 85974 77147 86009 77175
rect 86037 77147 86071 77175
rect 86099 77147 86134 77175
rect 85974 77113 86134 77147
rect 85974 77085 86009 77113
rect 86037 77085 86071 77113
rect 86099 77085 86134 77113
rect 85974 77051 86134 77085
rect 85974 77023 86009 77051
rect 86037 77023 86071 77051
rect 86099 77023 86134 77051
rect 85974 76989 86134 77023
rect 85974 76961 86009 76989
rect 86037 76961 86071 76989
rect 86099 76961 86134 76989
rect 85974 76944 86134 76961
rect 90474 77175 90634 77192
rect 90474 77147 90509 77175
rect 90537 77147 90571 77175
rect 90599 77147 90634 77175
rect 90474 77113 90634 77147
rect 90474 77085 90509 77113
rect 90537 77085 90571 77113
rect 90599 77085 90634 77113
rect 90474 77051 90634 77085
rect 90474 77023 90509 77051
rect 90537 77023 90571 77051
rect 90599 77023 90634 77051
rect 90474 76989 90634 77023
rect 90474 76961 90509 76989
rect 90537 76961 90571 76989
rect 90599 76961 90634 76989
rect 90474 76944 90634 76961
rect 88224 74175 88384 74192
rect 88224 74147 88259 74175
rect 88287 74147 88321 74175
rect 88349 74147 88384 74175
rect 88224 74113 88384 74147
rect 88224 74085 88259 74113
rect 88287 74085 88321 74113
rect 88349 74085 88384 74113
rect 88224 74051 88384 74085
rect 88224 74023 88259 74051
rect 88287 74023 88321 74051
rect 88349 74023 88384 74051
rect 88224 73989 88384 74023
rect 88224 73961 88259 73989
rect 88287 73961 88321 73989
rect 88349 73961 88384 73989
rect 88224 73944 88384 73961
rect 91577 74175 91887 82961
rect 92724 83175 92884 83192
rect 92724 83147 92759 83175
rect 92787 83147 92821 83175
rect 92849 83147 92884 83175
rect 92724 83113 92884 83147
rect 92724 83085 92759 83113
rect 92787 83085 92821 83113
rect 92849 83085 92884 83113
rect 92724 83051 92884 83085
rect 92724 83023 92759 83051
rect 92787 83023 92821 83051
rect 92849 83023 92884 83051
rect 92724 82989 92884 83023
rect 92724 82961 92759 82989
rect 92787 82961 92821 82989
rect 92849 82961 92884 82989
rect 92724 82944 92884 82961
rect 97224 83175 97384 83192
rect 97224 83147 97259 83175
rect 97287 83147 97321 83175
rect 97349 83147 97384 83175
rect 97224 83113 97384 83147
rect 97224 83085 97259 83113
rect 97287 83085 97321 83113
rect 97349 83085 97384 83113
rect 97224 83051 97384 83085
rect 97224 83023 97259 83051
rect 97287 83023 97321 83051
rect 97349 83023 97384 83051
rect 97224 82989 97384 83023
rect 97224 82961 97259 82989
rect 97287 82961 97321 82989
rect 97349 82961 97384 82989
rect 97224 82944 97384 82961
rect 101724 83175 101884 83192
rect 101724 83147 101759 83175
rect 101787 83147 101821 83175
rect 101849 83147 101884 83175
rect 101724 83113 101884 83147
rect 101724 83085 101759 83113
rect 101787 83085 101821 83113
rect 101849 83085 101884 83113
rect 101724 83051 101884 83085
rect 101724 83023 101759 83051
rect 101787 83023 101821 83051
rect 101849 83023 101884 83051
rect 101724 82989 101884 83023
rect 101724 82961 101759 82989
rect 101787 82961 101821 82989
rect 101849 82961 101884 82989
rect 101724 82944 101884 82961
rect 106224 83175 106384 83192
rect 106224 83147 106259 83175
rect 106287 83147 106321 83175
rect 106349 83147 106384 83175
rect 106224 83113 106384 83147
rect 106224 83085 106259 83113
rect 106287 83085 106321 83113
rect 106349 83085 106384 83113
rect 106224 83051 106384 83085
rect 106224 83023 106259 83051
rect 106287 83023 106321 83051
rect 106349 83023 106384 83051
rect 106224 82989 106384 83023
rect 106224 82961 106259 82989
rect 106287 82961 106321 82989
rect 106349 82961 106384 82989
rect 106224 82944 106384 82961
rect 110724 83175 110884 83192
rect 110724 83147 110759 83175
rect 110787 83147 110821 83175
rect 110849 83147 110884 83175
rect 110724 83113 110884 83147
rect 110724 83085 110759 83113
rect 110787 83085 110821 83113
rect 110849 83085 110884 83113
rect 110724 83051 110884 83085
rect 110724 83023 110759 83051
rect 110787 83023 110821 83051
rect 110849 83023 110884 83051
rect 110724 82989 110884 83023
rect 110724 82961 110759 82989
rect 110787 82961 110821 82989
rect 110849 82961 110884 82989
rect 110724 82944 110884 82961
rect 115224 83175 115384 83192
rect 115224 83147 115259 83175
rect 115287 83147 115321 83175
rect 115349 83147 115384 83175
rect 115224 83113 115384 83147
rect 115224 83085 115259 83113
rect 115287 83085 115321 83113
rect 115349 83085 115384 83113
rect 115224 83051 115384 83085
rect 115224 83023 115259 83051
rect 115287 83023 115321 83051
rect 115349 83023 115384 83051
rect 115224 82989 115384 83023
rect 115224 82961 115259 82989
rect 115287 82961 115321 82989
rect 115349 82961 115384 82989
rect 115224 82944 115384 82961
rect 94974 77175 95134 77192
rect 94974 77147 95009 77175
rect 95037 77147 95071 77175
rect 95099 77147 95134 77175
rect 94974 77113 95134 77147
rect 94974 77085 95009 77113
rect 95037 77085 95071 77113
rect 95099 77085 95134 77113
rect 94974 77051 95134 77085
rect 94974 77023 95009 77051
rect 95037 77023 95071 77051
rect 95099 77023 95134 77051
rect 94974 76989 95134 77023
rect 94974 76961 95009 76989
rect 95037 76961 95071 76989
rect 95099 76961 95134 76989
rect 94974 76944 95134 76961
rect 99474 77175 99634 77192
rect 99474 77147 99509 77175
rect 99537 77147 99571 77175
rect 99599 77147 99634 77175
rect 99474 77113 99634 77147
rect 99474 77085 99509 77113
rect 99537 77085 99571 77113
rect 99599 77085 99634 77113
rect 99474 77051 99634 77085
rect 99474 77023 99509 77051
rect 99537 77023 99571 77051
rect 99599 77023 99634 77051
rect 99474 76989 99634 77023
rect 99474 76961 99509 76989
rect 99537 76961 99571 76989
rect 99599 76961 99634 76989
rect 99474 76944 99634 76961
rect 103974 77175 104134 77192
rect 103974 77147 104009 77175
rect 104037 77147 104071 77175
rect 104099 77147 104134 77175
rect 103974 77113 104134 77147
rect 103974 77085 104009 77113
rect 104037 77085 104071 77113
rect 104099 77085 104134 77113
rect 103974 77051 104134 77085
rect 103974 77023 104009 77051
rect 104037 77023 104071 77051
rect 104099 77023 104134 77051
rect 103974 76989 104134 77023
rect 103974 76961 104009 76989
rect 104037 76961 104071 76989
rect 104099 76961 104134 76989
rect 103974 76944 104134 76961
rect 108474 77175 108634 77192
rect 108474 77147 108509 77175
rect 108537 77147 108571 77175
rect 108599 77147 108634 77175
rect 108474 77113 108634 77147
rect 108474 77085 108509 77113
rect 108537 77085 108571 77113
rect 108599 77085 108634 77113
rect 108474 77051 108634 77085
rect 108474 77023 108509 77051
rect 108537 77023 108571 77051
rect 108599 77023 108634 77051
rect 108474 76989 108634 77023
rect 108474 76961 108509 76989
rect 108537 76961 108571 76989
rect 108599 76961 108634 76989
rect 108474 76944 108634 76961
rect 112974 77175 113134 77192
rect 112974 77147 113009 77175
rect 113037 77147 113071 77175
rect 113099 77147 113134 77175
rect 112974 77113 113134 77147
rect 112974 77085 113009 77113
rect 113037 77085 113071 77113
rect 113099 77085 113134 77113
rect 112974 77051 113134 77085
rect 112974 77023 113009 77051
rect 113037 77023 113071 77051
rect 113099 77023 113134 77051
rect 112974 76989 113134 77023
rect 112974 76961 113009 76989
rect 113037 76961 113071 76989
rect 113099 76961 113134 76989
rect 112974 76944 113134 76961
rect 117474 77175 117634 77192
rect 117474 77147 117509 77175
rect 117537 77147 117571 77175
rect 117599 77147 117634 77175
rect 117474 77113 117634 77147
rect 117474 77085 117509 77113
rect 117537 77085 117571 77113
rect 117599 77085 117634 77113
rect 117474 77051 117634 77085
rect 117474 77023 117509 77051
rect 117537 77023 117571 77051
rect 117599 77023 117634 77051
rect 117474 76989 117634 77023
rect 117474 76961 117509 76989
rect 117537 76961 117571 76989
rect 117599 76961 117634 76989
rect 117474 76944 117634 76961
rect 120437 77175 120747 85961
rect 120437 77147 120485 77175
rect 120513 77147 120547 77175
rect 120575 77147 120609 77175
rect 120637 77147 120671 77175
rect 120699 77147 120747 77175
rect 120437 77113 120747 77147
rect 120437 77085 120485 77113
rect 120513 77085 120547 77113
rect 120575 77085 120609 77113
rect 120637 77085 120671 77113
rect 120699 77085 120747 77113
rect 120437 77051 120747 77085
rect 120437 77023 120485 77051
rect 120513 77023 120547 77051
rect 120575 77023 120609 77051
rect 120637 77023 120671 77051
rect 120699 77023 120747 77051
rect 120437 76989 120747 77023
rect 120437 76961 120485 76989
rect 120513 76961 120547 76989
rect 120575 76961 120609 76989
rect 120637 76961 120671 76989
rect 120699 76961 120747 76989
rect 91577 74147 91625 74175
rect 91653 74147 91687 74175
rect 91715 74147 91749 74175
rect 91777 74147 91811 74175
rect 91839 74147 91887 74175
rect 91577 74113 91887 74147
rect 91577 74085 91625 74113
rect 91653 74085 91687 74113
rect 91715 74085 91749 74113
rect 91777 74085 91811 74113
rect 91839 74085 91887 74113
rect 91577 74051 91887 74085
rect 91577 74023 91625 74051
rect 91653 74023 91687 74051
rect 91715 74023 91749 74051
rect 91777 74023 91811 74051
rect 91839 74023 91887 74051
rect 91577 73989 91887 74023
rect 91577 73961 91625 73989
rect 91653 73961 91687 73989
rect 91715 73961 91749 73989
rect 91777 73961 91811 73989
rect 91839 73961 91887 73989
rect 84437 68147 84485 68175
rect 84513 68147 84547 68175
rect 84575 68147 84609 68175
rect 84637 68147 84671 68175
rect 84699 68147 84747 68175
rect 84437 68113 84747 68147
rect 84437 68085 84485 68113
rect 84513 68085 84547 68113
rect 84575 68085 84609 68113
rect 84637 68085 84671 68113
rect 84699 68085 84747 68113
rect 84437 68051 84747 68085
rect 84437 68023 84485 68051
rect 84513 68023 84547 68051
rect 84575 68023 84609 68051
rect 84637 68023 84671 68051
rect 84699 68023 84747 68051
rect 84437 67989 84747 68023
rect 84437 67961 84485 67989
rect 84513 67961 84547 67989
rect 84575 67961 84609 67989
rect 84637 67961 84671 67989
rect 84699 67961 84747 67989
rect 82577 65147 82625 65175
rect 82653 65147 82687 65175
rect 82715 65147 82749 65175
rect 82777 65147 82811 65175
rect 82839 65147 82887 65175
rect 82577 65113 82887 65147
rect 82577 65085 82625 65113
rect 82653 65085 82687 65113
rect 82715 65085 82749 65113
rect 82777 65085 82811 65113
rect 82839 65085 82887 65113
rect 82577 65051 82887 65085
rect 82577 65023 82625 65051
rect 82653 65023 82687 65051
rect 82715 65023 82749 65051
rect 82777 65023 82811 65051
rect 82839 65023 82887 65051
rect 82577 64989 82887 65023
rect 82577 64961 82625 64989
rect 82653 64961 82687 64989
rect 82715 64961 82749 64989
rect 82777 64961 82811 64989
rect 82839 64961 82887 64989
rect 75437 59147 75485 59175
rect 75513 59147 75547 59175
rect 75575 59147 75609 59175
rect 75637 59147 75671 59175
rect 75699 59147 75747 59175
rect 75437 59113 75747 59147
rect 75437 59085 75485 59113
rect 75513 59085 75547 59113
rect 75575 59085 75609 59113
rect 75637 59085 75671 59113
rect 75699 59085 75747 59113
rect 75437 59051 75747 59085
rect 75437 59023 75485 59051
rect 75513 59023 75547 59051
rect 75575 59023 75609 59051
rect 75637 59023 75671 59051
rect 75699 59023 75747 59051
rect 75437 58989 75747 59023
rect 75437 58961 75485 58989
rect 75513 58961 75547 58989
rect 75575 58961 75609 58989
rect 75637 58961 75671 58989
rect 75699 58961 75747 58989
rect 73577 56147 73625 56175
rect 73653 56147 73687 56175
rect 73715 56147 73749 56175
rect 73777 56147 73811 56175
rect 73839 56147 73887 56175
rect 73577 56113 73887 56147
rect 73577 56085 73625 56113
rect 73653 56085 73687 56113
rect 73715 56085 73749 56113
rect 73777 56085 73811 56113
rect 73839 56085 73887 56113
rect 73577 56051 73887 56085
rect 73577 56023 73625 56051
rect 73653 56023 73687 56051
rect 73715 56023 73749 56051
rect 73777 56023 73811 56051
rect 73839 56023 73887 56051
rect 73577 55989 73887 56023
rect 73577 55961 73625 55989
rect 73653 55961 73687 55989
rect 73715 55961 73749 55989
rect 73777 55961 73811 55989
rect 73839 55961 73887 55989
rect 66437 50147 66485 50175
rect 66513 50147 66547 50175
rect 66575 50147 66609 50175
rect 66637 50147 66671 50175
rect 66699 50147 66747 50175
rect 66437 50113 66747 50147
rect 66437 50085 66485 50113
rect 66513 50085 66547 50113
rect 66575 50085 66609 50113
rect 66637 50085 66671 50113
rect 66699 50085 66747 50113
rect 66437 50051 66747 50085
rect 66437 50023 66485 50051
rect 66513 50023 66547 50051
rect 66575 50023 66609 50051
rect 66637 50023 66671 50051
rect 66699 50023 66747 50051
rect 66437 49989 66747 50023
rect 66437 49961 66485 49989
rect 66513 49961 66547 49989
rect 66575 49961 66609 49989
rect 66637 49961 66671 49989
rect 66699 49961 66747 49989
rect 66437 41175 66747 49961
rect 66437 41147 66485 41175
rect 66513 41147 66547 41175
rect 66575 41147 66609 41175
rect 66637 41147 66671 41175
rect 66699 41147 66747 41175
rect 66437 41113 66747 41147
rect 66437 41085 66485 41113
rect 66513 41085 66547 41113
rect 66575 41085 66609 41113
rect 66637 41085 66671 41113
rect 66699 41085 66747 41113
rect 66437 41051 66747 41085
rect 66437 41023 66485 41051
rect 66513 41023 66547 41051
rect 66575 41023 66609 41051
rect 66637 41023 66671 41051
rect 66699 41023 66747 41051
rect 66437 40989 66747 41023
rect 66437 40961 66485 40989
rect 66513 40961 66547 40989
rect 66575 40961 66609 40989
rect 66637 40961 66671 40989
rect 66699 40961 66747 40989
rect 66437 32175 66747 40961
rect 66437 32147 66485 32175
rect 66513 32147 66547 32175
rect 66575 32147 66609 32175
rect 66637 32147 66671 32175
rect 66699 32147 66747 32175
rect 66437 32113 66747 32147
rect 66437 32085 66485 32113
rect 66513 32085 66547 32113
rect 66575 32085 66609 32113
rect 66637 32085 66671 32113
rect 66699 32085 66747 32113
rect 66437 32051 66747 32085
rect 66437 32023 66485 32051
rect 66513 32023 66547 32051
rect 66575 32023 66609 32051
rect 66637 32023 66671 32051
rect 66699 32023 66747 32051
rect 66437 31989 66747 32023
rect 66437 31961 66485 31989
rect 66513 31961 66547 31989
rect 66575 31961 66609 31989
rect 66637 31961 66671 31989
rect 66699 31961 66747 31989
rect 66437 23175 66747 31961
rect 66437 23147 66485 23175
rect 66513 23147 66547 23175
rect 66575 23147 66609 23175
rect 66637 23147 66671 23175
rect 66699 23147 66747 23175
rect 66437 23113 66747 23147
rect 66437 23085 66485 23113
rect 66513 23085 66547 23113
rect 66575 23085 66609 23113
rect 66637 23085 66671 23113
rect 66699 23085 66747 23113
rect 66437 23051 66747 23085
rect 66437 23023 66485 23051
rect 66513 23023 66547 23051
rect 66575 23023 66609 23051
rect 66637 23023 66671 23051
rect 66699 23023 66747 23051
rect 66437 22989 66747 23023
rect 66437 22961 66485 22989
rect 66513 22961 66547 22989
rect 66575 22961 66609 22989
rect 66637 22961 66671 22989
rect 66699 22961 66747 22989
rect 66437 14175 66747 22961
rect 66437 14147 66485 14175
rect 66513 14147 66547 14175
rect 66575 14147 66609 14175
rect 66637 14147 66671 14175
rect 66699 14147 66747 14175
rect 66437 14113 66747 14147
rect 66437 14085 66485 14113
rect 66513 14085 66547 14113
rect 66575 14085 66609 14113
rect 66637 14085 66671 14113
rect 66699 14085 66747 14113
rect 66437 14051 66747 14085
rect 66437 14023 66485 14051
rect 66513 14023 66547 14051
rect 66575 14023 66609 14051
rect 66637 14023 66671 14051
rect 66699 14023 66747 14051
rect 66437 13989 66747 14023
rect 66437 13961 66485 13989
rect 66513 13961 66547 13989
rect 66575 13961 66609 13989
rect 66637 13961 66671 13989
rect 66699 13961 66747 13989
rect 66437 5175 66747 13961
rect 66437 5147 66485 5175
rect 66513 5147 66547 5175
rect 66575 5147 66609 5175
rect 66637 5147 66671 5175
rect 66699 5147 66747 5175
rect 66437 5113 66747 5147
rect 66437 5085 66485 5113
rect 66513 5085 66547 5113
rect 66575 5085 66609 5113
rect 66637 5085 66671 5113
rect 66699 5085 66747 5113
rect 66437 5051 66747 5085
rect 66437 5023 66485 5051
rect 66513 5023 66547 5051
rect 66575 5023 66609 5051
rect 66637 5023 66671 5051
rect 66699 5023 66747 5051
rect 66437 4989 66747 5023
rect 66437 4961 66485 4989
rect 66513 4961 66547 4989
rect 66575 4961 66609 4989
rect 66637 4961 66671 4989
rect 66699 4961 66747 4989
rect 66437 -560 66747 4961
rect 66437 -588 66485 -560
rect 66513 -588 66547 -560
rect 66575 -588 66609 -560
rect 66637 -588 66671 -560
rect 66699 -588 66747 -560
rect 66437 -622 66747 -588
rect 66437 -650 66485 -622
rect 66513 -650 66547 -622
rect 66575 -650 66609 -622
rect 66637 -650 66671 -622
rect 66699 -650 66747 -622
rect 66437 -684 66747 -650
rect 66437 -712 66485 -684
rect 66513 -712 66547 -684
rect 66575 -712 66609 -684
rect 66637 -712 66671 -684
rect 66699 -712 66747 -684
rect 66437 -746 66747 -712
rect 66437 -774 66485 -746
rect 66513 -774 66547 -746
rect 66575 -774 66609 -746
rect 66637 -774 66671 -746
rect 66699 -774 66747 -746
rect 66437 -822 66747 -774
rect 73577 47175 73887 55961
rect 74724 56175 74884 56192
rect 74724 56147 74759 56175
rect 74787 56147 74821 56175
rect 74849 56147 74884 56175
rect 74724 56113 74884 56147
rect 74724 56085 74759 56113
rect 74787 56085 74821 56113
rect 74849 56085 74884 56113
rect 74724 56051 74884 56085
rect 74724 56023 74759 56051
rect 74787 56023 74821 56051
rect 74849 56023 74884 56051
rect 74724 55989 74884 56023
rect 74724 55961 74759 55989
rect 74787 55961 74821 55989
rect 74849 55961 74884 55989
rect 74724 55944 74884 55961
rect 73577 47147 73625 47175
rect 73653 47147 73687 47175
rect 73715 47147 73749 47175
rect 73777 47147 73811 47175
rect 73839 47147 73887 47175
rect 73577 47113 73887 47147
rect 73577 47085 73625 47113
rect 73653 47085 73687 47113
rect 73715 47085 73749 47113
rect 73777 47085 73811 47113
rect 73839 47085 73887 47113
rect 73577 47051 73887 47085
rect 73577 47023 73625 47051
rect 73653 47023 73687 47051
rect 73715 47023 73749 47051
rect 73777 47023 73811 47051
rect 73839 47023 73887 47051
rect 73577 46989 73887 47023
rect 73577 46961 73625 46989
rect 73653 46961 73687 46989
rect 73715 46961 73749 46989
rect 73777 46961 73811 46989
rect 73839 46961 73887 46989
rect 73577 38175 73887 46961
rect 73577 38147 73625 38175
rect 73653 38147 73687 38175
rect 73715 38147 73749 38175
rect 73777 38147 73811 38175
rect 73839 38147 73887 38175
rect 73577 38113 73887 38147
rect 73577 38085 73625 38113
rect 73653 38085 73687 38113
rect 73715 38085 73749 38113
rect 73777 38085 73811 38113
rect 73839 38085 73887 38113
rect 73577 38051 73887 38085
rect 73577 38023 73625 38051
rect 73653 38023 73687 38051
rect 73715 38023 73749 38051
rect 73777 38023 73811 38051
rect 73839 38023 73887 38051
rect 73577 37989 73887 38023
rect 73577 37961 73625 37989
rect 73653 37961 73687 37989
rect 73715 37961 73749 37989
rect 73777 37961 73811 37989
rect 73839 37961 73887 37989
rect 73577 29175 73887 37961
rect 73577 29147 73625 29175
rect 73653 29147 73687 29175
rect 73715 29147 73749 29175
rect 73777 29147 73811 29175
rect 73839 29147 73887 29175
rect 73577 29113 73887 29147
rect 73577 29085 73625 29113
rect 73653 29085 73687 29113
rect 73715 29085 73749 29113
rect 73777 29085 73811 29113
rect 73839 29085 73887 29113
rect 73577 29051 73887 29085
rect 73577 29023 73625 29051
rect 73653 29023 73687 29051
rect 73715 29023 73749 29051
rect 73777 29023 73811 29051
rect 73839 29023 73887 29051
rect 73577 28989 73887 29023
rect 73577 28961 73625 28989
rect 73653 28961 73687 28989
rect 73715 28961 73749 28989
rect 73777 28961 73811 28989
rect 73839 28961 73887 28989
rect 73577 20175 73887 28961
rect 73577 20147 73625 20175
rect 73653 20147 73687 20175
rect 73715 20147 73749 20175
rect 73777 20147 73811 20175
rect 73839 20147 73887 20175
rect 73577 20113 73887 20147
rect 73577 20085 73625 20113
rect 73653 20085 73687 20113
rect 73715 20085 73749 20113
rect 73777 20085 73811 20113
rect 73839 20085 73887 20113
rect 73577 20051 73887 20085
rect 73577 20023 73625 20051
rect 73653 20023 73687 20051
rect 73715 20023 73749 20051
rect 73777 20023 73811 20051
rect 73839 20023 73887 20051
rect 73577 19989 73887 20023
rect 73577 19961 73625 19989
rect 73653 19961 73687 19989
rect 73715 19961 73749 19989
rect 73777 19961 73811 19989
rect 73839 19961 73887 19989
rect 73577 11175 73887 19961
rect 73577 11147 73625 11175
rect 73653 11147 73687 11175
rect 73715 11147 73749 11175
rect 73777 11147 73811 11175
rect 73839 11147 73887 11175
rect 73577 11113 73887 11147
rect 73577 11085 73625 11113
rect 73653 11085 73687 11113
rect 73715 11085 73749 11113
rect 73777 11085 73811 11113
rect 73839 11085 73887 11113
rect 73577 11051 73887 11085
rect 73577 11023 73625 11051
rect 73653 11023 73687 11051
rect 73715 11023 73749 11051
rect 73777 11023 73811 11051
rect 73839 11023 73887 11051
rect 73577 10989 73887 11023
rect 73577 10961 73625 10989
rect 73653 10961 73687 10989
rect 73715 10961 73749 10989
rect 73777 10961 73811 10989
rect 73839 10961 73887 10989
rect 73577 2175 73887 10961
rect 73577 2147 73625 2175
rect 73653 2147 73687 2175
rect 73715 2147 73749 2175
rect 73777 2147 73811 2175
rect 73839 2147 73887 2175
rect 73577 2113 73887 2147
rect 73577 2085 73625 2113
rect 73653 2085 73687 2113
rect 73715 2085 73749 2113
rect 73777 2085 73811 2113
rect 73839 2085 73887 2113
rect 73577 2051 73887 2085
rect 73577 2023 73625 2051
rect 73653 2023 73687 2051
rect 73715 2023 73749 2051
rect 73777 2023 73811 2051
rect 73839 2023 73887 2051
rect 73577 1989 73887 2023
rect 73577 1961 73625 1989
rect 73653 1961 73687 1989
rect 73715 1961 73749 1989
rect 73777 1961 73811 1989
rect 73839 1961 73887 1989
rect 73577 -80 73887 1961
rect 73577 -108 73625 -80
rect 73653 -108 73687 -80
rect 73715 -108 73749 -80
rect 73777 -108 73811 -80
rect 73839 -108 73887 -80
rect 73577 -142 73887 -108
rect 73577 -170 73625 -142
rect 73653 -170 73687 -142
rect 73715 -170 73749 -142
rect 73777 -170 73811 -142
rect 73839 -170 73887 -142
rect 73577 -204 73887 -170
rect 73577 -232 73625 -204
rect 73653 -232 73687 -204
rect 73715 -232 73749 -204
rect 73777 -232 73811 -204
rect 73839 -232 73887 -204
rect 73577 -266 73887 -232
rect 73577 -294 73625 -266
rect 73653 -294 73687 -266
rect 73715 -294 73749 -266
rect 73777 -294 73811 -266
rect 73839 -294 73887 -266
rect 73577 -822 73887 -294
rect 75437 50175 75747 58961
rect 76974 59175 77134 59192
rect 76974 59147 77009 59175
rect 77037 59147 77071 59175
rect 77099 59147 77134 59175
rect 76974 59113 77134 59147
rect 76974 59085 77009 59113
rect 77037 59085 77071 59113
rect 77099 59085 77134 59113
rect 76974 59051 77134 59085
rect 76974 59023 77009 59051
rect 77037 59023 77071 59051
rect 77099 59023 77134 59051
rect 76974 58989 77134 59023
rect 76974 58961 77009 58989
rect 77037 58961 77071 58989
rect 77099 58961 77134 58989
rect 76974 58944 77134 58961
rect 81474 59175 81634 59192
rect 81474 59147 81509 59175
rect 81537 59147 81571 59175
rect 81599 59147 81634 59175
rect 81474 59113 81634 59147
rect 81474 59085 81509 59113
rect 81537 59085 81571 59113
rect 81599 59085 81634 59113
rect 81474 59051 81634 59085
rect 81474 59023 81509 59051
rect 81537 59023 81571 59051
rect 81599 59023 81634 59051
rect 81474 58989 81634 59023
rect 81474 58961 81509 58989
rect 81537 58961 81571 58989
rect 81599 58961 81634 58989
rect 81474 58944 81634 58961
rect 79224 56175 79384 56192
rect 79224 56147 79259 56175
rect 79287 56147 79321 56175
rect 79349 56147 79384 56175
rect 79224 56113 79384 56147
rect 79224 56085 79259 56113
rect 79287 56085 79321 56113
rect 79349 56085 79384 56113
rect 79224 56051 79384 56085
rect 79224 56023 79259 56051
rect 79287 56023 79321 56051
rect 79349 56023 79384 56051
rect 79224 55989 79384 56023
rect 79224 55961 79259 55989
rect 79287 55961 79321 55989
rect 79349 55961 79384 55989
rect 79224 55944 79384 55961
rect 82577 56175 82887 64961
rect 83724 65175 83884 65192
rect 83724 65147 83759 65175
rect 83787 65147 83821 65175
rect 83849 65147 83884 65175
rect 83724 65113 83884 65147
rect 83724 65085 83759 65113
rect 83787 65085 83821 65113
rect 83849 65085 83884 65113
rect 83724 65051 83884 65085
rect 83724 65023 83759 65051
rect 83787 65023 83821 65051
rect 83849 65023 83884 65051
rect 83724 64989 83884 65023
rect 83724 64961 83759 64989
rect 83787 64961 83821 64989
rect 83849 64961 83884 64989
rect 83724 64944 83884 64961
rect 84437 59175 84747 67961
rect 85974 68175 86134 68192
rect 85974 68147 86009 68175
rect 86037 68147 86071 68175
rect 86099 68147 86134 68175
rect 85974 68113 86134 68147
rect 85974 68085 86009 68113
rect 86037 68085 86071 68113
rect 86099 68085 86134 68113
rect 85974 68051 86134 68085
rect 85974 68023 86009 68051
rect 86037 68023 86071 68051
rect 86099 68023 86134 68051
rect 85974 67989 86134 68023
rect 85974 67961 86009 67989
rect 86037 67961 86071 67989
rect 86099 67961 86134 67989
rect 85974 67944 86134 67961
rect 90474 68175 90634 68192
rect 90474 68147 90509 68175
rect 90537 68147 90571 68175
rect 90599 68147 90634 68175
rect 90474 68113 90634 68147
rect 90474 68085 90509 68113
rect 90537 68085 90571 68113
rect 90599 68085 90634 68113
rect 90474 68051 90634 68085
rect 90474 68023 90509 68051
rect 90537 68023 90571 68051
rect 90599 68023 90634 68051
rect 90474 67989 90634 68023
rect 90474 67961 90509 67989
rect 90537 67961 90571 67989
rect 90599 67961 90634 67989
rect 90474 67944 90634 67961
rect 88224 65175 88384 65192
rect 88224 65147 88259 65175
rect 88287 65147 88321 65175
rect 88349 65147 88384 65175
rect 88224 65113 88384 65147
rect 88224 65085 88259 65113
rect 88287 65085 88321 65113
rect 88349 65085 88384 65113
rect 88224 65051 88384 65085
rect 88224 65023 88259 65051
rect 88287 65023 88321 65051
rect 88349 65023 88384 65051
rect 88224 64989 88384 65023
rect 88224 64961 88259 64989
rect 88287 64961 88321 64989
rect 88349 64961 88384 64989
rect 88224 64944 88384 64961
rect 91577 65175 91887 73961
rect 92724 74175 92884 74192
rect 92724 74147 92759 74175
rect 92787 74147 92821 74175
rect 92849 74147 92884 74175
rect 92724 74113 92884 74147
rect 92724 74085 92759 74113
rect 92787 74085 92821 74113
rect 92849 74085 92884 74113
rect 92724 74051 92884 74085
rect 92724 74023 92759 74051
rect 92787 74023 92821 74051
rect 92849 74023 92884 74051
rect 92724 73989 92884 74023
rect 92724 73961 92759 73989
rect 92787 73961 92821 73989
rect 92849 73961 92884 73989
rect 92724 73944 92884 73961
rect 97224 74175 97384 74192
rect 97224 74147 97259 74175
rect 97287 74147 97321 74175
rect 97349 74147 97384 74175
rect 97224 74113 97384 74147
rect 97224 74085 97259 74113
rect 97287 74085 97321 74113
rect 97349 74085 97384 74113
rect 97224 74051 97384 74085
rect 97224 74023 97259 74051
rect 97287 74023 97321 74051
rect 97349 74023 97384 74051
rect 97224 73989 97384 74023
rect 97224 73961 97259 73989
rect 97287 73961 97321 73989
rect 97349 73961 97384 73989
rect 97224 73944 97384 73961
rect 101724 74175 101884 74192
rect 101724 74147 101759 74175
rect 101787 74147 101821 74175
rect 101849 74147 101884 74175
rect 101724 74113 101884 74147
rect 101724 74085 101759 74113
rect 101787 74085 101821 74113
rect 101849 74085 101884 74113
rect 101724 74051 101884 74085
rect 101724 74023 101759 74051
rect 101787 74023 101821 74051
rect 101849 74023 101884 74051
rect 101724 73989 101884 74023
rect 101724 73961 101759 73989
rect 101787 73961 101821 73989
rect 101849 73961 101884 73989
rect 101724 73944 101884 73961
rect 106224 74175 106384 74192
rect 106224 74147 106259 74175
rect 106287 74147 106321 74175
rect 106349 74147 106384 74175
rect 106224 74113 106384 74147
rect 106224 74085 106259 74113
rect 106287 74085 106321 74113
rect 106349 74085 106384 74113
rect 106224 74051 106384 74085
rect 106224 74023 106259 74051
rect 106287 74023 106321 74051
rect 106349 74023 106384 74051
rect 106224 73989 106384 74023
rect 106224 73961 106259 73989
rect 106287 73961 106321 73989
rect 106349 73961 106384 73989
rect 106224 73944 106384 73961
rect 110724 74175 110884 74192
rect 110724 74147 110759 74175
rect 110787 74147 110821 74175
rect 110849 74147 110884 74175
rect 110724 74113 110884 74147
rect 110724 74085 110759 74113
rect 110787 74085 110821 74113
rect 110849 74085 110884 74113
rect 110724 74051 110884 74085
rect 110724 74023 110759 74051
rect 110787 74023 110821 74051
rect 110849 74023 110884 74051
rect 110724 73989 110884 74023
rect 110724 73961 110759 73989
rect 110787 73961 110821 73989
rect 110849 73961 110884 73989
rect 110724 73944 110884 73961
rect 115224 74175 115384 74192
rect 115224 74147 115259 74175
rect 115287 74147 115321 74175
rect 115349 74147 115384 74175
rect 115224 74113 115384 74147
rect 115224 74085 115259 74113
rect 115287 74085 115321 74113
rect 115349 74085 115384 74113
rect 115224 74051 115384 74085
rect 115224 74023 115259 74051
rect 115287 74023 115321 74051
rect 115349 74023 115384 74051
rect 115224 73989 115384 74023
rect 115224 73961 115259 73989
rect 115287 73961 115321 73989
rect 115349 73961 115384 73989
rect 115224 73944 115384 73961
rect 94974 68175 95134 68192
rect 94974 68147 95009 68175
rect 95037 68147 95071 68175
rect 95099 68147 95134 68175
rect 94974 68113 95134 68147
rect 94974 68085 95009 68113
rect 95037 68085 95071 68113
rect 95099 68085 95134 68113
rect 94974 68051 95134 68085
rect 94974 68023 95009 68051
rect 95037 68023 95071 68051
rect 95099 68023 95134 68051
rect 94974 67989 95134 68023
rect 94974 67961 95009 67989
rect 95037 67961 95071 67989
rect 95099 67961 95134 67989
rect 94974 67944 95134 67961
rect 99474 68175 99634 68192
rect 99474 68147 99509 68175
rect 99537 68147 99571 68175
rect 99599 68147 99634 68175
rect 99474 68113 99634 68147
rect 99474 68085 99509 68113
rect 99537 68085 99571 68113
rect 99599 68085 99634 68113
rect 99474 68051 99634 68085
rect 99474 68023 99509 68051
rect 99537 68023 99571 68051
rect 99599 68023 99634 68051
rect 99474 67989 99634 68023
rect 99474 67961 99509 67989
rect 99537 67961 99571 67989
rect 99599 67961 99634 67989
rect 99474 67944 99634 67961
rect 103974 68175 104134 68192
rect 103974 68147 104009 68175
rect 104037 68147 104071 68175
rect 104099 68147 104134 68175
rect 103974 68113 104134 68147
rect 103974 68085 104009 68113
rect 104037 68085 104071 68113
rect 104099 68085 104134 68113
rect 103974 68051 104134 68085
rect 103974 68023 104009 68051
rect 104037 68023 104071 68051
rect 104099 68023 104134 68051
rect 103974 67989 104134 68023
rect 103974 67961 104009 67989
rect 104037 67961 104071 67989
rect 104099 67961 104134 67989
rect 103974 67944 104134 67961
rect 108474 68175 108634 68192
rect 108474 68147 108509 68175
rect 108537 68147 108571 68175
rect 108599 68147 108634 68175
rect 108474 68113 108634 68147
rect 108474 68085 108509 68113
rect 108537 68085 108571 68113
rect 108599 68085 108634 68113
rect 108474 68051 108634 68085
rect 108474 68023 108509 68051
rect 108537 68023 108571 68051
rect 108599 68023 108634 68051
rect 108474 67989 108634 68023
rect 108474 67961 108509 67989
rect 108537 67961 108571 67989
rect 108599 67961 108634 67989
rect 108474 67944 108634 67961
rect 112974 68175 113134 68192
rect 112974 68147 113009 68175
rect 113037 68147 113071 68175
rect 113099 68147 113134 68175
rect 112974 68113 113134 68147
rect 112974 68085 113009 68113
rect 113037 68085 113071 68113
rect 113099 68085 113134 68113
rect 112974 68051 113134 68085
rect 112974 68023 113009 68051
rect 113037 68023 113071 68051
rect 113099 68023 113134 68051
rect 112974 67989 113134 68023
rect 112974 67961 113009 67989
rect 113037 67961 113071 67989
rect 113099 67961 113134 67989
rect 112974 67944 113134 67961
rect 117474 68175 117634 68192
rect 117474 68147 117509 68175
rect 117537 68147 117571 68175
rect 117599 68147 117634 68175
rect 117474 68113 117634 68147
rect 117474 68085 117509 68113
rect 117537 68085 117571 68113
rect 117599 68085 117634 68113
rect 117474 68051 117634 68085
rect 117474 68023 117509 68051
rect 117537 68023 117571 68051
rect 117599 68023 117634 68051
rect 117474 67989 117634 68023
rect 117474 67961 117509 67989
rect 117537 67961 117571 67989
rect 117599 67961 117634 67989
rect 117474 67944 117634 67961
rect 120437 68175 120747 76961
rect 120437 68147 120485 68175
rect 120513 68147 120547 68175
rect 120575 68147 120609 68175
rect 120637 68147 120671 68175
rect 120699 68147 120747 68175
rect 120437 68113 120747 68147
rect 120437 68085 120485 68113
rect 120513 68085 120547 68113
rect 120575 68085 120609 68113
rect 120637 68085 120671 68113
rect 120699 68085 120747 68113
rect 120437 68051 120747 68085
rect 120437 68023 120485 68051
rect 120513 68023 120547 68051
rect 120575 68023 120609 68051
rect 120637 68023 120671 68051
rect 120699 68023 120747 68051
rect 120437 67989 120747 68023
rect 120437 67961 120485 67989
rect 120513 67961 120547 67989
rect 120575 67961 120609 67989
rect 120637 67961 120671 67989
rect 120699 67961 120747 67989
rect 91577 65147 91625 65175
rect 91653 65147 91687 65175
rect 91715 65147 91749 65175
rect 91777 65147 91811 65175
rect 91839 65147 91887 65175
rect 91577 65113 91887 65147
rect 91577 65085 91625 65113
rect 91653 65085 91687 65113
rect 91715 65085 91749 65113
rect 91777 65085 91811 65113
rect 91839 65085 91887 65113
rect 91577 65051 91887 65085
rect 91577 65023 91625 65051
rect 91653 65023 91687 65051
rect 91715 65023 91749 65051
rect 91777 65023 91811 65051
rect 91839 65023 91887 65051
rect 91577 64989 91887 65023
rect 91577 64961 91625 64989
rect 91653 64961 91687 64989
rect 91715 64961 91749 64989
rect 91777 64961 91811 64989
rect 91839 64961 91887 64989
rect 84437 59147 84485 59175
rect 84513 59147 84547 59175
rect 84575 59147 84609 59175
rect 84637 59147 84671 59175
rect 84699 59147 84747 59175
rect 84437 59113 84747 59147
rect 84437 59085 84485 59113
rect 84513 59085 84547 59113
rect 84575 59085 84609 59113
rect 84637 59085 84671 59113
rect 84699 59085 84747 59113
rect 84437 59051 84747 59085
rect 84437 59023 84485 59051
rect 84513 59023 84547 59051
rect 84575 59023 84609 59051
rect 84637 59023 84671 59051
rect 84699 59023 84747 59051
rect 84437 58989 84747 59023
rect 84437 58961 84485 58989
rect 84513 58961 84547 58989
rect 84575 58961 84609 58989
rect 84637 58961 84671 58989
rect 84699 58961 84747 58989
rect 82577 56147 82625 56175
rect 82653 56147 82687 56175
rect 82715 56147 82749 56175
rect 82777 56147 82811 56175
rect 82839 56147 82887 56175
rect 82577 56113 82887 56147
rect 82577 56085 82625 56113
rect 82653 56085 82687 56113
rect 82715 56085 82749 56113
rect 82777 56085 82811 56113
rect 82839 56085 82887 56113
rect 82577 56051 82887 56085
rect 82577 56023 82625 56051
rect 82653 56023 82687 56051
rect 82715 56023 82749 56051
rect 82777 56023 82811 56051
rect 82839 56023 82887 56051
rect 82577 55989 82887 56023
rect 82577 55961 82625 55989
rect 82653 55961 82687 55989
rect 82715 55961 82749 55989
rect 82777 55961 82811 55989
rect 82839 55961 82887 55989
rect 75437 50147 75485 50175
rect 75513 50147 75547 50175
rect 75575 50147 75609 50175
rect 75637 50147 75671 50175
rect 75699 50147 75747 50175
rect 75437 50113 75747 50147
rect 75437 50085 75485 50113
rect 75513 50085 75547 50113
rect 75575 50085 75609 50113
rect 75637 50085 75671 50113
rect 75699 50085 75747 50113
rect 75437 50051 75747 50085
rect 75437 50023 75485 50051
rect 75513 50023 75547 50051
rect 75575 50023 75609 50051
rect 75637 50023 75671 50051
rect 75699 50023 75747 50051
rect 75437 49989 75747 50023
rect 75437 49961 75485 49989
rect 75513 49961 75547 49989
rect 75575 49961 75609 49989
rect 75637 49961 75671 49989
rect 75699 49961 75747 49989
rect 75437 41175 75747 49961
rect 75437 41147 75485 41175
rect 75513 41147 75547 41175
rect 75575 41147 75609 41175
rect 75637 41147 75671 41175
rect 75699 41147 75747 41175
rect 75437 41113 75747 41147
rect 75437 41085 75485 41113
rect 75513 41085 75547 41113
rect 75575 41085 75609 41113
rect 75637 41085 75671 41113
rect 75699 41085 75747 41113
rect 75437 41051 75747 41085
rect 75437 41023 75485 41051
rect 75513 41023 75547 41051
rect 75575 41023 75609 41051
rect 75637 41023 75671 41051
rect 75699 41023 75747 41051
rect 75437 40989 75747 41023
rect 75437 40961 75485 40989
rect 75513 40961 75547 40989
rect 75575 40961 75609 40989
rect 75637 40961 75671 40989
rect 75699 40961 75747 40989
rect 75437 32175 75747 40961
rect 75437 32147 75485 32175
rect 75513 32147 75547 32175
rect 75575 32147 75609 32175
rect 75637 32147 75671 32175
rect 75699 32147 75747 32175
rect 75437 32113 75747 32147
rect 75437 32085 75485 32113
rect 75513 32085 75547 32113
rect 75575 32085 75609 32113
rect 75637 32085 75671 32113
rect 75699 32085 75747 32113
rect 75437 32051 75747 32085
rect 75437 32023 75485 32051
rect 75513 32023 75547 32051
rect 75575 32023 75609 32051
rect 75637 32023 75671 32051
rect 75699 32023 75747 32051
rect 75437 31989 75747 32023
rect 75437 31961 75485 31989
rect 75513 31961 75547 31989
rect 75575 31961 75609 31989
rect 75637 31961 75671 31989
rect 75699 31961 75747 31989
rect 75437 23175 75747 31961
rect 75437 23147 75485 23175
rect 75513 23147 75547 23175
rect 75575 23147 75609 23175
rect 75637 23147 75671 23175
rect 75699 23147 75747 23175
rect 75437 23113 75747 23147
rect 75437 23085 75485 23113
rect 75513 23085 75547 23113
rect 75575 23085 75609 23113
rect 75637 23085 75671 23113
rect 75699 23085 75747 23113
rect 75437 23051 75747 23085
rect 75437 23023 75485 23051
rect 75513 23023 75547 23051
rect 75575 23023 75609 23051
rect 75637 23023 75671 23051
rect 75699 23023 75747 23051
rect 75437 22989 75747 23023
rect 75437 22961 75485 22989
rect 75513 22961 75547 22989
rect 75575 22961 75609 22989
rect 75637 22961 75671 22989
rect 75699 22961 75747 22989
rect 75437 14175 75747 22961
rect 75437 14147 75485 14175
rect 75513 14147 75547 14175
rect 75575 14147 75609 14175
rect 75637 14147 75671 14175
rect 75699 14147 75747 14175
rect 75437 14113 75747 14147
rect 75437 14085 75485 14113
rect 75513 14085 75547 14113
rect 75575 14085 75609 14113
rect 75637 14085 75671 14113
rect 75699 14085 75747 14113
rect 75437 14051 75747 14085
rect 75437 14023 75485 14051
rect 75513 14023 75547 14051
rect 75575 14023 75609 14051
rect 75637 14023 75671 14051
rect 75699 14023 75747 14051
rect 75437 13989 75747 14023
rect 75437 13961 75485 13989
rect 75513 13961 75547 13989
rect 75575 13961 75609 13989
rect 75637 13961 75671 13989
rect 75699 13961 75747 13989
rect 75437 5175 75747 13961
rect 75437 5147 75485 5175
rect 75513 5147 75547 5175
rect 75575 5147 75609 5175
rect 75637 5147 75671 5175
rect 75699 5147 75747 5175
rect 75437 5113 75747 5147
rect 75437 5085 75485 5113
rect 75513 5085 75547 5113
rect 75575 5085 75609 5113
rect 75637 5085 75671 5113
rect 75699 5085 75747 5113
rect 75437 5051 75747 5085
rect 75437 5023 75485 5051
rect 75513 5023 75547 5051
rect 75575 5023 75609 5051
rect 75637 5023 75671 5051
rect 75699 5023 75747 5051
rect 75437 4989 75747 5023
rect 75437 4961 75485 4989
rect 75513 4961 75547 4989
rect 75575 4961 75609 4989
rect 75637 4961 75671 4989
rect 75699 4961 75747 4989
rect 75437 -560 75747 4961
rect 75437 -588 75485 -560
rect 75513 -588 75547 -560
rect 75575 -588 75609 -560
rect 75637 -588 75671 -560
rect 75699 -588 75747 -560
rect 75437 -622 75747 -588
rect 75437 -650 75485 -622
rect 75513 -650 75547 -622
rect 75575 -650 75609 -622
rect 75637 -650 75671 -622
rect 75699 -650 75747 -622
rect 75437 -684 75747 -650
rect 75437 -712 75485 -684
rect 75513 -712 75547 -684
rect 75575 -712 75609 -684
rect 75637 -712 75671 -684
rect 75699 -712 75747 -684
rect 75437 -746 75747 -712
rect 75437 -774 75485 -746
rect 75513 -774 75547 -746
rect 75575 -774 75609 -746
rect 75637 -774 75671 -746
rect 75699 -774 75747 -746
rect 75437 -822 75747 -774
rect 82577 47175 82887 55961
rect 83724 56175 83884 56192
rect 83724 56147 83759 56175
rect 83787 56147 83821 56175
rect 83849 56147 83884 56175
rect 83724 56113 83884 56147
rect 83724 56085 83759 56113
rect 83787 56085 83821 56113
rect 83849 56085 83884 56113
rect 83724 56051 83884 56085
rect 83724 56023 83759 56051
rect 83787 56023 83821 56051
rect 83849 56023 83884 56051
rect 83724 55989 83884 56023
rect 83724 55961 83759 55989
rect 83787 55961 83821 55989
rect 83849 55961 83884 55989
rect 83724 55944 83884 55961
rect 82577 47147 82625 47175
rect 82653 47147 82687 47175
rect 82715 47147 82749 47175
rect 82777 47147 82811 47175
rect 82839 47147 82887 47175
rect 82577 47113 82887 47147
rect 82577 47085 82625 47113
rect 82653 47085 82687 47113
rect 82715 47085 82749 47113
rect 82777 47085 82811 47113
rect 82839 47085 82887 47113
rect 82577 47051 82887 47085
rect 82577 47023 82625 47051
rect 82653 47023 82687 47051
rect 82715 47023 82749 47051
rect 82777 47023 82811 47051
rect 82839 47023 82887 47051
rect 82577 46989 82887 47023
rect 82577 46961 82625 46989
rect 82653 46961 82687 46989
rect 82715 46961 82749 46989
rect 82777 46961 82811 46989
rect 82839 46961 82887 46989
rect 82577 38175 82887 46961
rect 82577 38147 82625 38175
rect 82653 38147 82687 38175
rect 82715 38147 82749 38175
rect 82777 38147 82811 38175
rect 82839 38147 82887 38175
rect 82577 38113 82887 38147
rect 82577 38085 82625 38113
rect 82653 38085 82687 38113
rect 82715 38085 82749 38113
rect 82777 38085 82811 38113
rect 82839 38085 82887 38113
rect 82577 38051 82887 38085
rect 82577 38023 82625 38051
rect 82653 38023 82687 38051
rect 82715 38023 82749 38051
rect 82777 38023 82811 38051
rect 82839 38023 82887 38051
rect 82577 37989 82887 38023
rect 82577 37961 82625 37989
rect 82653 37961 82687 37989
rect 82715 37961 82749 37989
rect 82777 37961 82811 37989
rect 82839 37961 82887 37989
rect 82577 29175 82887 37961
rect 82577 29147 82625 29175
rect 82653 29147 82687 29175
rect 82715 29147 82749 29175
rect 82777 29147 82811 29175
rect 82839 29147 82887 29175
rect 82577 29113 82887 29147
rect 82577 29085 82625 29113
rect 82653 29085 82687 29113
rect 82715 29085 82749 29113
rect 82777 29085 82811 29113
rect 82839 29085 82887 29113
rect 82577 29051 82887 29085
rect 82577 29023 82625 29051
rect 82653 29023 82687 29051
rect 82715 29023 82749 29051
rect 82777 29023 82811 29051
rect 82839 29023 82887 29051
rect 82577 28989 82887 29023
rect 82577 28961 82625 28989
rect 82653 28961 82687 28989
rect 82715 28961 82749 28989
rect 82777 28961 82811 28989
rect 82839 28961 82887 28989
rect 82577 20175 82887 28961
rect 82577 20147 82625 20175
rect 82653 20147 82687 20175
rect 82715 20147 82749 20175
rect 82777 20147 82811 20175
rect 82839 20147 82887 20175
rect 82577 20113 82887 20147
rect 82577 20085 82625 20113
rect 82653 20085 82687 20113
rect 82715 20085 82749 20113
rect 82777 20085 82811 20113
rect 82839 20085 82887 20113
rect 82577 20051 82887 20085
rect 82577 20023 82625 20051
rect 82653 20023 82687 20051
rect 82715 20023 82749 20051
rect 82777 20023 82811 20051
rect 82839 20023 82887 20051
rect 82577 19989 82887 20023
rect 82577 19961 82625 19989
rect 82653 19961 82687 19989
rect 82715 19961 82749 19989
rect 82777 19961 82811 19989
rect 82839 19961 82887 19989
rect 82577 11175 82887 19961
rect 82577 11147 82625 11175
rect 82653 11147 82687 11175
rect 82715 11147 82749 11175
rect 82777 11147 82811 11175
rect 82839 11147 82887 11175
rect 82577 11113 82887 11147
rect 82577 11085 82625 11113
rect 82653 11085 82687 11113
rect 82715 11085 82749 11113
rect 82777 11085 82811 11113
rect 82839 11085 82887 11113
rect 82577 11051 82887 11085
rect 82577 11023 82625 11051
rect 82653 11023 82687 11051
rect 82715 11023 82749 11051
rect 82777 11023 82811 11051
rect 82839 11023 82887 11051
rect 82577 10989 82887 11023
rect 82577 10961 82625 10989
rect 82653 10961 82687 10989
rect 82715 10961 82749 10989
rect 82777 10961 82811 10989
rect 82839 10961 82887 10989
rect 82577 2175 82887 10961
rect 82577 2147 82625 2175
rect 82653 2147 82687 2175
rect 82715 2147 82749 2175
rect 82777 2147 82811 2175
rect 82839 2147 82887 2175
rect 82577 2113 82887 2147
rect 82577 2085 82625 2113
rect 82653 2085 82687 2113
rect 82715 2085 82749 2113
rect 82777 2085 82811 2113
rect 82839 2085 82887 2113
rect 82577 2051 82887 2085
rect 82577 2023 82625 2051
rect 82653 2023 82687 2051
rect 82715 2023 82749 2051
rect 82777 2023 82811 2051
rect 82839 2023 82887 2051
rect 82577 1989 82887 2023
rect 82577 1961 82625 1989
rect 82653 1961 82687 1989
rect 82715 1961 82749 1989
rect 82777 1961 82811 1989
rect 82839 1961 82887 1989
rect 82577 -80 82887 1961
rect 82577 -108 82625 -80
rect 82653 -108 82687 -80
rect 82715 -108 82749 -80
rect 82777 -108 82811 -80
rect 82839 -108 82887 -80
rect 82577 -142 82887 -108
rect 82577 -170 82625 -142
rect 82653 -170 82687 -142
rect 82715 -170 82749 -142
rect 82777 -170 82811 -142
rect 82839 -170 82887 -142
rect 82577 -204 82887 -170
rect 82577 -232 82625 -204
rect 82653 -232 82687 -204
rect 82715 -232 82749 -204
rect 82777 -232 82811 -204
rect 82839 -232 82887 -204
rect 82577 -266 82887 -232
rect 82577 -294 82625 -266
rect 82653 -294 82687 -266
rect 82715 -294 82749 -266
rect 82777 -294 82811 -266
rect 82839 -294 82887 -266
rect 82577 -822 82887 -294
rect 84437 50175 84747 58961
rect 85974 59175 86134 59192
rect 85974 59147 86009 59175
rect 86037 59147 86071 59175
rect 86099 59147 86134 59175
rect 85974 59113 86134 59147
rect 85974 59085 86009 59113
rect 86037 59085 86071 59113
rect 86099 59085 86134 59113
rect 85974 59051 86134 59085
rect 85974 59023 86009 59051
rect 86037 59023 86071 59051
rect 86099 59023 86134 59051
rect 85974 58989 86134 59023
rect 85974 58961 86009 58989
rect 86037 58961 86071 58989
rect 86099 58961 86134 58989
rect 85974 58944 86134 58961
rect 90474 59175 90634 59192
rect 90474 59147 90509 59175
rect 90537 59147 90571 59175
rect 90599 59147 90634 59175
rect 90474 59113 90634 59147
rect 90474 59085 90509 59113
rect 90537 59085 90571 59113
rect 90599 59085 90634 59113
rect 90474 59051 90634 59085
rect 90474 59023 90509 59051
rect 90537 59023 90571 59051
rect 90599 59023 90634 59051
rect 90474 58989 90634 59023
rect 90474 58961 90509 58989
rect 90537 58961 90571 58989
rect 90599 58961 90634 58989
rect 90474 58944 90634 58961
rect 88224 56175 88384 56192
rect 88224 56147 88259 56175
rect 88287 56147 88321 56175
rect 88349 56147 88384 56175
rect 88224 56113 88384 56147
rect 88224 56085 88259 56113
rect 88287 56085 88321 56113
rect 88349 56085 88384 56113
rect 88224 56051 88384 56085
rect 88224 56023 88259 56051
rect 88287 56023 88321 56051
rect 88349 56023 88384 56051
rect 88224 55989 88384 56023
rect 88224 55961 88259 55989
rect 88287 55961 88321 55989
rect 88349 55961 88384 55989
rect 88224 55944 88384 55961
rect 91577 56175 91887 64961
rect 92724 65175 92884 65192
rect 92724 65147 92759 65175
rect 92787 65147 92821 65175
rect 92849 65147 92884 65175
rect 92724 65113 92884 65147
rect 92724 65085 92759 65113
rect 92787 65085 92821 65113
rect 92849 65085 92884 65113
rect 92724 65051 92884 65085
rect 92724 65023 92759 65051
rect 92787 65023 92821 65051
rect 92849 65023 92884 65051
rect 92724 64989 92884 65023
rect 92724 64961 92759 64989
rect 92787 64961 92821 64989
rect 92849 64961 92884 64989
rect 92724 64944 92884 64961
rect 97224 65175 97384 65192
rect 97224 65147 97259 65175
rect 97287 65147 97321 65175
rect 97349 65147 97384 65175
rect 97224 65113 97384 65147
rect 97224 65085 97259 65113
rect 97287 65085 97321 65113
rect 97349 65085 97384 65113
rect 97224 65051 97384 65085
rect 97224 65023 97259 65051
rect 97287 65023 97321 65051
rect 97349 65023 97384 65051
rect 97224 64989 97384 65023
rect 97224 64961 97259 64989
rect 97287 64961 97321 64989
rect 97349 64961 97384 64989
rect 97224 64944 97384 64961
rect 101724 65175 101884 65192
rect 101724 65147 101759 65175
rect 101787 65147 101821 65175
rect 101849 65147 101884 65175
rect 101724 65113 101884 65147
rect 101724 65085 101759 65113
rect 101787 65085 101821 65113
rect 101849 65085 101884 65113
rect 101724 65051 101884 65085
rect 101724 65023 101759 65051
rect 101787 65023 101821 65051
rect 101849 65023 101884 65051
rect 101724 64989 101884 65023
rect 101724 64961 101759 64989
rect 101787 64961 101821 64989
rect 101849 64961 101884 64989
rect 101724 64944 101884 64961
rect 106224 65175 106384 65192
rect 106224 65147 106259 65175
rect 106287 65147 106321 65175
rect 106349 65147 106384 65175
rect 106224 65113 106384 65147
rect 106224 65085 106259 65113
rect 106287 65085 106321 65113
rect 106349 65085 106384 65113
rect 106224 65051 106384 65085
rect 106224 65023 106259 65051
rect 106287 65023 106321 65051
rect 106349 65023 106384 65051
rect 106224 64989 106384 65023
rect 106224 64961 106259 64989
rect 106287 64961 106321 64989
rect 106349 64961 106384 64989
rect 106224 64944 106384 64961
rect 110724 65175 110884 65192
rect 110724 65147 110759 65175
rect 110787 65147 110821 65175
rect 110849 65147 110884 65175
rect 110724 65113 110884 65147
rect 110724 65085 110759 65113
rect 110787 65085 110821 65113
rect 110849 65085 110884 65113
rect 110724 65051 110884 65085
rect 110724 65023 110759 65051
rect 110787 65023 110821 65051
rect 110849 65023 110884 65051
rect 110724 64989 110884 65023
rect 110724 64961 110759 64989
rect 110787 64961 110821 64989
rect 110849 64961 110884 64989
rect 110724 64944 110884 64961
rect 115224 65175 115384 65192
rect 115224 65147 115259 65175
rect 115287 65147 115321 65175
rect 115349 65147 115384 65175
rect 115224 65113 115384 65147
rect 115224 65085 115259 65113
rect 115287 65085 115321 65113
rect 115349 65085 115384 65113
rect 115224 65051 115384 65085
rect 115224 65023 115259 65051
rect 115287 65023 115321 65051
rect 115349 65023 115384 65051
rect 115224 64989 115384 65023
rect 115224 64961 115259 64989
rect 115287 64961 115321 64989
rect 115349 64961 115384 64989
rect 115224 64944 115384 64961
rect 94974 59175 95134 59192
rect 94974 59147 95009 59175
rect 95037 59147 95071 59175
rect 95099 59147 95134 59175
rect 94974 59113 95134 59147
rect 94974 59085 95009 59113
rect 95037 59085 95071 59113
rect 95099 59085 95134 59113
rect 94974 59051 95134 59085
rect 94974 59023 95009 59051
rect 95037 59023 95071 59051
rect 95099 59023 95134 59051
rect 94974 58989 95134 59023
rect 94974 58961 95009 58989
rect 95037 58961 95071 58989
rect 95099 58961 95134 58989
rect 94974 58944 95134 58961
rect 99474 59175 99634 59192
rect 99474 59147 99509 59175
rect 99537 59147 99571 59175
rect 99599 59147 99634 59175
rect 99474 59113 99634 59147
rect 99474 59085 99509 59113
rect 99537 59085 99571 59113
rect 99599 59085 99634 59113
rect 99474 59051 99634 59085
rect 99474 59023 99509 59051
rect 99537 59023 99571 59051
rect 99599 59023 99634 59051
rect 99474 58989 99634 59023
rect 99474 58961 99509 58989
rect 99537 58961 99571 58989
rect 99599 58961 99634 58989
rect 99474 58944 99634 58961
rect 103974 59175 104134 59192
rect 103974 59147 104009 59175
rect 104037 59147 104071 59175
rect 104099 59147 104134 59175
rect 103974 59113 104134 59147
rect 103974 59085 104009 59113
rect 104037 59085 104071 59113
rect 104099 59085 104134 59113
rect 103974 59051 104134 59085
rect 103974 59023 104009 59051
rect 104037 59023 104071 59051
rect 104099 59023 104134 59051
rect 103974 58989 104134 59023
rect 103974 58961 104009 58989
rect 104037 58961 104071 58989
rect 104099 58961 104134 58989
rect 103974 58944 104134 58961
rect 108474 59175 108634 59192
rect 108474 59147 108509 59175
rect 108537 59147 108571 59175
rect 108599 59147 108634 59175
rect 108474 59113 108634 59147
rect 108474 59085 108509 59113
rect 108537 59085 108571 59113
rect 108599 59085 108634 59113
rect 108474 59051 108634 59085
rect 108474 59023 108509 59051
rect 108537 59023 108571 59051
rect 108599 59023 108634 59051
rect 108474 58989 108634 59023
rect 108474 58961 108509 58989
rect 108537 58961 108571 58989
rect 108599 58961 108634 58989
rect 108474 58944 108634 58961
rect 112974 59175 113134 59192
rect 112974 59147 113009 59175
rect 113037 59147 113071 59175
rect 113099 59147 113134 59175
rect 112974 59113 113134 59147
rect 112974 59085 113009 59113
rect 113037 59085 113071 59113
rect 113099 59085 113134 59113
rect 112974 59051 113134 59085
rect 112974 59023 113009 59051
rect 113037 59023 113071 59051
rect 113099 59023 113134 59051
rect 112974 58989 113134 59023
rect 112974 58961 113009 58989
rect 113037 58961 113071 58989
rect 113099 58961 113134 58989
rect 112974 58944 113134 58961
rect 117474 59175 117634 59192
rect 117474 59147 117509 59175
rect 117537 59147 117571 59175
rect 117599 59147 117634 59175
rect 117474 59113 117634 59147
rect 117474 59085 117509 59113
rect 117537 59085 117571 59113
rect 117599 59085 117634 59113
rect 117474 59051 117634 59085
rect 117474 59023 117509 59051
rect 117537 59023 117571 59051
rect 117599 59023 117634 59051
rect 117474 58989 117634 59023
rect 117474 58961 117509 58989
rect 117537 58961 117571 58989
rect 117599 58961 117634 58989
rect 117474 58944 117634 58961
rect 120437 59175 120747 67961
rect 120437 59147 120485 59175
rect 120513 59147 120547 59175
rect 120575 59147 120609 59175
rect 120637 59147 120671 59175
rect 120699 59147 120747 59175
rect 120437 59113 120747 59147
rect 120437 59085 120485 59113
rect 120513 59085 120547 59113
rect 120575 59085 120609 59113
rect 120637 59085 120671 59113
rect 120699 59085 120747 59113
rect 120437 59051 120747 59085
rect 120437 59023 120485 59051
rect 120513 59023 120547 59051
rect 120575 59023 120609 59051
rect 120637 59023 120671 59051
rect 120699 59023 120747 59051
rect 120437 58989 120747 59023
rect 120437 58961 120485 58989
rect 120513 58961 120547 58989
rect 120575 58961 120609 58989
rect 120637 58961 120671 58989
rect 120699 58961 120747 58989
rect 91577 56147 91625 56175
rect 91653 56147 91687 56175
rect 91715 56147 91749 56175
rect 91777 56147 91811 56175
rect 91839 56147 91887 56175
rect 91577 56113 91887 56147
rect 91577 56085 91625 56113
rect 91653 56085 91687 56113
rect 91715 56085 91749 56113
rect 91777 56085 91811 56113
rect 91839 56085 91887 56113
rect 91577 56051 91887 56085
rect 91577 56023 91625 56051
rect 91653 56023 91687 56051
rect 91715 56023 91749 56051
rect 91777 56023 91811 56051
rect 91839 56023 91887 56051
rect 91577 55989 91887 56023
rect 91577 55961 91625 55989
rect 91653 55961 91687 55989
rect 91715 55961 91749 55989
rect 91777 55961 91811 55989
rect 91839 55961 91887 55989
rect 84437 50147 84485 50175
rect 84513 50147 84547 50175
rect 84575 50147 84609 50175
rect 84637 50147 84671 50175
rect 84699 50147 84747 50175
rect 84437 50113 84747 50147
rect 84437 50085 84485 50113
rect 84513 50085 84547 50113
rect 84575 50085 84609 50113
rect 84637 50085 84671 50113
rect 84699 50085 84747 50113
rect 84437 50051 84747 50085
rect 84437 50023 84485 50051
rect 84513 50023 84547 50051
rect 84575 50023 84609 50051
rect 84637 50023 84671 50051
rect 84699 50023 84747 50051
rect 84437 49989 84747 50023
rect 84437 49961 84485 49989
rect 84513 49961 84547 49989
rect 84575 49961 84609 49989
rect 84637 49961 84671 49989
rect 84699 49961 84747 49989
rect 84437 41175 84747 49961
rect 84437 41147 84485 41175
rect 84513 41147 84547 41175
rect 84575 41147 84609 41175
rect 84637 41147 84671 41175
rect 84699 41147 84747 41175
rect 84437 41113 84747 41147
rect 84437 41085 84485 41113
rect 84513 41085 84547 41113
rect 84575 41085 84609 41113
rect 84637 41085 84671 41113
rect 84699 41085 84747 41113
rect 84437 41051 84747 41085
rect 84437 41023 84485 41051
rect 84513 41023 84547 41051
rect 84575 41023 84609 41051
rect 84637 41023 84671 41051
rect 84699 41023 84747 41051
rect 84437 40989 84747 41023
rect 84437 40961 84485 40989
rect 84513 40961 84547 40989
rect 84575 40961 84609 40989
rect 84637 40961 84671 40989
rect 84699 40961 84747 40989
rect 84437 32175 84747 40961
rect 84437 32147 84485 32175
rect 84513 32147 84547 32175
rect 84575 32147 84609 32175
rect 84637 32147 84671 32175
rect 84699 32147 84747 32175
rect 84437 32113 84747 32147
rect 84437 32085 84485 32113
rect 84513 32085 84547 32113
rect 84575 32085 84609 32113
rect 84637 32085 84671 32113
rect 84699 32085 84747 32113
rect 84437 32051 84747 32085
rect 84437 32023 84485 32051
rect 84513 32023 84547 32051
rect 84575 32023 84609 32051
rect 84637 32023 84671 32051
rect 84699 32023 84747 32051
rect 84437 31989 84747 32023
rect 84437 31961 84485 31989
rect 84513 31961 84547 31989
rect 84575 31961 84609 31989
rect 84637 31961 84671 31989
rect 84699 31961 84747 31989
rect 84437 23175 84747 31961
rect 84437 23147 84485 23175
rect 84513 23147 84547 23175
rect 84575 23147 84609 23175
rect 84637 23147 84671 23175
rect 84699 23147 84747 23175
rect 84437 23113 84747 23147
rect 84437 23085 84485 23113
rect 84513 23085 84547 23113
rect 84575 23085 84609 23113
rect 84637 23085 84671 23113
rect 84699 23085 84747 23113
rect 84437 23051 84747 23085
rect 84437 23023 84485 23051
rect 84513 23023 84547 23051
rect 84575 23023 84609 23051
rect 84637 23023 84671 23051
rect 84699 23023 84747 23051
rect 84437 22989 84747 23023
rect 84437 22961 84485 22989
rect 84513 22961 84547 22989
rect 84575 22961 84609 22989
rect 84637 22961 84671 22989
rect 84699 22961 84747 22989
rect 84437 14175 84747 22961
rect 84437 14147 84485 14175
rect 84513 14147 84547 14175
rect 84575 14147 84609 14175
rect 84637 14147 84671 14175
rect 84699 14147 84747 14175
rect 84437 14113 84747 14147
rect 84437 14085 84485 14113
rect 84513 14085 84547 14113
rect 84575 14085 84609 14113
rect 84637 14085 84671 14113
rect 84699 14085 84747 14113
rect 84437 14051 84747 14085
rect 84437 14023 84485 14051
rect 84513 14023 84547 14051
rect 84575 14023 84609 14051
rect 84637 14023 84671 14051
rect 84699 14023 84747 14051
rect 84437 13989 84747 14023
rect 84437 13961 84485 13989
rect 84513 13961 84547 13989
rect 84575 13961 84609 13989
rect 84637 13961 84671 13989
rect 84699 13961 84747 13989
rect 84437 5175 84747 13961
rect 84437 5147 84485 5175
rect 84513 5147 84547 5175
rect 84575 5147 84609 5175
rect 84637 5147 84671 5175
rect 84699 5147 84747 5175
rect 84437 5113 84747 5147
rect 84437 5085 84485 5113
rect 84513 5085 84547 5113
rect 84575 5085 84609 5113
rect 84637 5085 84671 5113
rect 84699 5085 84747 5113
rect 84437 5051 84747 5085
rect 84437 5023 84485 5051
rect 84513 5023 84547 5051
rect 84575 5023 84609 5051
rect 84637 5023 84671 5051
rect 84699 5023 84747 5051
rect 84437 4989 84747 5023
rect 84437 4961 84485 4989
rect 84513 4961 84547 4989
rect 84575 4961 84609 4989
rect 84637 4961 84671 4989
rect 84699 4961 84747 4989
rect 84437 -560 84747 4961
rect 84437 -588 84485 -560
rect 84513 -588 84547 -560
rect 84575 -588 84609 -560
rect 84637 -588 84671 -560
rect 84699 -588 84747 -560
rect 84437 -622 84747 -588
rect 84437 -650 84485 -622
rect 84513 -650 84547 -622
rect 84575 -650 84609 -622
rect 84637 -650 84671 -622
rect 84699 -650 84747 -622
rect 84437 -684 84747 -650
rect 84437 -712 84485 -684
rect 84513 -712 84547 -684
rect 84575 -712 84609 -684
rect 84637 -712 84671 -684
rect 84699 -712 84747 -684
rect 84437 -746 84747 -712
rect 84437 -774 84485 -746
rect 84513 -774 84547 -746
rect 84575 -774 84609 -746
rect 84637 -774 84671 -746
rect 84699 -774 84747 -746
rect 84437 -822 84747 -774
rect 91577 47175 91887 55961
rect 92724 56175 92884 56192
rect 92724 56147 92759 56175
rect 92787 56147 92821 56175
rect 92849 56147 92884 56175
rect 92724 56113 92884 56147
rect 92724 56085 92759 56113
rect 92787 56085 92821 56113
rect 92849 56085 92884 56113
rect 92724 56051 92884 56085
rect 92724 56023 92759 56051
rect 92787 56023 92821 56051
rect 92849 56023 92884 56051
rect 92724 55989 92884 56023
rect 92724 55961 92759 55989
rect 92787 55961 92821 55989
rect 92849 55961 92884 55989
rect 92724 55944 92884 55961
rect 97224 56175 97384 56192
rect 97224 56147 97259 56175
rect 97287 56147 97321 56175
rect 97349 56147 97384 56175
rect 97224 56113 97384 56147
rect 97224 56085 97259 56113
rect 97287 56085 97321 56113
rect 97349 56085 97384 56113
rect 97224 56051 97384 56085
rect 97224 56023 97259 56051
rect 97287 56023 97321 56051
rect 97349 56023 97384 56051
rect 97224 55989 97384 56023
rect 97224 55961 97259 55989
rect 97287 55961 97321 55989
rect 97349 55961 97384 55989
rect 97224 55944 97384 55961
rect 101724 56175 101884 56192
rect 101724 56147 101759 56175
rect 101787 56147 101821 56175
rect 101849 56147 101884 56175
rect 101724 56113 101884 56147
rect 101724 56085 101759 56113
rect 101787 56085 101821 56113
rect 101849 56085 101884 56113
rect 101724 56051 101884 56085
rect 101724 56023 101759 56051
rect 101787 56023 101821 56051
rect 101849 56023 101884 56051
rect 101724 55989 101884 56023
rect 101724 55961 101759 55989
rect 101787 55961 101821 55989
rect 101849 55961 101884 55989
rect 101724 55944 101884 55961
rect 106224 56175 106384 56192
rect 106224 56147 106259 56175
rect 106287 56147 106321 56175
rect 106349 56147 106384 56175
rect 106224 56113 106384 56147
rect 106224 56085 106259 56113
rect 106287 56085 106321 56113
rect 106349 56085 106384 56113
rect 106224 56051 106384 56085
rect 106224 56023 106259 56051
rect 106287 56023 106321 56051
rect 106349 56023 106384 56051
rect 106224 55989 106384 56023
rect 106224 55961 106259 55989
rect 106287 55961 106321 55989
rect 106349 55961 106384 55989
rect 106224 55944 106384 55961
rect 110724 56175 110884 56192
rect 110724 56147 110759 56175
rect 110787 56147 110821 56175
rect 110849 56147 110884 56175
rect 110724 56113 110884 56147
rect 110724 56085 110759 56113
rect 110787 56085 110821 56113
rect 110849 56085 110884 56113
rect 110724 56051 110884 56085
rect 110724 56023 110759 56051
rect 110787 56023 110821 56051
rect 110849 56023 110884 56051
rect 110724 55989 110884 56023
rect 110724 55961 110759 55989
rect 110787 55961 110821 55989
rect 110849 55961 110884 55989
rect 110724 55944 110884 55961
rect 115224 56175 115384 56192
rect 115224 56147 115259 56175
rect 115287 56147 115321 56175
rect 115349 56147 115384 56175
rect 115224 56113 115384 56147
rect 115224 56085 115259 56113
rect 115287 56085 115321 56113
rect 115349 56085 115384 56113
rect 115224 56051 115384 56085
rect 115224 56023 115259 56051
rect 115287 56023 115321 56051
rect 115349 56023 115384 56051
rect 115224 55989 115384 56023
rect 115224 55961 115259 55989
rect 115287 55961 115321 55989
rect 115349 55961 115384 55989
rect 115224 55944 115384 55961
rect 120437 50175 120747 58961
rect 120437 50147 120485 50175
rect 120513 50147 120547 50175
rect 120575 50147 120609 50175
rect 120637 50147 120671 50175
rect 120699 50147 120747 50175
rect 120437 50113 120747 50147
rect 120437 50085 120485 50113
rect 120513 50085 120547 50113
rect 120575 50085 120609 50113
rect 120637 50085 120671 50113
rect 120699 50085 120747 50113
rect 120437 50051 120747 50085
rect 120437 50023 120485 50051
rect 120513 50023 120547 50051
rect 120575 50023 120609 50051
rect 120637 50023 120671 50051
rect 120699 50023 120747 50051
rect 120437 49989 120747 50023
rect 120437 49961 120485 49989
rect 120513 49961 120547 49989
rect 120575 49961 120609 49989
rect 120637 49961 120671 49989
rect 120699 49961 120747 49989
rect 91577 47147 91625 47175
rect 91653 47147 91687 47175
rect 91715 47147 91749 47175
rect 91777 47147 91811 47175
rect 91839 47147 91887 47175
rect 91577 47113 91887 47147
rect 91577 47085 91625 47113
rect 91653 47085 91687 47113
rect 91715 47085 91749 47113
rect 91777 47085 91811 47113
rect 91839 47085 91887 47113
rect 91577 47051 91887 47085
rect 91577 47023 91625 47051
rect 91653 47023 91687 47051
rect 91715 47023 91749 47051
rect 91777 47023 91811 47051
rect 91839 47023 91887 47051
rect 91577 46989 91887 47023
rect 91577 46961 91625 46989
rect 91653 46961 91687 46989
rect 91715 46961 91749 46989
rect 91777 46961 91811 46989
rect 91839 46961 91887 46989
rect 91577 38175 91887 46961
rect 91577 38147 91625 38175
rect 91653 38147 91687 38175
rect 91715 38147 91749 38175
rect 91777 38147 91811 38175
rect 91839 38147 91887 38175
rect 91577 38113 91887 38147
rect 91577 38085 91625 38113
rect 91653 38085 91687 38113
rect 91715 38085 91749 38113
rect 91777 38085 91811 38113
rect 91839 38085 91887 38113
rect 91577 38051 91887 38085
rect 91577 38023 91625 38051
rect 91653 38023 91687 38051
rect 91715 38023 91749 38051
rect 91777 38023 91811 38051
rect 91839 38023 91887 38051
rect 91577 37989 91887 38023
rect 91577 37961 91625 37989
rect 91653 37961 91687 37989
rect 91715 37961 91749 37989
rect 91777 37961 91811 37989
rect 91839 37961 91887 37989
rect 91577 29175 91887 37961
rect 91577 29147 91625 29175
rect 91653 29147 91687 29175
rect 91715 29147 91749 29175
rect 91777 29147 91811 29175
rect 91839 29147 91887 29175
rect 91577 29113 91887 29147
rect 91577 29085 91625 29113
rect 91653 29085 91687 29113
rect 91715 29085 91749 29113
rect 91777 29085 91811 29113
rect 91839 29085 91887 29113
rect 91577 29051 91887 29085
rect 91577 29023 91625 29051
rect 91653 29023 91687 29051
rect 91715 29023 91749 29051
rect 91777 29023 91811 29051
rect 91839 29023 91887 29051
rect 91577 28989 91887 29023
rect 91577 28961 91625 28989
rect 91653 28961 91687 28989
rect 91715 28961 91749 28989
rect 91777 28961 91811 28989
rect 91839 28961 91887 28989
rect 91577 20175 91887 28961
rect 91577 20147 91625 20175
rect 91653 20147 91687 20175
rect 91715 20147 91749 20175
rect 91777 20147 91811 20175
rect 91839 20147 91887 20175
rect 91577 20113 91887 20147
rect 91577 20085 91625 20113
rect 91653 20085 91687 20113
rect 91715 20085 91749 20113
rect 91777 20085 91811 20113
rect 91839 20085 91887 20113
rect 91577 20051 91887 20085
rect 91577 20023 91625 20051
rect 91653 20023 91687 20051
rect 91715 20023 91749 20051
rect 91777 20023 91811 20051
rect 91839 20023 91887 20051
rect 91577 19989 91887 20023
rect 91577 19961 91625 19989
rect 91653 19961 91687 19989
rect 91715 19961 91749 19989
rect 91777 19961 91811 19989
rect 91839 19961 91887 19989
rect 91577 11175 91887 19961
rect 91577 11147 91625 11175
rect 91653 11147 91687 11175
rect 91715 11147 91749 11175
rect 91777 11147 91811 11175
rect 91839 11147 91887 11175
rect 91577 11113 91887 11147
rect 91577 11085 91625 11113
rect 91653 11085 91687 11113
rect 91715 11085 91749 11113
rect 91777 11085 91811 11113
rect 91839 11085 91887 11113
rect 91577 11051 91887 11085
rect 91577 11023 91625 11051
rect 91653 11023 91687 11051
rect 91715 11023 91749 11051
rect 91777 11023 91811 11051
rect 91839 11023 91887 11051
rect 91577 10989 91887 11023
rect 91577 10961 91625 10989
rect 91653 10961 91687 10989
rect 91715 10961 91749 10989
rect 91777 10961 91811 10989
rect 91839 10961 91887 10989
rect 91577 2175 91887 10961
rect 91577 2147 91625 2175
rect 91653 2147 91687 2175
rect 91715 2147 91749 2175
rect 91777 2147 91811 2175
rect 91839 2147 91887 2175
rect 91577 2113 91887 2147
rect 91577 2085 91625 2113
rect 91653 2085 91687 2113
rect 91715 2085 91749 2113
rect 91777 2085 91811 2113
rect 91839 2085 91887 2113
rect 91577 2051 91887 2085
rect 91577 2023 91625 2051
rect 91653 2023 91687 2051
rect 91715 2023 91749 2051
rect 91777 2023 91811 2051
rect 91839 2023 91887 2051
rect 91577 1989 91887 2023
rect 91577 1961 91625 1989
rect 91653 1961 91687 1989
rect 91715 1961 91749 1989
rect 91777 1961 91811 1989
rect 91839 1961 91887 1989
rect 91577 -80 91887 1961
rect 91577 -108 91625 -80
rect 91653 -108 91687 -80
rect 91715 -108 91749 -80
rect 91777 -108 91811 -80
rect 91839 -108 91887 -80
rect 91577 -142 91887 -108
rect 91577 -170 91625 -142
rect 91653 -170 91687 -142
rect 91715 -170 91749 -142
rect 91777 -170 91811 -142
rect 91839 -170 91887 -142
rect 91577 -204 91887 -170
rect 91577 -232 91625 -204
rect 91653 -232 91687 -204
rect 91715 -232 91749 -204
rect 91777 -232 91811 -204
rect 91839 -232 91887 -204
rect 91577 -266 91887 -232
rect 91577 -294 91625 -266
rect 91653 -294 91687 -266
rect 91715 -294 91749 -266
rect 91777 -294 91811 -266
rect 91839 -294 91887 -266
rect 91577 -822 91887 -294
rect 93437 41175 93747 49317
rect 93437 41147 93485 41175
rect 93513 41147 93547 41175
rect 93575 41147 93609 41175
rect 93637 41147 93671 41175
rect 93699 41147 93747 41175
rect 93437 41113 93747 41147
rect 93437 41085 93485 41113
rect 93513 41085 93547 41113
rect 93575 41085 93609 41113
rect 93637 41085 93671 41113
rect 93699 41085 93747 41113
rect 93437 41051 93747 41085
rect 93437 41023 93485 41051
rect 93513 41023 93547 41051
rect 93575 41023 93609 41051
rect 93637 41023 93671 41051
rect 93699 41023 93747 41051
rect 93437 40989 93747 41023
rect 93437 40961 93485 40989
rect 93513 40961 93547 40989
rect 93575 40961 93609 40989
rect 93637 40961 93671 40989
rect 93699 40961 93747 40989
rect 93437 32175 93747 40961
rect 93437 32147 93485 32175
rect 93513 32147 93547 32175
rect 93575 32147 93609 32175
rect 93637 32147 93671 32175
rect 93699 32147 93747 32175
rect 93437 32113 93747 32147
rect 93437 32085 93485 32113
rect 93513 32085 93547 32113
rect 93575 32085 93609 32113
rect 93637 32085 93671 32113
rect 93699 32085 93747 32113
rect 93437 32051 93747 32085
rect 93437 32023 93485 32051
rect 93513 32023 93547 32051
rect 93575 32023 93609 32051
rect 93637 32023 93671 32051
rect 93699 32023 93747 32051
rect 93437 31989 93747 32023
rect 93437 31961 93485 31989
rect 93513 31961 93547 31989
rect 93575 31961 93609 31989
rect 93637 31961 93671 31989
rect 93699 31961 93747 31989
rect 93437 23175 93747 31961
rect 93437 23147 93485 23175
rect 93513 23147 93547 23175
rect 93575 23147 93609 23175
rect 93637 23147 93671 23175
rect 93699 23147 93747 23175
rect 93437 23113 93747 23147
rect 93437 23085 93485 23113
rect 93513 23085 93547 23113
rect 93575 23085 93609 23113
rect 93637 23085 93671 23113
rect 93699 23085 93747 23113
rect 93437 23051 93747 23085
rect 93437 23023 93485 23051
rect 93513 23023 93547 23051
rect 93575 23023 93609 23051
rect 93637 23023 93671 23051
rect 93699 23023 93747 23051
rect 93437 22989 93747 23023
rect 93437 22961 93485 22989
rect 93513 22961 93547 22989
rect 93575 22961 93609 22989
rect 93637 22961 93671 22989
rect 93699 22961 93747 22989
rect 93437 14175 93747 22961
rect 93437 14147 93485 14175
rect 93513 14147 93547 14175
rect 93575 14147 93609 14175
rect 93637 14147 93671 14175
rect 93699 14147 93747 14175
rect 93437 14113 93747 14147
rect 93437 14085 93485 14113
rect 93513 14085 93547 14113
rect 93575 14085 93609 14113
rect 93637 14085 93671 14113
rect 93699 14085 93747 14113
rect 93437 14051 93747 14085
rect 93437 14023 93485 14051
rect 93513 14023 93547 14051
rect 93575 14023 93609 14051
rect 93637 14023 93671 14051
rect 93699 14023 93747 14051
rect 93437 13989 93747 14023
rect 93437 13961 93485 13989
rect 93513 13961 93547 13989
rect 93575 13961 93609 13989
rect 93637 13961 93671 13989
rect 93699 13961 93747 13989
rect 93437 5175 93747 13961
rect 93437 5147 93485 5175
rect 93513 5147 93547 5175
rect 93575 5147 93609 5175
rect 93637 5147 93671 5175
rect 93699 5147 93747 5175
rect 93437 5113 93747 5147
rect 93437 5085 93485 5113
rect 93513 5085 93547 5113
rect 93575 5085 93609 5113
rect 93637 5085 93671 5113
rect 93699 5085 93747 5113
rect 93437 5051 93747 5085
rect 93437 5023 93485 5051
rect 93513 5023 93547 5051
rect 93575 5023 93609 5051
rect 93637 5023 93671 5051
rect 93699 5023 93747 5051
rect 93437 4989 93747 5023
rect 93437 4961 93485 4989
rect 93513 4961 93547 4989
rect 93575 4961 93609 4989
rect 93637 4961 93671 4989
rect 93699 4961 93747 4989
rect 93437 -560 93747 4961
rect 93437 -588 93485 -560
rect 93513 -588 93547 -560
rect 93575 -588 93609 -560
rect 93637 -588 93671 -560
rect 93699 -588 93747 -560
rect 93437 -622 93747 -588
rect 93437 -650 93485 -622
rect 93513 -650 93547 -622
rect 93575 -650 93609 -622
rect 93637 -650 93671 -622
rect 93699 -650 93747 -622
rect 93437 -684 93747 -650
rect 93437 -712 93485 -684
rect 93513 -712 93547 -684
rect 93575 -712 93609 -684
rect 93637 -712 93671 -684
rect 93699 -712 93747 -684
rect 93437 -746 93747 -712
rect 93437 -774 93485 -746
rect 93513 -774 93547 -746
rect 93575 -774 93609 -746
rect 93637 -774 93671 -746
rect 93699 -774 93747 -746
rect 93437 -822 93747 -774
rect 100577 47175 100887 49317
rect 100577 47147 100625 47175
rect 100653 47147 100687 47175
rect 100715 47147 100749 47175
rect 100777 47147 100811 47175
rect 100839 47147 100887 47175
rect 100577 47113 100887 47147
rect 100577 47085 100625 47113
rect 100653 47085 100687 47113
rect 100715 47085 100749 47113
rect 100777 47085 100811 47113
rect 100839 47085 100887 47113
rect 100577 47051 100887 47085
rect 100577 47023 100625 47051
rect 100653 47023 100687 47051
rect 100715 47023 100749 47051
rect 100777 47023 100811 47051
rect 100839 47023 100887 47051
rect 100577 46989 100887 47023
rect 100577 46961 100625 46989
rect 100653 46961 100687 46989
rect 100715 46961 100749 46989
rect 100777 46961 100811 46989
rect 100839 46961 100887 46989
rect 100577 38175 100887 46961
rect 100577 38147 100625 38175
rect 100653 38147 100687 38175
rect 100715 38147 100749 38175
rect 100777 38147 100811 38175
rect 100839 38147 100887 38175
rect 100577 38113 100887 38147
rect 100577 38085 100625 38113
rect 100653 38085 100687 38113
rect 100715 38085 100749 38113
rect 100777 38085 100811 38113
rect 100839 38085 100887 38113
rect 100577 38051 100887 38085
rect 100577 38023 100625 38051
rect 100653 38023 100687 38051
rect 100715 38023 100749 38051
rect 100777 38023 100811 38051
rect 100839 38023 100887 38051
rect 100577 37989 100887 38023
rect 100577 37961 100625 37989
rect 100653 37961 100687 37989
rect 100715 37961 100749 37989
rect 100777 37961 100811 37989
rect 100839 37961 100887 37989
rect 100577 29175 100887 37961
rect 100577 29147 100625 29175
rect 100653 29147 100687 29175
rect 100715 29147 100749 29175
rect 100777 29147 100811 29175
rect 100839 29147 100887 29175
rect 100577 29113 100887 29147
rect 100577 29085 100625 29113
rect 100653 29085 100687 29113
rect 100715 29085 100749 29113
rect 100777 29085 100811 29113
rect 100839 29085 100887 29113
rect 100577 29051 100887 29085
rect 100577 29023 100625 29051
rect 100653 29023 100687 29051
rect 100715 29023 100749 29051
rect 100777 29023 100811 29051
rect 100839 29023 100887 29051
rect 100577 28989 100887 29023
rect 100577 28961 100625 28989
rect 100653 28961 100687 28989
rect 100715 28961 100749 28989
rect 100777 28961 100811 28989
rect 100839 28961 100887 28989
rect 100577 20175 100887 28961
rect 100577 20147 100625 20175
rect 100653 20147 100687 20175
rect 100715 20147 100749 20175
rect 100777 20147 100811 20175
rect 100839 20147 100887 20175
rect 100577 20113 100887 20147
rect 100577 20085 100625 20113
rect 100653 20085 100687 20113
rect 100715 20085 100749 20113
rect 100777 20085 100811 20113
rect 100839 20085 100887 20113
rect 100577 20051 100887 20085
rect 100577 20023 100625 20051
rect 100653 20023 100687 20051
rect 100715 20023 100749 20051
rect 100777 20023 100811 20051
rect 100839 20023 100887 20051
rect 100577 19989 100887 20023
rect 100577 19961 100625 19989
rect 100653 19961 100687 19989
rect 100715 19961 100749 19989
rect 100777 19961 100811 19989
rect 100839 19961 100887 19989
rect 100577 11175 100887 19961
rect 100577 11147 100625 11175
rect 100653 11147 100687 11175
rect 100715 11147 100749 11175
rect 100777 11147 100811 11175
rect 100839 11147 100887 11175
rect 100577 11113 100887 11147
rect 100577 11085 100625 11113
rect 100653 11085 100687 11113
rect 100715 11085 100749 11113
rect 100777 11085 100811 11113
rect 100839 11085 100887 11113
rect 100577 11051 100887 11085
rect 100577 11023 100625 11051
rect 100653 11023 100687 11051
rect 100715 11023 100749 11051
rect 100777 11023 100811 11051
rect 100839 11023 100887 11051
rect 100577 10989 100887 11023
rect 100577 10961 100625 10989
rect 100653 10961 100687 10989
rect 100715 10961 100749 10989
rect 100777 10961 100811 10989
rect 100839 10961 100887 10989
rect 100577 2175 100887 10961
rect 100577 2147 100625 2175
rect 100653 2147 100687 2175
rect 100715 2147 100749 2175
rect 100777 2147 100811 2175
rect 100839 2147 100887 2175
rect 100577 2113 100887 2147
rect 100577 2085 100625 2113
rect 100653 2085 100687 2113
rect 100715 2085 100749 2113
rect 100777 2085 100811 2113
rect 100839 2085 100887 2113
rect 100577 2051 100887 2085
rect 100577 2023 100625 2051
rect 100653 2023 100687 2051
rect 100715 2023 100749 2051
rect 100777 2023 100811 2051
rect 100839 2023 100887 2051
rect 100577 1989 100887 2023
rect 100577 1961 100625 1989
rect 100653 1961 100687 1989
rect 100715 1961 100749 1989
rect 100777 1961 100811 1989
rect 100839 1961 100887 1989
rect 100577 -80 100887 1961
rect 100577 -108 100625 -80
rect 100653 -108 100687 -80
rect 100715 -108 100749 -80
rect 100777 -108 100811 -80
rect 100839 -108 100887 -80
rect 100577 -142 100887 -108
rect 100577 -170 100625 -142
rect 100653 -170 100687 -142
rect 100715 -170 100749 -142
rect 100777 -170 100811 -142
rect 100839 -170 100887 -142
rect 100577 -204 100887 -170
rect 100577 -232 100625 -204
rect 100653 -232 100687 -204
rect 100715 -232 100749 -204
rect 100777 -232 100811 -204
rect 100839 -232 100887 -204
rect 100577 -266 100887 -232
rect 100577 -294 100625 -266
rect 100653 -294 100687 -266
rect 100715 -294 100749 -266
rect 100777 -294 100811 -266
rect 100839 -294 100887 -266
rect 100577 -822 100887 -294
rect 102437 41175 102747 49317
rect 102437 41147 102485 41175
rect 102513 41147 102547 41175
rect 102575 41147 102609 41175
rect 102637 41147 102671 41175
rect 102699 41147 102747 41175
rect 102437 41113 102747 41147
rect 102437 41085 102485 41113
rect 102513 41085 102547 41113
rect 102575 41085 102609 41113
rect 102637 41085 102671 41113
rect 102699 41085 102747 41113
rect 102437 41051 102747 41085
rect 102437 41023 102485 41051
rect 102513 41023 102547 41051
rect 102575 41023 102609 41051
rect 102637 41023 102671 41051
rect 102699 41023 102747 41051
rect 102437 40989 102747 41023
rect 102437 40961 102485 40989
rect 102513 40961 102547 40989
rect 102575 40961 102609 40989
rect 102637 40961 102671 40989
rect 102699 40961 102747 40989
rect 102437 32175 102747 40961
rect 102437 32147 102485 32175
rect 102513 32147 102547 32175
rect 102575 32147 102609 32175
rect 102637 32147 102671 32175
rect 102699 32147 102747 32175
rect 102437 32113 102747 32147
rect 102437 32085 102485 32113
rect 102513 32085 102547 32113
rect 102575 32085 102609 32113
rect 102637 32085 102671 32113
rect 102699 32085 102747 32113
rect 102437 32051 102747 32085
rect 102437 32023 102485 32051
rect 102513 32023 102547 32051
rect 102575 32023 102609 32051
rect 102637 32023 102671 32051
rect 102699 32023 102747 32051
rect 102437 31989 102747 32023
rect 102437 31961 102485 31989
rect 102513 31961 102547 31989
rect 102575 31961 102609 31989
rect 102637 31961 102671 31989
rect 102699 31961 102747 31989
rect 102437 23175 102747 31961
rect 102437 23147 102485 23175
rect 102513 23147 102547 23175
rect 102575 23147 102609 23175
rect 102637 23147 102671 23175
rect 102699 23147 102747 23175
rect 102437 23113 102747 23147
rect 102437 23085 102485 23113
rect 102513 23085 102547 23113
rect 102575 23085 102609 23113
rect 102637 23085 102671 23113
rect 102699 23085 102747 23113
rect 102437 23051 102747 23085
rect 102437 23023 102485 23051
rect 102513 23023 102547 23051
rect 102575 23023 102609 23051
rect 102637 23023 102671 23051
rect 102699 23023 102747 23051
rect 102437 22989 102747 23023
rect 102437 22961 102485 22989
rect 102513 22961 102547 22989
rect 102575 22961 102609 22989
rect 102637 22961 102671 22989
rect 102699 22961 102747 22989
rect 102437 14175 102747 22961
rect 102437 14147 102485 14175
rect 102513 14147 102547 14175
rect 102575 14147 102609 14175
rect 102637 14147 102671 14175
rect 102699 14147 102747 14175
rect 102437 14113 102747 14147
rect 102437 14085 102485 14113
rect 102513 14085 102547 14113
rect 102575 14085 102609 14113
rect 102637 14085 102671 14113
rect 102699 14085 102747 14113
rect 102437 14051 102747 14085
rect 102437 14023 102485 14051
rect 102513 14023 102547 14051
rect 102575 14023 102609 14051
rect 102637 14023 102671 14051
rect 102699 14023 102747 14051
rect 102437 13989 102747 14023
rect 102437 13961 102485 13989
rect 102513 13961 102547 13989
rect 102575 13961 102609 13989
rect 102637 13961 102671 13989
rect 102699 13961 102747 13989
rect 102437 5175 102747 13961
rect 102437 5147 102485 5175
rect 102513 5147 102547 5175
rect 102575 5147 102609 5175
rect 102637 5147 102671 5175
rect 102699 5147 102747 5175
rect 102437 5113 102747 5147
rect 102437 5085 102485 5113
rect 102513 5085 102547 5113
rect 102575 5085 102609 5113
rect 102637 5085 102671 5113
rect 102699 5085 102747 5113
rect 102437 5051 102747 5085
rect 102437 5023 102485 5051
rect 102513 5023 102547 5051
rect 102575 5023 102609 5051
rect 102637 5023 102671 5051
rect 102699 5023 102747 5051
rect 102437 4989 102747 5023
rect 102437 4961 102485 4989
rect 102513 4961 102547 4989
rect 102575 4961 102609 4989
rect 102637 4961 102671 4989
rect 102699 4961 102747 4989
rect 102437 -560 102747 4961
rect 102437 -588 102485 -560
rect 102513 -588 102547 -560
rect 102575 -588 102609 -560
rect 102637 -588 102671 -560
rect 102699 -588 102747 -560
rect 102437 -622 102747 -588
rect 102437 -650 102485 -622
rect 102513 -650 102547 -622
rect 102575 -650 102609 -622
rect 102637 -650 102671 -622
rect 102699 -650 102747 -622
rect 102437 -684 102747 -650
rect 102437 -712 102485 -684
rect 102513 -712 102547 -684
rect 102575 -712 102609 -684
rect 102637 -712 102671 -684
rect 102699 -712 102747 -684
rect 102437 -746 102747 -712
rect 102437 -774 102485 -746
rect 102513 -774 102547 -746
rect 102575 -774 102609 -746
rect 102637 -774 102671 -746
rect 102699 -774 102747 -746
rect 102437 -822 102747 -774
rect 109577 47175 109887 49317
rect 109577 47147 109625 47175
rect 109653 47147 109687 47175
rect 109715 47147 109749 47175
rect 109777 47147 109811 47175
rect 109839 47147 109887 47175
rect 109577 47113 109887 47147
rect 109577 47085 109625 47113
rect 109653 47085 109687 47113
rect 109715 47085 109749 47113
rect 109777 47085 109811 47113
rect 109839 47085 109887 47113
rect 109577 47051 109887 47085
rect 109577 47023 109625 47051
rect 109653 47023 109687 47051
rect 109715 47023 109749 47051
rect 109777 47023 109811 47051
rect 109839 47023 109887 47051
rect 109577 46989 109887 47023
rect 109577 46961 109625 46989
rect 109653 46961 109687 46989
rect 109715 46961 109749 46989
rect 109777 46961 109811 46989
rect 109839 46961 109887 46989
rect 109577 38175 109887 46961
rect 109577 38147 109625 38175
rect 109653 38147 109687 38175
rect 109715 38147 109749 38175
rect 109777 38147 109811 38175
rect 109839 38147 109887 38175
rect 109577 38113 109887 38147
rect 109577 38085 109625 38113
rect 109653 38085 109687 38113
rect 109715 38085 109749 38113
rect 109777 38085 109811 38113
rect 109839 38085 109887 38113
rect 109577 38051 109887 38085
rect 109577 38023 109625 38051
rect 109653 38023 109687 38051
rect 109715 38023 109749 38051
rect 109777 38023 109811 38051
rect 109839 38023 109887 38051
rect 109577 37989 109887 38023
rect 109577 37961 109625 37989
rect 109653 37961 109687 37989
rect 109715 37961 109749 37989
rect 109777 37961 109811 37989
rect 109839 37961 109887 37989
rect 109577 29175 109887 37961
rect 109577 29147 109625 29175
rect 109653 29147 109687 29175
rect 109715 29147 109749 29175
rect 109777 29147 109811 29175
rect 109839 29147 109887 29175
rect 109577 29113 109887 29147
rect 109577 29085 109625 29113
rect 109653 29085 109687 29113
rect 109715 29085 109749 29113
rect 109777 29085 109811 29113
rect 109839 29085 109887 29113
rect 109577 29051 109887 29085
rect 109577 29023 109625 29051
rect 109653 29023 109687 29051
rect 109715 29023 109749 29051
rect 109777 29023 109811 29051
rect 109839 29023 109887 29051
rect 109577 28989 109887 29023
rect 109577 28961 109625 28989
rect 109653 28961 109687 28989
rect 109715 28961 109749 28989
rect 109777 28961 109811 28989
rect 109839 28961 109887 28989
rect 109577 20175 109887 28961
rect 109577 20147 109625 20175
rect 109653 20147 109687 20175
rect 109715 20147 109749 20175
rect 109777 20147 109811 20175
rect 109839 20147 109887 20175
rect 109577 20113 109887 20147
rect 109577 20085 109625 20113
rect 109653 20085 109687 20113
rect 109715 20085 109749 20113
rect 109777 20085 109811 20113
rect 109839 20085 109887 20113
rect 109577 20051 109887 20085
rect 109577 20023 109625 20051
rect 109653 20023 109687 20051
rect 109715 20023 109749 20051
rect 109777 20023 109811 20051
rect 109839 20023 109887 20051
rect 109577 19989 109887 20023
rect 109577 19961 109625 19989
rect 109653 19961 109687 19989
rect 109715 19961 109749 19989
rect 109777 19961 109811 19989
rect 109839 19961 109887 19989
rect 109577 11175 109887 19961
rect 109577 11147 109625 11175
rect 109653 11147 109687 11175
rect 109715 11147 109749 11175
rect 109777 11147 109811 11175
rect 109839 11147 109887 11175
rect 109577 11113 109887 11147
rect 109577 11085 109625 11113
rect 109653 11085 109687 11113
rect 109715 11085 109749 11113
rect 109777 11085 109811 11113
rect 109839 11085 109887 11113
rect 109577 11051 109887 11085
rect 109577 11023 109625 11051
rect 109653 11023 109687 11051
rect 109715 11023 109749 11051
rect 109777 11023 109811 11051
rect 109839 11023 109887 11051
rect 109577 10989 109887 11023
rect 109577 10961 109625 10989
rect 109653 10961 109687 10989
rect 109715 10961 109749 10989
rect 109777 10961 109811 10989
rect 109839 10961 109887 10989
rect 109577 2175 109887 10961
rect 109577 2147 109625 2175
rect 109653 2147 109687 2175
rect 109715 2147 109749 2175
rect 109777 2147 109811 2175
rect 109839 2147 109887 2175
rect 109577 2113 109887 2147
rect 109577 2085 109625 2113
rect 109653 2085 109687 2113
rect 109715 2085 109749 2113
rect 109777 2085 109811 2113
rect 109839 2085 109887 2113
rect 109577 2051 109887 2085
rect 109577 2023 109625 2051
rect 109653 2023 109687 2051
rect 109715 2023 109749 2051
rect 109777 2023 109811 2051
rect 109839 2023 109887 2051
rect 109577 1989 109887 2023
rect 109577 1961 109625 1989
rect 109653 1961 109687 1989
rect 109715 1961 109749 1989
rect 109777 1961 109811 1989
rect 109839 1961 109887 1989
rect 109577 -80 109887 1961
rect 109577 -108 109625 -80
rect 109653 -108 109687 -80
rect 109715 -108 109749 -80
rect 109777 -108 109811 -80
rect 109839 -108 109887 -80
rect 109577 -142 109887 -108
rect 109577 -170 109625 -142
rect 109653 -170 109687 -142
rect 109715 -170 109749 -142
rect 109777 -170 109811 -142
rect 109839 -170 109887 -142
rect 109577 -204 109887 -170
rect 109577 -232 109625 -204
rect 109653 -232 109687 -204
rect 109715 -232 109749 -204
rect 109777 -232 109811 -204
rect 109839 -232 109887 -204
rect 109577 -266 109887 -232
rect 109577 -294 109625 -266
rect 109653 -294 109687 -266
rect 109715 -294 109749 -266
rect 109777 -294 109811 -266
rect 109839 -294 109887 -266
rect 109577 -822 109887 -294
rect 111437 41175 111747 49317
rect 111437 41147 111485 41175
rect 111513 41147 111547 41175
rect 111575 41147 111609 41175
rect 111637 41147 111671 41175
rect 111699 41147 111747 41175
rect 111437 41113 111747 41147
rect 111437 41085 111485 41113
rect 111513 41085 111547 41113
rect 111575 41085 111609 41113
rect 111637 41085 111671 41113
rect 111699 41085 111747 41113
rect 111437 41051 111747 41085
rect 111437 41023 111485 41051
rect 111513 41023 111547 41051
rect 111575 41023 111609 41051
rect 111637 41023 111671 41051
rect 111699 41023 111747 41051
rect 111437 40989 111747 41023
rect 111437 40961 111485 40989
rect 111513 40961 111547 40989
rect 111575 40961 111609 40989
rect 111637 40961 111671 40989
rect 111699 40961 111747 40989
rect 111437 32175 111747 40961
rect 111437 32147 111485 32175
rect 111513 32147 111547 32175
rect 111575 32147 111609 32175
rect 111637 32147 111671 32175
rect 111699 32147 111747 32175
rect 111437 32113 111747 32147
rect 111437 32085 111485 32113
rect 111513 32085 111547 32113
rect 111575 32085 111609 32113
rect 111637 32085 111671 32113
rect 111699 32085 111747 32113
rect 111437 32051 111747 32085
rect 111437 32023 111485 32051
rect 111513 32023 111547 32051
rect 111575 32023 111609 32051
rect 111637 32023 111671 32051
rect 111699 32023 111747 32051
rect 111437 31989 111747 32023
rect 111437 31961 111485 31989
rect 111513 31961 111547 31989
rect 111575 31961 111609 31989
rect 111637 31961 111671 31989
rect 111699 31961 111747 31989
rect 111437 23175 111747 31961
rect 111437 23147 111485 23175
rect 111513 23147 111547 23175
rect 111575 23147 111609 23175
rect 111637 23147 111671 23175
rect 111699 23147 111747 23175
rect 111437 23113 111747 23147
rect 111437 23085 111485 23113
rect 111513 23085 111547 23113
rect 111575 23085 111609 23113
rect 111637 23085 111671 23113
rect 111699 23085 111747 23113
rect 111437 23051 111747 23085
rect 111437 23023 111485 23051
rect 111513 23023 111547 23051
rect 111575 23023 111609 23051
rect 111637 23023 111671 23051
rect 111699 23023 111747 23051
rect 111437 22989 111747 23023
rect 111437 22961 111485 22989
rect 111513 22961 111547 22989
rect 111575 22961 111609 22989
rect 111637 22961 111671 22989
rect 111699 22961 111747 22989
rect 111437 14175 111747 22961
rect 111437 14147 111485 14175
rect 111513 14147 111547 14175
rect 111575 14147 111609 14175
rect 111637 14147 111671 14175
rect 111699 14147 111747 14175
rect 111437 14113 111747 14147
rect 111437 14085 111485 14113
rect 111513 14085 111547 14113
rect 111575 14085 111609 14113
rect 111637 14085 111671 14113
rect 111699 14085 111747 14113
rect 111437 14051 111747 14085
rect 111437 14023 111485 14051
rect 111513 14023 111547 14051
rect 111575 14023 111609 14051
rect 111637 14023 111671 14051
rect 111699 14023 111747 14051
rect 111437 13989 111747 14023
rect 111437 13961 111485 13989
rect 111513 13961 111547 13989
rect 111575 13961 111609 13989
rect 111637 13961 111671 13989
rect 111699 13961 111747 13989
rect 111437 5175 111747 13961
rect 111437 5147 111485 5175
rect 111513 5147 111547 5175
rect 111575 5147 111609 5175
rect 111637 5147 111671 5175
rect 111699 5147 111747 5175
rect 111437 5113 111747 5147
rect 111437 5085 111485 5113
rect 111513 5085 111547 5113
rect 111575 5085 111609 5113
rect 111637 5085 111671 5113
rect 111699 5085 111747 5113
rect 111437 5051 111747 5085
rect 111437 5023 111485 5051
rect 111513 5023 111547 5051
rect 111575 5023 111609 5051
rect 111637 5023 111671 5051
rect 111699 5023 111747 5051
rect 111437 4989 111747 5023
rect 111437 4961 111485 4989
rect 111513 4961 111547 4989
rect 111575 4961 111609 4989
rect 111637 4961 111671 4989
rect 111699 4961 111747 4989
rect 111437 -560 111747 4961
rect 111437 -588 111485 -560
rect 111513 -588 111547 -560
rect 111575 -588 111609 -560
rect 111637 -588 111671 -560
rect 111699 -588 111747 -560
rect 111437 -622 111747 -588
rect 111437 -650 111485 -622
rect 111513 -650 111547 -622
rect 111575 -650 111609 -622
rect 111637 -650 111671 -622
rect 111699 -650 111747 -622
rect 111437 -684 111747 -650
rect 111437 -712 111485 -684
rect 111513 -712 111547 -684
rect 111575 -712 111609 -684
rect 111637 -712 111671 -684
rect 111699 -712 111747 -684
rect 111437 -746 111747 -712
rect 111437 -774 111485 -746
rect 111513 -774 111547 -746
rect 111575 -774 111609 -746
rect 111637 -774 111671 -746
rect 111699 -774 111747 -746
rect 111437 -822 111747 -774
rect 118577 47175 118887 49317
rect 118577 47147 118625 47175
rect 118653 47147 118687 47175
rect 118715 47147 118749 47175
rect 118777 47147 118811 47175
rect 118839 47147 118887 47175
rect 118577 47113 118887 47147
rect 118577 47085 118625 47113
rect 118653 47085 118687 47113
rect 118715 47085 118749 47113
rect 118777 47085 118811 47113
rect 118839 47085 118887 47113
rect 118577 47051 118887 47085
rect 118577 47023 118625 47051
rect 118653 47023 118687 47051
rect 118715 47023 118749 47051
rect 118777 47023 118811 47051
rect 118839 47023 118887 47051
rect 118577 46989 118887 47023
rect 118577 46961 118625 46989
rect 118653 46961 118687 46989
rect 118715 46961 118749 46989
rect 118777 46961 118811 46989
rect 118839 46961 118887 46989
rect 118577 38175 118887 46961
rect 118577 38147 118625 38175
rect 118653 38147 118687 38175
rect 118715 38147 118749 38175
rect 118777 38147 118811 38175
rect 118839 38147 118887 38175
rect 118577 38113 118887 38147
rect 118577 38085 118625 38113
rect 118653 38085 118687 38113
rect 118715 38085 118749 38113
rect 118777 38085 118811 38113
rect 118839 38085 118887 38113
rect 118577 38051 118887 38085
rect 118577 38023 118625 38051
rect 118653 38023 118687 38051
rect 118715 38023 118749 38051
rect 118777 38023 118811 38051
rect 118839 38023 118887 38051
rect 118577 37989 118887 38023
rect 118577 37961 118625 37989
rect 118653 37961 118687 37989
rect 118715 37961 118749 37989
rect 118777 37961 118811 37989
rect 118839 37961 118887 37989
rect 118577 29175 118887 37961
rect 118577 29147 118625 29175
rect 118653 29147 118687 29175
rect 118715 29147 118749 29175
rect 118777 29147 118811 29175
rect 118839 29147 118887 29175
rect 118577 29113 118887 29147
rect 118577 29085 118625 29113
rect 118653 29085 118687 29113
rect 118715 29085 118749 29113
rect 118777 29085 118811 29113
rect 118839 29085 118887 29113
rect 118577 29051 118887 29085
rect 118577 29023 118625 29051
rect 118653 29023 118687 29051
rect 118715 29023 118749 29051
rect 118777 29023 118811 29051
rect 118839 29023 118887 29051
rect 118577 28989 118887 29023
rect 118577 28961 118625 28989
rect 118653 28961 118687 28989
rect 118715 28961 118749 28989
rect 118777 28961 118811 28989
rect 118839 28961 118887 28989
rect 118577 20175 118887 28961
rect 118577 20147 118625 20175
rect 118653 20147 118687 20175
rect 118715 20147 118749 20175
rect 118777 20147 118811 20175
rect 118839 20147 118887 20175
rect 118577 20113 118887 20147
rect 118577 20085 118625 20113
rect 118653 20085 118687 20113
rect 118715 20085 118749 20113
rect 118777 20085 118811 20113
rect 118839 20085 118887 20113
rect 118577 20051 118887 20085
rect 118577 20023 118625 20051
rect 118653 20023 118687 20051
rect 118715 20023 118749 20051
rect 118777 20023 118811 20051
rect 118839 20023 118887 20051
rect 118577 19989 118887 20023
rect 118577 19961 118625 19989
rect 118653 19961 118687 19989
rect 118715 19961 118749 19989
rect 118777 19961 118811 19989
rect 118839 19961 118887 19989
rect 118577 11175 118887 19961
rect 118577 11147 118625 11175
rect 118653 11147 118687 11175
rect 118715 11147 118749 11175
rect 118777 11147 118811 11175
rect 118839 11147 118887 11175
rect 118577 11113 118887 11147
rect 118577 11085 118625 11113
rect 118653 11085 118687 11113
rect 118715 11085 118749 11113
rect 118777 11085 118811 11113
rect 118839 11085 118887 11113
rect 118577 11051 118887 11085
rect 118577 11023 118625 11051
rect 118653 11023 118687 11051
rect 118715 11023 118749 11051
rect 118777 11023 118811 11051
rect 118839 11023 118887 11051
rect 118577 10989 118887 11023
rect 118577 10961 118625 10989
rect 118653 10961 118687 10989
rect 118715 10961 118749 10989
rect 118777 10961 118811 10989
rect 118839 10961 118887 10989
rect 118577 2175 118887 10961
rect 118577 2147 118625 2175
rect 118653 2147 118687 2175
rect 118715 2147 118749 2175
rect 118777 2147 118811 2175
rect 118839 2147 118887 2175
rect 118577 2113 118887 2147
rect 118577 2085 118625 2113
rect 118653 2085 118687 2113
rect 118715 2085 118749 2113
rect 118777 2085 118811 2113
rect 118839 2085 118887 2113
rect 118577 2051 118887 2085
rect 118577 2023 118625 2051
rect 118653 2023 118687 2051
rect 118715 2023 118749 2051
rect 118777 2023 118811 2051
rect 118839 2023 118887 2051
rect 118577 1989 118887 2023
rect 118577 1961 118625 1989
rect 118653 1961 118687 1989
rect 118715 1961 118749 1989
rect 118777 1961 118811 1989
rect 118839 1961 118887 1989
rect 118577 -80 118887 1961
rect 118577 -108 118625 -80
rect 118653 -108 118687 -80
rect 118715 -108 118749 -80
rect 118777 -108 118811 -80
rect 118839 -108 118887 -80
rect 118577 -142 118887 -108
rect 118577 -170 118625 -142
rect 118653 -170 118687 -142
rect 118715 -170 118749 -142
rect 118777 -170 118811 -142
rect 118839 -170 118887 -142
rect 118577 -204 118887 -170
rect 118577 -232 118625 -204
rect 118653 -232 118687 -204
rect 118715 -232 118749 -204
rect 118777 -232 118811 -204
rect 118839 -232 118887 -204
rect 118577 -266 118887 -232
rect 118577 -294 118625 -266
rect 118653 -294 118687 -266
rect 118715 -294 118749 -266
rect 118777 -294 118811 -266
rect 118839 -294 118887 -266
rect 118577 -822 118887 -294
rect 120437 41175 120747 49961
rect 120437 41147 120485 41175
rect 120513 41147 120547 41175
rect 120575 41147 120609 41175
rect 120637 41147 120671 41175
rect 120699 41147 120747 41175
rect 120437 41113 120747 41147
rect 120437 41085 120485 41113
rect 120513 41085 120547 41113
rect 120575 41085 120609 41113
rect 120637 41085 120671 41113
rect 120699 41085 120747 41113
rect 120437 41051 120747 41085
rect 120437 41023 120485 41051
rect 120513 41023 120547 41051
rect 120575 41023 120609 41051
rect 120637 41023 120671 41051
rect 120699 41023 120747 41051
rect 120437 40989 120747 41023
rect 120437 40961 120485 40989
rect 120513 40961 120547 40989
rect 120575 40961 120609 40989
rect 120637 40961 120671 40989
rect 120699 40961 120747 40989
rect 120437 32175 120747 40961
rect 120437 32147 120485 32175
rect 120513 32147 120547 32175
rect 120575 32147 120609 32175
rect 120637 32147 120671 32175
rect 120699 32147 120747 32175
rect 120437 32113 120747 32147
rect 120437 32085 120485 32113
rect 120513 32085 120547 32113
rect 120575 32085 120609 32113
rect 120637 32085 120671 32113
rect 120699 32085 120747 32113
rect 120437 32051 120747 32085
rect 120437 32023 120485 32051
rect 120513 32023 120547 32051
rect 120575 32023 120609 32051
rect 120637 32023 120671 32051
rect 120699 32023 120747 32051
rect 120437 31989 120747 32023
rect 120437 31961 120485 31989
rect 120513 31961 120547 31989
rect 120575 31961 120609 31989
rect 120637 31961 120671 31989
rect 120699 31961 120747 31989
rect 120437 23175 120747 31961
rect 120437 23147 120485 23175
rect 120513 23147 120547 23175
rect 120575 23147 120609 23175
rect 120637 23147 120671 23175
rect 120699 23147 120747 23175
rect 120437 23113 120747 23147
rect 120437 23085 120485 23113
rect 120513 23085 120547 23113
rect 120575 23085 120609 23113
rect 120637 23085 120671 23113
rect 120699 23085 120747 23113
rect 120437 23051 120747 23085
rect 120437 23023 120485 23051
rect 120513 23023 120547 23051
rect 120575 23023 120609 23051
rect 120637 23023 120671 23051
rect 120699 23023 120747 23051
rect 120437 22989 120747 23023
rect 120437 22961 120485 22989
rect 120513 22961 120547 22989
rect 120575 22961 120609 22989
rect 120637 22961 120671 22989
rect 120699 22961 120747 22989
rect 120437 14175 120747 22961
rect 120437 14147 120485 14175
rect 120513 14147 120547 14175
rect 120575 14147 120609 14175
rect 120637 14147 120671 14175
rect 120699 14147 120747 14175
rect 120437 14113 120747 14147
rect 120437 14085 120485 14113
rect 120513 14085 120547 14113
rect 120575 14085 120609 14113
rect 120637 14085 120671 14113
rect 120699 14085 120747 14113
rect 120437 14051 120747 14085
rect 120437 14023 120485 14051
rect 120513 14023 120547 14051
rect 120575 14023 120609 14051
rect 120637 14023 120671 14051
rect 120699 14023 120747 14051
rect 120437 13989 120747 14023
rect 120437 13961 120485 13989
rect 120513 13961 120547 13989
rect 120575 13961 120609 13989
rect 120637 13961 120671 13989
rect 120699 13961 120747 13989
rect 120437 5175 120747 13961
rect 120437 5147 120485 5175
rect 120513 5147 120547 5175
rect 120575 5147 120609 5175
rect 120637 5147 120671 5175
rect 120699 5147 120747 5175
rect 120437 5113 120747 5147
rect 120437 5085 120485 5113
rect 120513 5085 120547 5113
rect 120575 5085 120609 5113
rect 120637 5085 120671 5113
rect 120699 5085 120747 5113
rect 120437 5051 120747 5085
rect 120437 5023 120485 5051
rect 120513 5023 120547 5051
rect 120575 5023 120609 5051
rect 120637 5023 120671 5051
rect 120699 5023 120747 5051
rect 120437 4989 120747 5023
rect 120437 4961 120485 4989
rect 120513 4961 120547 4989
rect 120575 4961 120609 4989
rect 120637 4961 120671 4989
rect 120699 4961 120747 4989
rect 120437 -560 120747 4961
rect 120437 -588 120485 -560
rect 120513 -588 120547 -560
rect 120575 -588 120609 -560
rect 120637 -588 120671 -560
rect 120699 -588 120747 -560
rect 120437 -622 120747 -588
rect 120437 -650 120485 -622
rect 120513 -650 120547 -622
rect 120575 -650 120609 -622
rect 120637 -650 120671 -622
rect 120699 -650 120747 -622
rect 120437 -684 120747 -650
rect 120437 -712 120485 -684
rect 120513 -712 120547 -684
rect 120575 -712 120609 -684
rect 120637 -712 120671 -684
rect 120699 -712 120747 -684
rect 120437 -746 120747 -712
rect 120437 -774 120485 -746
rect 120513 -774 120547 -746
rect 120575 -774 120609 -746
rect 120637 -774 120671 -746
rect 120699 -774 120747 -746
rect 120437 -822 120747 -774
rect 127577 119175 127887 124261
rect 127577 119147 127625 119175
rect 127653 119147 127687 119175
rect 127715 119147 127749 119175
rect 127777 119147 127811 119175
rect 127839 119147 127887 119175
rect 127577 119113 127887 119147
rect 127577 119085 127625 119113
rect 127653 119085 127687 119113
rect 127715 119085 127749 119113
rect 127777 119085 127811 119113
rect 127839 119085 127887 119113
rect 127577 119051 127887 119085
rect 127577 119023 127625 119051
rect 127653 119023 127687 119051
rect 127715 119023 127749 119051
rect 127777 119023 127811 119051
rect 127839 119023 127887 119051
rect 127577 118989 127887 119023
rect 127577 118961 127625 118989
rect 127653 118961 127687 118989
rect 127715 118961 127749 118989
rect 127777 118961 127811 118989
rect 127839 118961 127887 118989
rect 127577 110175 127887 118961
rect 127577 110147 127625 110175
rect 127653 110147 127687 110175
rect 127715 110147 127749 110175
rect 127777 110147 127811 110175
rect 127839 110147 127887 110175
rect 127577 110113 127887 110147
rect 127577 110085 127625 110113
rect 127653 110085 127687 110113
rect 127715 110085 127749 110113
rect 127777 110085 127811 110113
rect 127839 110085 127887 110113
rect 127577 110051 127887 110085
rect 127577 110023 127625 110051
rect 127653 110023 127687 110051
rect 127715 110023 127749 110051
rect 127777 110023 127811 110051
rect 127839 110023 127887 110051
rect 127577 109989 127887 110023
rect 127577 109961 127625 109989
rect 127653 109961 127687 109989
rect 127715 109961 127749 109989
rect 127777 109961 127811 109989
rect 127839 109961 127887 109989
rect 127577 101175 127887 109961
rect 127577 101147 127625 101175
rect 127653 101147 127687 101175
rect 127715 101147 127749 101175
rect 127777 101147 127811 101175
rect 127839 101147 127887 101175
rect 127577 101113 127887 101147
rect 127577 101085 127625 101113
rect 127653 101085 127687 101113
rect 127715 101085 127749 101113
rect 127777 101085 127811 101113
rect 127839 101085 127887 101113
rect 127577 101051 127887 101085
rect 127577 101023 127625 101051
rect 127653 101023 127687 101051
rect 127715 101023 127749 101051
rect 127777 101023 127811 101051
rect 127839 101023 127887 101051
rect 127577 100989 127887 101023
rect 127577 100961 127625 100989
rect 127653 100961 127687 100989
rect 127715 100961 127749 100989
rect 127777 100961 127811 100989
rect 127839 100961 127887 100989
rect 127577 92175 127887 100961
rect 127577 92147 127625 92175
rect 127653 92147 127687 92175
rect 127715 92147 127749 92175
rect 127777 92147 127811 92175
rect 127839 92147 127887 92175
rect 127577 92113 127887 92147
rect 127577 92085 127625 92113
rect 127653 92085 127687 92113
rect 127715 92085 127749 92113
rect 127777 92085 127811 92113
rect 127839 92085 127887 92113
rect 127577 92051 127887 92085
rect 127577 92023 127625 92051
rect 127653 92023 127687 92051
rect 127715 92023 127749 92051
rect 127777 92023 127811 92051
rect 127839 92023 127887 92051
rect 127577 91989 127887 92023
rect 127577 91961 127625 91989
rect 127653 91961 127687 91989
rect 127715 91961 127749 91989
rect 127777 91961 127811 91989
rect 127839 91961 127887 91989
rect 127577 83175 127887 91961
rect 127577 83147 127625 83175
rect 127653 83147 127687 83175
rect 127715 83147 127749 83175
rect 127777 83147 127811 83175
rect 127839 83147 127887 83175
rect 127577 83113 127887 83147
rect 127577 83085 127625 83113
rect 127653 83085 127687 83113
rect 127715 83085 127749 83113
rect 127777 83085 127811 83113
rect 127839 83085 127887 83113
rect 127577 83051 127887 83085
rect 127577 83023 127625 83051
rect 127653 83023 127687 83051
rect 127715 83023 127749 83051
rect 127777 83023 127811 83051
rect 127839 83023 127887 83051
rect 127577 82989 127887 83023
rect 127577 82961 127625 82989
rect 127653 82961 127687 82989
rect 127715 82961 127749 82989
rect 127777 82961 127811 82989
rect 127839 82961 127887 82989
rect 127577 74175 127887 82961
rect 127577 74147 127625 74175
rect 127653 74147 127687 74175
rect 127715 74147 127749 74175
rect 127777 74147 127811 74175
rect 127839 74147 127887 74175
rect 127577 74113 127887 74147
rect 127577 74085 127625 74113
rect 127653 74085 127687 74113
rect 127715 74085 127749 74113
rect 127777 74085 127811 74113
rect 127839 74085 127887 74113
rect 127577 74051 127887 74085
rect 127577 74023 127625 74051
rect 127653 74023 127687 74051
rect 127715 74023 127749 74051
rect 127777 74023 127811 74051
rect 127839 74023 127887 74051
rect 127577 73989 127887 74023
rect 127577 73961 127625 73989
rect 127653 73961 127687 73989
rect 127715 73961 127749 73989
rect 127777 73961 127811 73989
rect 127839 73961 127887 73989
rect 127577 65175 127887 73961
rect 127577 65147 127625 65175
rect 127653 65147 127687 65175
rect 127715 65147 127749 65175
rect 127777 65147 127811 65175
rect 127839 65147 127887 65175
rect 127577 65113 127887 65147
rect 127577 65085 127625 65113
rect 127653 65085 127687 65113
rect 127715 65085 127749 65113
rect 127777 65085 127811 65113
rect 127839 65085 127887 65113
rect 127577 65051 127887 65085
rect 127577 65023 127625 65051
rect 127653 65023 127687 65051
rect 127715 65023 127749 65051
rect 127777 65023 127811 65051
rect 127839 65023 127887 65051
rect 127577 64989 127887 65023
rect 127577 64961 127625 64989
rect 127653 64961 127687 64989
rect 127715 64961 127749 64989
rect 127777 64961 127811 64989
rect 127839 64961 127887 64989
rect 127577 56175 127887 64961
rect 127577 56147 127625 56175
rect 127653 56147 127687 56175
rect 127715 56147 127749 56175
rect 127777 56147 127811 56175
rect 127839 56147 127887 56175
rect 127577 56113 127887 56147
rect 127577 56085 127625 56113
rect 127653 56085 127687 56113
rect 127715 56085 127749 56113
rect 127777 56085 127811 56113
rect 127839 56085 127887 56113
rect 127577 56051 127887 56085
rect 127577 56023 127625 56051
rect 127653 56023 127687 56051
rect 127715 56023 127749 56051
rect 127777 56023 127811 56051
rect 127839 56023 127887 56051
rect 127577 55989 127887 56023
rect 127577 55961 127625 55989
rect 127653 55961 127687 55989
rect 127715 55961 127749 55989
rect 127777 55961 127811 55989
rect 127839 55961 127887 55989
rect 127577 47175 127887 55961
rect 127577 47147 127625 47175
rect 127653 47147 127687 47175
rect 127715 47147 127749 47175
rect 127777 47147 127811 47175
rect 127839 47147 127887 47175
rect 127577 47113 127887 47147
rect 127577 47085 127625 47113
rect 127653 47085 127687 47113
rect 127715 47085 127749 47113
rect 127777 47085 127811 47113
rect 127839 47085 127887 47113
rect 127577 47051 127887 47085
rect 127577 47023 127625 47051
rect 127653 47023 127687 47051
rect 127715 47023 127749 47051
rect 127777 47023 127811 47051
rect 127839 47023 127887 47051
rect 127577 46989 127887 47023
rect 127577 46961 127625 46989
rect 127653 46961 127687 46989
rect 127715 46961 127749 46989
rect 127777 46961 127811 46989
rect 127839 46961 127887 46989
rect 127577 38175 127887 46961
rect 127577 38147 127625 38175
rect 127653 38147 127687 38175
rect 127715 38147 127749 38175
rect 127777 38147 127811 38175
rect 127839 38147 127887 38175
rect 127577 38113 127887 38147
rect 127577 38085 127625 38113
rect 127653 38085 127687 38113
rect 127715 38085 127749 38113
rect 127777 38085 127811 38113
rect 127839 38085 127887 38113
rect 127577 38051 127887 38085
rect 127577 38023 127625 38051
rect 127653 38023 127687 38051
rect 127715 38023 127749 38051
rect 127777 38023 127811 38051
rect 127839 38023 127887 38051
rect 127577 37989 127887 38023
rect 127577 37961 127625 37989
rect 127653 37961 127687 37989
rect 127715 37961 127749 37989
rect 127777 37961 127811 37989
rect 127839 37961 127887 37989
rect 127577 29175 127887 37961
rect 127577 29147 127625 29175
rect 127653 29147 127687 29175
rect 127715 29147 127749 29175
rect 127777 29147 127811 29175
rect 127839 29147 127887 29175
rect 127577 29113 127887 29147
rect 127577 29085 127625 29113
rect 127653 29085 127687 29113
rect 127715 29085 127749 29113
rect 127777 29085 127811 29113
rect 127839 29085 127887 29113
rect 127577 29051 127887 29085
rect 127577 29023 127625 29051
rect 127653 29023 127687 29051
rect 127715 29023 127749 29051
rect 127777 29023 127811 29051
rect 127839 29023 127887 29051
rect 127577 28989 127887 29023
rect 127577 28961 127625 28989
rect 127653 28961 127687 28989
rect 127715 28961 127749 28989
rect 127777 28961 127811 28989
rect 127839 28961 127887 28989
rect 127577 20175 127887 28961
rect 127577 20147 127625 20175
rect 127653 20147 127687 20175
rect 127715 20147 127749 20175
rect 127777 20147 127811 20175
rect 127839 20147 127887 20175
rect 127577 20113 127887 20147
rect 127577 20085 127625 20113
rect 127653 20085 127687 20113
rect 127715 20085 127749 20113
rect 127777 20085 127811 20113
rect 127839 20085 127887 20113
rect 127577 20051 127887 20085
rect 127577 20023 127625 20051
rect 127653 20023 127687 20051
rect 127715 20023 127749 20051
rect 127777 20023 127811 20051
rect 127839 20023 127887 20051
rect 127577 19989 127887 20023
rect 127577 19961 127625 19989
rect 127653 19961 127687 19989
rect 127715 19961 127749 19989
rect 127777 19961 127811 19989
rect 127839 19961 127887 19989
rect 127577 11175 127887 19961
rect 127577 11147 127625 11175
rect 127653 11147 127687 11175
rect 127715 11147 127749 11175
rect 127777 11147 127811 11175
rect 127839 11147 127887 11175
rect 127577 11113 127887 11147
rect 127577 11085 127625 11113
rect 127653 11085 127687 11113
rect 127715 11085 127749 11113
rect 127777 11085 127811 11113
rect 127839 11085 127887 11113
rect 127577 11051 127887 11085
rect 127577 11023 127625 11051
rect 127653 11023 127687 11051
rect 127715 11023 127749 11051
rect 127777 11023 127811 11051
rect 127839 11023 127887 11051
rect 127577 10989 127887 11023
rect 127577 10961 127625 10989
rect 127653 10961 127687 10989
rect 127715 10961 127749 10989
rect 127777 10961 127811 10989
rect 127839 10961 127887 10989
rect 127577 2175 127887 10961
rect 127577 2147 127625 2175
rect 127653 2147 127687 2175
rect 127715 2147 127749 2175
rect 127777 2147 127811 2175
rect 127839 2147 127887 2175
rect 127577 2113 127887 2147
rect 127577 2085 127625 2113
rect 127653 2085 127687 2113
rect 127715 2085 127749 2113
rect 127777 2085 127811 2113
rect 127839 2085 127887 2113
rect 127577 2051 127887 2085
rect 127577 2023 127625 2051
rect 127653 2023 127687 2051
rect 127715 2023 127749 2051
rect 127777 2023 127811 2051
rect 127839 2023 127887 2051
rect 127577 1989 127887 2023
rect 127577 1961 127625 1989
rect 127653 1961 127687 1989
rect 127715 1961 127749 1989
rect 127777 1961 127811 1989
rect 127839 1961 127887 1989
rect 127577 -80 127887 1961
rect 127577 -108 127625 -80
rect 127653 -108 127687 -80
rect 127715 -108 127749 -80
rect 127777 -108 127811 -80
rect 127839 -108 127887 -80
rect 127577 -142 127887 -108
rect 127577 -170 127625 -142
rect 127653 -170 127687 -142
rect 127715 -170 127749 -142
rect 127777 -170 127811 -142
rect 127839 -170 127887 -142
rect 127577 -204 127887 -170
rect 127577 -232 127625 -204
rect 127653 -232 127687 -204
rect 127715 -232 127749 -204
rect 127777 -232 127811 -204
rect 127839 -232 127887 -204
rect 127577 -266 127887 -232
rect 127577 -294 127625 -266
rect 127653 -294 127687 -266
rect 127715 -294 127749 -266
rect 127777 -294 127811 -266
rect 127839 -294 127887 -266
rect 127577 -822 127887 -294
rect 129437 122175 129747 124261
rect 129437 122147 129485 122175
rect 129513 122147 129547 122175
rect 129575 122147 129609 122175
rect 129637 122147 129671 122175
rect 129699 122147 129747 122175
rect 129437 122113 129747 122147
rect 129437 122085 129485 122113
rect 129513 122085 129547 122113
rect 129575 122085 129609 122113
rect 129637 122085 129671 122113
rect 129699 122085 129747 122113
rect 129437 122051 129747 122085
rect 129437 122023 129485 122051
rect 129513 122023 129547 122051
rect 129575 122023 129609 122051
rect 129637 122023 129671 122051
rect 129699 122023 129747 122051
rect 129437 121989 129747 122023
rect 129437 121961 129485 121989
rect 129513 121961 129547 121989
rect 129575 121961 129609 121989
rect 129637 121961 129671 121989
rect 129699 121961 129747 121989
rect 129437 113175 129747 121961
rect 129437 113147 129485 113175
rect 129513 113147 129547 113175
rect 129575 113147 129609 113175
rect 129637 113147 129671 113175
rect 129699 113147 129747 113175
rect 129437 113113 129747 113147
rect 129437 113085 129485 113113
rect 129513 113085 129547 113113
rect 129575 113085 129609 113113
rect 129637 113085 129671 113113
rect 129699 113085 129747 113113
rect 129437 113051 129747 113085
rect 129437 113023 129485 113051
rect 129513 113023 129547 113051
rect 129575 113023 129609 113051
rect 129637 113023 129671 113051
rect 129699 113023 129747 113051
rect 129437 112989 129747 113023
rect 129437 112961 129485 112989
rect 129513 112961 129547 112989
rect 129575 112961 129609 112989
rect 129637 112961 129671 112989
rect 129699 112961 129747 112989
rect 129437 104175 129747 112961
rect 129437 104147 129485 104175
rect 129513 104147 129547 104175
rect 129575 104147 129609 104175
rect 129637 104147 129671 104175
rect 129699 104147 129747 104175
rect 129437 104113 129747 104147
rect 129437 104085 129485 104113
rect 129513 104085 129547 104113
rect 129575 104085 129609 104113
rect 129637 104085 129671 104113
rect 129699 104085 129747 104113
rect 129437 104051 129747 104085
rect 129437 104023 129485 104051
rect 129513 104023 129547 104051
rect 129575 104023 129609 104051
rect 129637 104023 129671 104051
rect 129699 104023 129747 104051
rect 129437 103989 129747 104023
rect 129437 103961 129485 103989
rect 129513 103961 129547 103989
rect 129575 103961 129609 103989
rect 129637 103961 129671 103989
rect 129699 103961 129747 103989
rect 129437 95175 129747 103961
rect 129437 95147 129485 95175
rect 129513 95147 129547 95175
rect 129575 95147 129609 95175
rect 129637 95147 129671 95175
rect 129699 95147 129747 95175
rect 129437 95113 129747 95147
rect 129437 95085 129485 95113
rect 129513 95085 129547 95113
rect 129575 95085 129609 95113
rect 129637 95085 129671 95113
rect 129699 95085 129747 95113
rect 129437 95051 129747 95085
rect 129437 95023 129485 95051
rect 129513 95023 129547 95051
rect 129575 95023 129609 95051
rect 129637 95023 129671 95051
rect 129699 95023 129747 95051
rect 129437 94989 129747 95023
rect 129437 94961 129485 94989
rect 129513 94961 129547 94989
rect 129575 94961 129609 94989
rect 129637 94961 129671 94989
rect 129699 94961 129747 94989
rect 129437 86175 129747 94961
rect 129437 86147 129485 86175
rect 129513 86147 129547 86175
rect 129575 86147 129609 86175
rect 129637 86147 129671 86175
rect 129699 86147 129747 86175
rect 129437 86113 129747 86147
rect 129437 86085 129485 86113
rect 129513 86085 129547 86113
rect 129575 86085 129609 86113
rect 129637 86085 129671 86113
rect 129699 86085 129747 86113
rect 129437 86051 129747 86085
rect 129437 86023 129485 86051
rect 129513 86023 129547 86051
rect 129575 86023 129609 86051
rect 129637 86023 129671 86051
rect 129699 86023 129747 86051
rect 129437 85989 129747 86023
rect 129437 85961 129485 85989
rect 129513 85961 129547 85989
rect 129575 85961 129609 85989
rect 129637 85961 129671 85989
rect 129699 85961 129747 85989
rect 129437 77175 129747 85961
rect 129437 77147 129485 77175
rect 129513 77147 129547 77175
rect 129575 77147 129609 77175
rect 129637 77147 129671 77175
rect 129699 77147 129747 77175
rect 129437 77113 129747 77147
rect 129437 77085 129485 77113
rect 129513 77085 129547 77113
rect 129575 77085 129609 77113
rect 129637 77085 129671 77113
rect 129699 77085 129747 77113
rect 129437 77051 129747 77085
rect 129437 77023 129485 77051
rect 129513 77023 129547 77051
rect 129575 77023 129609 77051
rect 129637 77023 129671 77051
rect 129699 77023 129747 77051
rect 129437 76989 129747 77023
rect 129437 76961 129485 76989
rect 129513 76961 129547 76989
rect 129575 76961 129609 76989
rect 129637 76961 129671 76989
rect 129699 76961 129747 76989
rect 129437 68175 129747 76961
rect 129437 68147 129485 68175
rect 129513 68147 129547 68175
rect 129575 68147 129609 68175
rect 129637 68147 129671 68175
rect 129699 68147 129747 68175
rect 129437 68113 129747 68147
rect 129437 68085 129485 68113
rect 129513 68085 129547 68113
rect 129575 68085 129609 68113
rect 129637 68085 129671 68113
rect 129699 68085 129747 68113
rect 129437 68051 129747 68085
rect 129437 68023 129485 68051
rect 129513 68023 129547 68051
rect 129575 68023 129609 68051
rect 129637 68023 129671 68051
rect 129699 68023 129747 68051
rect 129437 67989 129747 68023
rect 129437 67961 129485 67989
rect 129513 67961 129547 67989
rect 129575 67961 129609 67989
rect 129637 67961 129671 67989
rect 129699 67961 129747 67989
rect 129437 59175 129747 67961
rect 129437 59147 129485 59175
rect 129513 59147 129547 59175
rect 129575 59147 129609 59175
rect 129637 59147 129671 59175
rect 129699 59147 129747 59175
rect 129437 59113 129747 59147
rect 129437 59085 129485 59113
rect 129513 59085 129547 59113
rect 129575 59085 129609 59113
rect 129637 59085 129671 59113
rect 129699 59085 129747 59113
rect 129437 59051 129747 59085
rect 129437 59023 129485 59051
rect 129513 59023 129547 59051
rect 129575 59023 129609 59051
rect 129637 59023 129671 59051
rect 129699 59023 129747 59051
rect 129437 58989 129747 59023
rect 129437 58961 129485 58989
rect 129513 58961 129547 58989
rect 129575 58961 129609 58989
rect 129637 58961 129671 58989
rect 129699 58961 129747 58989
rect 129437 50175 129747 58961
rect 129437 50147 129485 50175
rect 129513 50147 129547 50175
rect 129575 50147 129609 50175
rect 129637 50147 129671 50175
rect 129699 50147 129747 50175
rect 129437 50113 129747 50147
rect 129437 50085 129485 50113
rect 129513 50085 129547 50113
rect 129575 50085 129609 50113
rect 129637 50085 129671 50113
rect 129699 50085 129747 50113
rect 129437 50051 129747 50085
rect 129437 50023 129485 50051
rect 129513 50023 129547 50051
rect 129575 50023 129609 50051
rect 129637 50023 129671 50051
rect 129699 50023 129747 50051
rect 129437 49989 129747 50023
rect 129437 49961 129485 49989
rect 129513 49961 129547 49989
rect 129575 49961 129609 49989
rect 129637 49961 129671 49989
rect 129699 49961 129747 49989
rect 129437 41175 129747 49961
rect 129437 41147 129485 41175
rect 129513 41147 129547 41175
rect 129575 41147 129609 41175
rect 129637 41147 129671 41175
rect 129699 41147 129747 41175
rect 129437 41113 129747 41147
rect 129437 41085 129485 41113
rect 129513 41085 129547 41113
rect 129575 41085 129609 41113
rect 129637 41085 129671 41113
rect 129699 41085 129747 41113
rect 129437 41051 129747 41085
rect 129437 41023 129485 41051
rect 129513 41023 129547 41051
rect 129575 41023 129609 41051
rect 129637 41023 129671 41051
rect 129699 41023 129747 41051
rect 129437 40989 129747 41023
rect 129437 40961 129485 40989
rect 129513 40961 129547 40989
rect 129575 40961 129609 40989
rect 129637 40961 129671 40989
rect 129699 40961 129747 40989
rect 129437 32175 129747 40961
rect 129437 32147 129485 32175
rect 129513 32147 129547 32175
rect 129575 32147 129609 32175
rect 129637 32147 129671 32175
rect 129699 32147 129747 32175
rect 129437 32113 129747 32147
rect 129437 32085 129485 32113
rect 129513 32085 129547 32113
rect 129575 32085 129609 32113
rect 129637 32085 129671 32113
rect 129699 32085 129747 32113
rect 129437 32051 129747 32085
rect 129437 32023 129485 32051
rect 129513 32023 129547 32051
rect 129575 32023 129609 32051
rect 129637 32023 129671 32051
rect 129699 32023 129747 32051
rect 129437 31989 129747 32023
rect 129437 31961 129485 31989
rect 129513 31961 129547 31989
rect 129575 31961 129609 31989
rect 129637 31961 129671 31989
rect 129699 31961 129747 31989
rect 129437 23175 129747 31961
rect 129437 23147 129485 23175
rect 129513 23147 129547 23175
rect 129575 23147 129609 23175
rect 129637 23147 129671 23175
rect 129699 23147 129747 23175
rect 129437 23113 129747 23147
rect 129437 23085 129485 23113
rect 129513 23085 129547 23113
rect 129575 23085 129609 23113
rect 129637 23085 129671 23113
rect 129699 23085 129747 23113
rect 129437 23051 129747 23085
rect 129437 23023 129485 23051
rect 129513 23023 129547 23051
rect 129575 23023 129609 23051
rect 129637 23023 129671 23051
rect 129699 23023 129747 23051
rect 129437 22989 129747 23023
rect 129437 22961 129485 22989
rect 129513 22961 129547 22989
rect 129575 22961 129609 22989
rect 129637 22961 129671 22989
rect 129699 22961 129747 22989
rect 129437 14175 129747 22961
rect 129437 14147 129485 14175
rect 129513 14147 129547 14175
rect 129575 14147 129609 14175
rect 129637 14147 129671 14175
rect 129699 14147 129747 14175
rect 129437 14113 129747 14147
rect 129437 14085 129485 14113
rect 129513 14085 129547 14113
rect 129575 14085 129609 14113
rect 129637 14085 129671 14113
rect 129699 14085 129747 14113
rect 129437 14051 129747 14085
rect 129437 14023 129485 14051
rect 129513 14023 129547 14051
rect 129575 14023 129609 14051
rect 129637 14023 129671 14051
rect 129699 14023 129747 14051
rect 129437 13989 129747 14023
rect 129437 13961 129485 13989
rect 129513 13961 129547 13989
rect 129575 13961 129609 13989
rect 129637 13961 129671 13989
rect 129699 13961 129747 13989
rect 129437 5175 129747 13961
rect 129437 5147 129485 5175
rect 129513 5147 129547 5175
rect 129575 5147 129609 5175
rect 129637 5147 129671 5175
rect 129699 5147 129747 5175
rect 129437 5113 129747 5147
rect 129437 5085 129485 5113
rect 129513 5085 129547 5113
rect 129575 5085 129609 5113
rect 129637 5085 129671 5113
rect 129699 5085 129747 5113
rect 129437 5051 129747 5085
rect 129437 5023 129485 5051
rect 129513 5023 129547 5051
rect 129575 5023 129609 5051
rect 129637 5023 129671 5051
rect 129699 5023 129747 5051
rect 129437 4989 129747 5023
rect 129437 4961 129485 4989
rect 129513 4961 129547 4989
rect 129575 4961 129609 4989
rect 129637 4961 129671 4989
rect 129699 4961 129747 4989
rect 129437 -560 129747 4961
rect 129437 -588 129485 -560
rect 129513 -588 129547 -560
rect 129575 -588 129609 -560
rect 129637 -588 129671 -560
rect 129699 -588 129747 -560
rect 129437 -622 129747 -588
rect 129437 -650 129485 -622
rect 129513 -650 129547 -622
rect 129575 -650 129609 -622
rect 129637 -650 129671 -622
rect 129699 -650 129747 -622
rect 129437 -684 129747 -650
rect 129437 -712 129485 -684
rect 129513 -712 129547 -684
rect 129575 -712 129609 -684
rect 129637 -712 129671 -684
rect 129699 -712 129747 -684
rect 129437 -746 129747 -712
rect 129437 -774 129485 -746
rect 129513 -774 129547 -746
rect 129575 -774 129609 -746
rect 129637 -774 129671 -746
rect 129699 -774 129747 -746
rect 129437 -822 129747 -774
rect 136577 119175 136887 124261
rect 136577 119147 136625 119175
rect 136653 119147 136687 119175
rect 136715 119147 136749 119175
rect 136777 119147 136811 119175
rect 136839 119147 136887 119175
rect 136577 119113 136887 119147
rect 136577 119085 136625 119113
rect 136653 119085 136687 119113
rect 136715 119085 136749 119113
rect 136777 119085 136811 119113
rect 136839 119085 136887 119113
rect 136577 119051 136887 119085
rect 136577 119023 136625 119051
rect 136653 119023 136687 119051
rect 136715 119023 136749 119051
rect 136777 119023 136811 119051
rect 136839 119023 136887 119051
rect 136577 118989 136887 119023
rect 136577 118961 136625 118989
rect 136653 118961 136687 118989
rect 136715 118961 136749 118989
rect 136777 118961 136811 118989
rect 136839 118961 136887 118989
rect 136577 110175 136887 118961
rect 136577 110147 136625 110175
rect 136653 110147 136687 110175
rect 136715 110147 136749 110175
rect 136777 110147 136811 110175
rect 136839 110147 136887 110175
rect 136577 110113 136887 110147
rect 136577 110085 136625 110113
rect 136653 110085 136687 110113
rect 136715 110085 136749 110113
rect 136777 110085 136811 110113
rect 136839 110085 136887 110113
rect 136577 110051 136887 110085
rect 136577 110023 136625 110051
rect 136653 110023 136687 110051
rect 136715 110023 136749 110051
rect 136777 110023 136811 110051
rect 136839 110023 136887 110051
rect 136577 109989 136887 110023
rect 136577 109961 136625 109989
rect 136653 109961 136687 109989
rect 136715 109961 136749 109989
rect 136777 109961 136811 109989
rect 136839 109961 136887 109989
rect 136577 101175 136887 109961
rect 136577 101147 136625 101175
rect 136653 101147 136687 101175
rect 136715 101147 136749 101175
rect 136777 101147 136811 101175
rect 136839 101147 136887 101175
rect 136577 101113 136887 101147
rect 136577 101085 136625 101113
rect 136653 101085 136687 101113
rect 136715 101085 136749 101113
rect 136777 101085 136811 101113
rect 136839 101085 136887 101113
rect 136577 101051 136887 101085
rect 136577 101023 136625 101051
rect 136653 101023 136687 101051
rect 136715 101023 136749 101051
rect 136777 101023 136811 101051
rect 136839 101023 136887 101051
rect 136577 100989 136887 101023
rect 136577 100961 136625 100989
rect 136653 100961 136687 100989
rect 136715 100961 136749 100989
rect 136777 100961 136811 100989
rect 136839 100961 136887 100989
rect 136577 92175 136887 100961
rect 136577 92147 136625 92175
rect 136653 92147 136687 92175
rect 136715 92147 136749 92175
rect 136777 92147 136811 92175
rect 136839 92147 136887 92175
rect 136577 92113 136887 92147
rect 136577 92085 136625 92113
rect 136653 92085 136687 92113
rect 136715 92085 136749 92113
rect 136777 92085 136811 92113
rect 136839 92085 136887 92113
rect 136577 92051 136887 92085
rect 136577 92023 136625 92051
rect 136653 92023 136687 92051
rect 136715 92023 136749 92051
rect 136777 92023 136811 92051
rect 136839 92023 136887 92051
rect 136577 91989 136887 92023
rect 136577 91961 136625 91989
rect 136653 91961 136687 91989
rect 136715 91961 136749 91989
rect 136777 91961 136811 91989
rect 136839 91961 136887 91989
rect 136577 83175 136887 91961
rect 136577 83147 136625 83175
rect 136653 83147 136687 83175
rect 136715 83147 136749 83175
rect 136777 83147 136811 83175
rect 136839 83147 136887 83175
rect 136577 83113 136887 83147
rect 136577 83085 136625 83113
rect 136653 83085 136687 83113
rect 136715 83085 136749 83113
rect 136777 83085 136811 83113
rect 136839 83085 136887 83113
rect 136577 83051 136887 83085
rect 136577 83023 136625 83051
rect 136653 83023 136687 83051
rect 136715 83023 136749 83051
rect 136777 83023 136811 83051
rect 136839 83023 136887 83051
rect 136577 82989 136887 83023
rect 136577 82961 136625 82989
rect 136653 82961 136687 82989
rect 136715 82961 136749 82989
rect 136777 82961 136811 82989
rect 136839 82961 136887 82989
rect 136577 74175 136887 82961
rect 136577 74147 136625 74175
rect 136653 74147 136687 74175
rect 136715 74147 136749 74175
rect 136777 74147 136811 74175
rect 136839 74147 136887 74175
rect 136577 74113 136887 74147
rect 136577 74085 136625 74113
rect 136653 74085 136687 74113
rect 136715 74085 136749 74113
rect 136777 74085 136811 74113
rect 136839 74085 136887 74113
rect 136577 74051 136887 74085
rect 136577 74023 136625 74051
rect 136653 74023 136687 74051
rect 136715 74023 136749 74051
rect 136777 74023 136811 74051
rect 136839 74023 136887 74051
rect 136577 73989 136887 74023
rect 136577 73961 136625 73989
rect 136653 73961 136687 73989
rect 136715 73961 136749 73989
rect 136777 73961 136811 73989
rect 136839 73961 136887 73989
rect 136577 65175 136887 73961
rect 136577 65147 136625 65175
rect 136653 65147 136687 65175
rect 136715 65147 136749 65175
rect 136777 65147 136811 65175
rect 136839 65147 136887 65175
rect 136577 65113 136887 65147
rect 136577 65085 136625 65113
rect 136653 65085 136687 65113
rect 136715 65085 136749 65113
rect 136777 65085 136811 65113
rect 136839 65085 136887 65113
rect 136577 65051 136887 65085
rect 136577 65023 136625 65051
rect 136653 65023 136687 65051
rect 136715 65023 136749 65051
rect 136777 65023 136811 65051
rect 136839 65023 136887 65051
rect 136577 64989 136887 65023
rect 136577 64961 136625 64989
rect 136653 64961 136687 64989
rect 136715 64961 136749 64989
rect 136777 64961 136811 64989
rect 136839 64961 136887 64989
rect 136577 56175 136887 64961
rect 136577 56147 136625 56175
rect 136653 56147 136687 56175
rect 136715 56147 136749 56175
rect 136777 56147 136811 56175
rect 136839 56147 136887 56175
rect 136577 56113 136887 56147
rect 136577 56085 136625 56113
rect 136653 56085 136687 56113
rect 136715 56085 136749 56113
rect 136777 56085 136811 56113
rect 136839 56085 136887 56113
rect 136577 56051 136887 56085
rect 136577 56023 136625 56051
rect 136653 56023 136687 56051
rect 136715 56023 136749 56051
rect 136777 56023 136811 56051
rect 136839 56023 136887 56051
rect 136577 55989 136887 56023
rect 136577 55961 136625 55989
rect 136653 55961 136687 55989
rect 136715 55961 136749 55989
rect 136777 55961 136811 55989
rect 136839 55961 136887 55989
rect 136577 47175 136887 55961
rect 136577 47147 136625 47175
rect 136653 47147 136687 47175
rect 136715 47147 136749 47175
rect 136777 47147 136811 47175
rect 136839 47147 136887 47175
rect 136577 47113 136887 47147
rect 136577 47085 136625 47113
rect 136653 47085 136687 47113
rect 136715 47085 136749 47113
rect 136777 47085 136811 47113
rect 136839 47085 136887 47113
rect 136577 47051 136887 47085
rect 136577 47023 136625 47051
rect 136653 47023 136687 47051
rect 136715 47023 136749 47051
rect 136777 47023 136811 47051
rect 136839 47023 136887 47051
rect 136577 46989 136887 47023
rect 136577 46961 136625 46989
rect 136653 46961 136687 46989
rect 136715 46961 136749 46989
rect 136777 46961 136811 46989
rect 136839 46961 136887 46989
rect 136577 38175 136887 46961
rect 136577 38147 136625 38175
rect 136653 38147 136687 38175
rect 136715 38147 136749 38175
rect 136777 38147 136811 38175
rect 136839 38147 136887 38175
rect 136577 38113 136887 38147
rect 136577 38085 136625 38113
rect 136653 38085 136687 38113
rect 136715 38085 136749 38113
rect 136777 38085 136811 38113
rect 136839 38085 136887 38113
rect 136577 38051 136887 38085
rect 136577 38023 136625 38051
rect 136653 38023 136687 38051
rect 136715 38023 136749 38051
rect 136777 38023 136811 38051
rect 136839 38023 136887 38051
rect 136577 37989 136887 38023
rect 136577 37961 136625 37989
rect 136653 37961 136687 37989
rect 136715 37961 136749 37989
rect 136777 37961 136811 37989
rect 136839 37961 136887 37989
rect 136577 29175 136887 37961
rect 136577 29147 136625 29175
rect 136653 29147 136687 29175
rect 136715 29147 136749 29175
rect 136777 29147 136811 29175
rect 136839 29147 136887 29175
rect 136577 29113 136887 29147
rect 136577 29085 136625 29113
rect 136653 29085 136687 29113
rect 136715 29085 136749 29113
rect 136777 29085 136811 29113
rect 136839 29085 136887 29113
rect 136577 29051 136887 29085
rect 136577 29023 136625 29051
rect 136653 29023 136687 29051
rect 136715 29023 136749 29051
rect 136777 29023 136811 29051
rect 136839 29023 136887 29051
rect 136577 28989 136887 29023
rect 136577 28961 136625 28989
rect 136653 28961 136687 28989
rect 136715 28961 136749 28989
rect 136777 28961 136811 28989
rect 136839 28961 136887 28989
rect 136577 20175 136887 28961
rect 136577 20147 136625 20175
rect 136653 20147 136687 20175
rect 136715 20147 136749 20175
rect 136777 20147 136811 20175
rect 136839 20147 136887 20175
rect 136577 20113 136887 20147
rect 136577 20085 136625 20113
rect 136653 20085 136687 20113
rect 136715 20085 136749 20113
rect 136777 20085 136811 20113
rect 136839 20085 136887 20113
rect 136577 20051 136887 20085
rect 136577 20023 136625 20051
rect 136653 20023 136687 20051
rect 136715 20023 136749 20051
rect 136777 20023 136811 20051
rect 136839 20023 136887 20051
rect 136577 19989 136887 20023
rect 136577 19961 136625 19989
rect 136653 19961 136687 19989
rect 136715 19961 136749 19989
rect 136777 19961 136811 19989
rect 136839 19961 136887 19989
rect 136577 11175 136887 19961
rect 136577 11147 136625 11175
rect 136653 11147 136687 11175
rect 136715 11147 136749 11175
rect 136777 11147 136811 11175
rect 136839 11147 136887 11175
rect 136577 11113 136887 11147
rect 136577 11085 136625 11113
rect 136653 11085 136687 11113
rect 136715 11085 136749 11113
rect 136777 11085 136811 11113
rect 136839 11085 136887 11113
rect 136577 11051 136887 11085
rect 136577 11023 136625 11051
rect 136653 11023 136687 11051
rect 136715 11023 136749 11051
rect 136777 11023 136811 11051
rect 136839 11023 136887 11051
rect 136577 10989 136887 11023
rect 136577 10961 136625 10989
rect 136653 10961 136687 10989
rect 136715 10961 136749 10989
rect 136777 10961 136811 10989
rect 136839 10961 136887 10989
rect 136577 2175 136887 10961
rect 136577 2147 136625 2175
rect 136653 2147 136687 2175
rect 136715 2147 136749 2175
rect 136777 2147 136811 2175
rect 136839 2147 136887 2175
rect 136577 2113 136887 2147
rect 136577 2085 136625 2113
rect 136653 2085 136687 2113
rect 136715 2085 136749 2113
rect 136777 2085 136811 2113
rect 136839 2085 136887 2113
rect 136577 2051 136887 2085
rect 136577 2023 136625 2051
rect 136653 2023 136687 2051
rect 136715 2023 136749 2051
rect 136777 2023 136811 2051
rect 136839 2023 136887 2051
rect 136577 1989 136887 2023
rect 136577 1961 136625 1989
rect 136653 1961 136687 1989
rect 136715 1961 136749 1989
rect 136777 1961 136811 1989
rect 136839 1961 136887 1989
rect 136577 -80 136887 1961
rect 136577 -108 136625 -80
rect 136653 -108 136687 -80
rect 136715 -108 136749 -80
rect 136777 -108 136811 -80
rect 136839 -108 136887 -80
rect 136577 -142 136887 -108
rect 136577 -170 136625 -142
rect 136653 -170 136687 -142
rect 136715 -170 136749 -142
rect 136777 -170 136811 -142
rect 136839 -170 136887 -142
rect 136577 -204 136887 -170
rect 136577 -232 136625 -204
rect 136653 -232 136687 -204
rect 136715 -232 136749 -204
rect 136777 -232 136811 -204
rect 136839 -232 136887 -204
rect 136577 -266 136887 -232
rect 136577 -294 136625 -266
rect 136653 -294 136687 -266
rect 136715 -294 136749 -266
rect 136777 -294 136811 -266
rect 136839 -294 136887 -266
rect 136577 -822 136887 -294
rect 138437 122175 138747 124261
rect 138437 122147 138485 122175
rect 138513 122147 138547 122175
rect 138575 122147 138609 122175
rect 138637 122147 138671 122175
rect 138699 122147 138747 122175
rect 138437 122113 138747 122147
rect 138437 122085 138485 122113
rect 138513 122085 138547 122113
rect 138575 122085 138609 122113
rect 138637 122085 138671 122113
rect 138699 122085 138747 122113
rect 138437 122051 138747 122085
rect 138437 122023 138485 122051
rect 138513 122023 138547 122051
rect 138575 122023 138609 122051
rect 138637 122023 138671 122051
rect 138699 122023 138747 122051
rect 138437 121989 138747 122023
rect 138437 121961 138485 121989
rect 138513 121961 138547 121989
rect 138575 121961 138609 121989
rect 138637 121961 138671 121989
rect 138699 121961 138747 121989
rect 138437 113175 138747 121961
rect 138437 113147 138485 113175
rect 138513 113147 138547 113175
rect 138575 113147 138609 113175
rect 138637 113147 138671 113175
rect 138699 113147 138747 113175
rect 138437 113113 138747 113147
rect 138437 113085 138485 113113
rect 138513 113085 138547 113113
rect 138575 113085 138609 113113
rect 138637 113085 138671 113113
rect 138699 113085 138747 113113
rect 138437 113051 138747 113085
rect 138437 113023 138485 113051
rect 138513 113023 138547 113051
rect 138575 113023 138609 113051
rect 138637 113023 138671 113051
rect 138699 113023 138747 113051
rect 138437 112989 138747 113023
rect 138437 112961 138485 112989
rect 138513 112961 138547 112989
rect 138575 112961 138609 112989
rect 138637 112961 138671 112989
rect 138699 112961 138747 112989
rect 138437 104175 138747 112961
rect 138437 104147 138485 104175
rect 138513 104147 138547 104175
rect 138575 104147 138609 104175
rect 138637 104147 138671 104175
rect 138699 104147 138747 104175
rect 138437 104113 138747 104147
rect 138437 104085 138485 104113
rect 138513 104085 138547 104113
rect 138575 104085 138609 104113
rect 138637 104085 138671 104113
rect 138699 104085 138747 104113
rect 138437 104051 138747 104085
rect 138437 104023 138485 104051
rect 138513 104023 138547 104051
rect 138575 104023 138609 104051
rect 138637 104023 138671 104051
rect 138699 104023 138747 104051
rect 138437 103989 138747 104023
rect 138437 103961 138485 103989
rect 138513 103961 138547 103989
rect 138575 103961 138609 103989
rect 138637 103961 138671 103989
rect 138699 103961 138747 103989
rect 138437 95175 138747 103961
rect 138437 95147 138485 95175
rect 138513 95147 138547 95175
rect 138575 95147 138609 95175
rect 138637 95147 138671 95175
rect 138699 95147 138747 95175
rect 138437 95113 138747 95147
rect 138437 95085 138485 95113
rect 138513 95085 138547 95113
rect 138575 95085 138609 95113
rect 138637 95085 138671 95113
rect 138699 95085 138747 95113
rect 138437 95051 138747 95085
rect 138437 95023 138485 95051
rect 138513 95023 138547 95051
rect 138575 95023 138609 95051
rect 138637 95023 138671 95051
rect 138699 95023 138747 95051
rect 138437 94989 138747 95023
rect 138437 94961 138485 94989
rect 138513 94961 138547 94989
rect 138575 94961 138609 94989
rect 138637 94961 138671 94989
rect 138699 94961 138747 94989
rect 138437 86175 138747 94961
rect 138437 86147 138485 86175
rect 138513 86147 138547 86175
rect 138575 86147 138609 86175
rect 138637 86147 138671 86175
rect 138699 86147 138747 86175
rect 138437 86113 138747 86147
rect 138437 86085 138485 86113
rect 138513 86085 138547 86113
rect 138575 86085 138609 86113
rect 138637 86085 138671 86113
rect 138699 86085 138747 86113
rect 138437 86051 138747 86085
rect 138437 86023 138485 86051
rect 138513 86023 138547 86051
rect 138575 86023 138609 86051
rect 138637 86023 138671 86051
rect 138699 86023 138747 86051
rect 138437 85989 138747 86023
rect 138437 85961 138485 85989
rect 138513 85961 138547 85989
rect 138575 85961 138609 85989
rect 138637 85961 138671 85989
rect 138699 85961 138747 85989
rect 138437 77175 138747 85961
rect 138437 77147 138485 77175
rect 138513 77147 138547 77175
rect 138575 77147 138609 77175
rect 138637 77147 138671 77175
rect 138699 77147 138747 77175
rect 138437 77113 138747 77147
rect 138437 77085 138485 77113
rect 138513 77085 138547 77113
rect 138575 77085 138609 77113
rect 138637 77085 138671 77113
rect 138699 77085 138747 77113
rect 138437 77051 138747 77085
rect 138437 77023 138485 77051
rect 138513 77023 138547 77051
rect 138575 77023 138609 77051
rect 138637 77023 138671 77051
rect 138699 77023 138747 77051
rect 138437 76989 138747 77023
rect 138437 76961 138485 76989
rect 138513 76961 138547 76989
rect 138575 76961 138609 76989
rect 138637 76961 138671 76989
rect 138699 76961 138747 76989
rect 138437 68175 138747 76961
rect 138437 68147 138485 68175
rect 138513 68147 138547 68175
rect 138575 68147 138609 68175
rect 138637 68147 138671 68175
rect 138699 68147 138747 68175
rect 138437 68113 138747 68147
rect 138437 68085 138485 68113
rect 138513 68085 138547 68113
rect 138575 68085 138609 68113
rect 138637 68085 138671 68113
rect 138699 68085 138747 68113
rect 138437 68051 138747 68085
rect 138437 68023 138485 68051
rect 138513 68023 138547 68051
rect 138575 68023 138609 68051
rect 138637 68023 138671 68051
rect 138699 68023 138747 68051
rect 138437 67989 138747 68023
rect 138437 67961 138485 67989
rect 138513 67961 138547 67989
rect 138575 67961 138609 67989
rect 138637 67961 138671 67989
rect 138699 67961 138747 67989
rect 138437 59175 138747 67961
rect 138437 59147 138485 59175
rect 138513 59147 138547 59175
rect 138575 59147 138609 59175
rect 138637 59147 138671 59175
rect 138699 59147 138747 59175
rect 138437 59113 138747 59147
rect 138437 59085 138485 59113
rect 138513 59085 138547 59113
rect 138575 59085 138609 59113
rect 138637 59085 138671 59113
rect 138699 59085 138747 59113
rect 138437 59051 138747 59085
rect 138437 59023 138485 59051
rect 138513 59023 138547 59051
rect 138575 59023 138609 59051
rect 138637 59023 138671 59051
rect 138699 59023 138747 59051
rect 138437 58989 138747 59023
rect 138437 58961 138485 58989
rect 138513 58961 138547 58989
rect 138575 58961 138609 58989
rect 138637 58961 138671 58989
rect 138699 58961 138747 58989
rect 138437 50175 138747 58961
rect 138437 50147 138485 50175
rect 138513 50147 138547 50175
rect 138575 50147 138609 50175
rect 138637 50147 138671 50175
rect 138699 50147 138747 50175
rect 138437 50113 138747 50147
rect 138437 50085 138485 50113
rect 138513 50085 138547 50113
rect 138575 50085 138609 50113
rect 138637 50085 138671 50113
rect 138699 50085 138747 50113
rect 138437 50051 138747 50085
rect 138437 50023 138485 50051
rect 138513 50023 138547 50051
rect 138575 50023 138609 50051
rect 138637 50023 138671 50051
rect 138699 50023 138747 50051
rect 138437 49989 138747 50023
rect 138437 49961 138485 49989
rect 138513 49961 138547 49989
rect 138575 49961 138609 49989
rect 138637 49961 138671 49989
rect 138699 49961 138747 49989
rect 138437 41175 138747 49961
rect 138437 41147 138485 41175
rect 138513 41147 138547 41175
rect 138575 41147 138609 41175
rect 138637 41147 138671 41175
rect 138699 41147 138747 41175
rect 138437 41113 138747 41147
rect 138437 41085 138485 41113
rect 138513 41085 138547 41113
rect 138575 41085 138609 41113
rect 138637 41085 138671 41113
rect 138699 41085 138747 41113
rect 138437 41051 138747 41085
rect 138437 41023 138485 41051
rect 138513 41023 138547 41051
rect 138575 41023 138609 41051
rect 138637 41023 138671 41051
rect 138699 41023 138747 41051
rect 138437 40989 138747 41023
rect 138437 40961 138485 40989
rect 138513 40961 138547 40989
rect 138575 40961 138609 40989
rect 138637 40961 138671 40989
rect 138699 40961 138747 40989
rect 138437 32175 138747 40961
rect 138437 32147 138485 32175
rect 138513 32147 138547 32175
rect 138575 32147 138609 32175
rect 138637 32147 138671 32175
rect 138699 32147 138747 32175
rect 138437 32113 138747 32147
rect 138437 32085 138485 32113
rect 138513 32085 138547 32113
rect 138575 32085 138609 32113
rect 138637 32085 138671 32113
rect 138699 32085 138747 32113
rect 138437 32051 138747 32085
rect 138437 32023 138485 32051
rect 138513 32023 138547 32051
rect 138575 32023 138609 32051
rect 138637 32023 138671 32051
rect 138699 32023 138747 32051
rect 138437 31989 138747 32023
rect 138437 31961 138485 31989
rect 138513 31961 138547 31989
rect 138575 31961 138609 31989
rect 138637 31961 138671 31989
rect 138699 31961 138747 31989
rect 138437 23175 138747 31961
rect 138437 23147 138485 23175
rect 138513 23147 138547 23175
rect 138575 23147 138609 23175
rect 138637 23147 138671 23175
rect 138699 23147 138747 23175
rect 138437 23113 138747 23147
rect 138437 23085 138485 23113
rect 138513 23085 138547 23113
rect 138575 23085 138609 23113
rect 138637 23085 138671 23113
rect 138699 23085 138747 23113
rect 138437 23051 138747 23085
rect 138437 23023 138485 23051
rect 138513 23023 138547 23051
rect 138575 23023 138609 23051
rect 138637 23023 138671 23051
rect 138699 23023 138747 23051
rect 138437 22989 138747 23023
rect 138437 22961 138485 22989
rect 138513 22961 138547 22989
rect 138575 22961 138609 22989
rect 138637 22961 138671 22989
rect 138699 22961 138747 22989
rect 138437 14175 138747 22961
rect 138437 14147 138485 14175
rect 138513 14147 138547 14175
rect 138575 14147 138609 14175
rect 138637 14147 138671 14175
rect 138699 14147 138747 14175
rect 138437 14113 138747 14147
rect 138437 14085 138485 14113
rect 138513 14085 138547 14113
rect 138575 14085 138609 14113
rect 138637 14085 138671 14113
rect 138699 14085 138747 14113
rect 138437 14051 138747 14085
rect 138437 14023 138485 14051
rect 138513 14023 138547 14051
rect 138575 14023 138609 14051
rect 138637 14023 138671 14051
rect 138699 14023 138747 14051
rect 138437 13989 138747 14023
rect 138437 13961 138485 13989
rect 138513 13961 138547 13989
rect 138575 13961 138609 13989
rect 138637 13961 138671 13989
rect 138699 13961 138747 13989
rect 138437 5175 138747 13961
rect 138437 5147 138485 5175
rect 138513 5147 138547 5175
rect 138575 5147 138609 5175
rect 138637 5147 138671 5175
rect 138699 5147 138747 5175
rect 138437 5113 138747 5147
rect 138437 5085 138485 5113
rect 138513 5085 138547 5113
rect 138575 5085 138609 5113
rect 138637 5085 138671 5113
rect 138699 5085 138747 5113
rect 138437 5051 138747 5085
rect 138437 5023 138485 5051
rect 138513 5023 138547 5051
rect 138575 5023 138609 5051
rect 138637 5023 138671 5051
rect 138699 5023 138747 5051
rect 138437 4989 138747 5023
rect 138437 4961 138485 4989
rect 138513 4961 138547 4989
rect 138575 4961 138609 4989
rect 138637 4961 138671 4989
rect 138699 4961 138747 4989
rect 138437 -560 138747 4961
rect 138437 -588 138485 -560
rect 138513 -588 138547 -560
rect 138575 -588 138609 -560
rect 138637 -588 138671 -560
rect 138699 -588 138747 -560
rect 138437 -622 138747 -588
rect 138437 -650 138485 -622
rect 138513 -650 138547 -622
rect 138575 -650 138609 -622
rect 138637 -650 138671 -622
rect 138699 -650 138747 -622
rect 138437 -684 138747 -650
rect 138437 -712 138485 -684
rect 138513 -712 138547 -684
rect 138575 -712 138609 -684
rect 138637 -712 138671 -684
rect 138699 -712 138747 -684
rect 138437 -746 138747 -712
rect 138437 -774 138485 -746
rect 138513 -774 138547 -746
rect 138575 -774 138609 -746
rect 138637 -774 138671 -746
rect 138699 -774 138747 -746
rect 138437 -822 138747 -774
rect 145577 119175 145887 124261
rect 145577 119147 145625 119175
rect 145653 119147 145687 119175
rect 145715 119147 145749 119175
rect 145777 119147 145811 119175
rect 145839 119147 145887 119175
rect 145577 119113 145887 119147
rect 145577 119085 145625 119113
rect 145653 119085 145687 119113
rect 145715 119085 145749 119113
rect 145777 119085 145811 119113
rect 145839 119085 145887 119113
rect 145577 119051 145887 119085
rect 145577 119023 145625 119051
rect 145653 119023 145687 119051
rect 145715 119023 145749 119051
rect 145777 119023 145811 119051
rect 145839 119023 145887 119051
rect 145577 118989 145887 119023
rect 145577 118961 145625 118989
rect 145653 118961 145687 118989
rect 145715 118961 145749 118989
rect 145777 118961 145811 118989
rect 145839 118961 145887 118989
rect 145577 110175 145887 118961
rect 145577 110147 145625 110175
rect 145653 110147 145687 110175
rect 145715 110147 145749 110175
rect 145777 110147 145811 110175
rect 145839 110147 145887 110175
rect 145577 110113 145887 110147
rect 145577 110085 145625 110113
rect 145653 110085 145687 110113
rect 145715 110085 145749 110113
rect 145777 110085 145811 110113
rect 145839 110085 145887 110113
rect 145577 110051 145887 110085
rect 145577 110023 145625 110051
rect 145653 110023 145687 110051
rect 145715 110023 145749 110051
rect 145777 110023 145811 110051
rect 145839 110023 145887 110051
rect 145577 109989 145887 110023
rect 145577 109961 145625 109989
rect 145653 109961 145687 109989
rect 145715 109961 145749 109989
rect 145777 109961 145811 109989
rect 145839 109961 145887 109989
rect 145577 101175 145887 109961
rect 145577 101147 145625 101175
rect 145653 101147 145687 101175
rect 145715 101147 145749 101175
rect 145777 101147 145811 101175
rect 145839 101147 145887 101175
rect 145577 101113 145887 101147
rect 145577 101085 145625 101113
rect 145653 101085 145687 101113
rect 145715 101085 145749 101113
rect 145777 101085 145811 101113
rect 145839 101085 145887 101113
rect 145577 101051 145887 101085
rect 145577 101023 145625 101051
rect 145653 101023 145687 101051
rect 145715 101023 145749 101051
rect 145777 101023 145811 101051
rect 145839 101023 145887 101051
rect 145577 100989 145887 101023
rect 145577 100961 145625 100989
rect 145653 100961 145687 100989
rect 145715 100961 145749 100989
rect 145777 100961 145811 100989
rect 145839 100961 145887 100989
rect 145577 92175 145887 100961
rect 145577 92147 145625 92175
rect 145653 92147 145687 92175
rect 145715 92147 145749 92175
rect 145777 92147 145811 92175
rect 145839 92147 145887 92175
rect 145577 92113 145887 92147
rect 145577 92085 145625 92113
rect 145653 92085 145687 92113
rect 145715 92085 145749 92113
rect 145777 92085 145811 92113
rect 145839 92085 145887 92113
rect 145577 92051 145887 92085
rect 145577 92023 145625 92051
rect 145653 92023 145687 92051
rect 145715 92023 145749 92051
rect 145777 92023 145811 92051
rect 145839 92023 145887 92051
rect 145577 91989 145887 92023
rect 145577 91961 145625 91989
rect 145653 91961 145687 91989
rect 145715 91961 145749 91989
rect 145777 91961 145811 91989
rect 145839 91961 145887 91989
rect 145577 83175 145887 91961
rect 145577 83147 145625 83175
rect 145653 83147 145687 83175
rect 145715 83147 145749 83175
rect 145777 83147 145811 83175
rect 145839 83147 145887 83175
rect 145577 83113 145887 83147
rect 145577 83085 145625 83113
rect 145653 83085 145687 83113
rect 145715 83085 145749 83113
rect 145777 83085 145811 83113
rect 145839 83085 145887 83113
rect 145577 83051 145887 83085
rect 145577 83023 145625 83051
rect 145653 83023 145687 83051
rect 145715 83023 145749 83051
rect 145777 83023 145811 83051
rect 145839 83023 145887 83051
rect 145577 82989 145887 83023
rect 145577 82961 145625 82989
rect 145653 82961 145687 82989
rect 145715 82961 145749 82989
rect 145777 82961 145811 82989
rect 145839 82961 145887 82989
rect 145577 74175 145887 82961
rect 145577 74147 145625 74175
rect 145653 74147 145687 74175
rect 145715 74147 145749 74175
rect 145777 74147 145811 74175
rect 145839 74147 145887 74175
rect 145577 74113 145887 74147
rect 145577 74085 145625 74113
rect 145653 74085 145687 74113
rect 145715 74085 145749 74113
rect 145777 74085 145811 74113
rect 145839 74085 145887 74113
rect 145577 74051 145887 74085
rect 145577 74023 145625 74051
rect 145653 74023 145687 74051
rect 145715 74023 145749 74051
rect 145777 74023 145811 74051
rect 145839 74023 145887 74051
rect 145577 73989 145887 74023
rect 145577 73961 145625 73989
rect 145653 73961 145687 73989
rect 145715 73961 145749 73989
rect 145777 73961 145811 73989
rect 145839 73961 145887 73989
rect 145577 65175 145887 73961
rect 145577 65147 145625 65175
rect 145653 65147 145687 65175
rect 145715 65147 145749 65175
rect 145777 65147 145811 65175
rect 145839 65147 145887 65175
rect 145577 65113 145887 65147
rect 145577 65085 145625 65113
rect 145653 65085 145687 65113
rect 145715 65085 145749 65113
rect 145777 65085 145811 65113
rect 145839 65085 145887 65113
rect 145577 65051 145887 65085
rect 145577 65023 145625 65051
rect 145653 65023 145687 65051
rect 145715 65023 145749 65051
rect 145777 65023 145811 65051
rect 145839 65023 145887 65051
rect 145577 64989 145887 65023
rect 145577 64961 145625 64989
rect 145653 64961 145687 64989
rect 145715 64961 145749 64989
rect 145777 64961 145811 64989
rect 145839 64961 145887 64989
rect 145577 56175 145887 64961
rect 145577 56147 145625 56175
rect 145653 56147 145687 56175
rect 145715 56147 145749 56175
rect 145777 56147 145811 56175
rect 145839 56147 145887 56175
rect 145577 56113 145887 56147
rect 145577 56085 145625 56113
rect 145653 56085 145687 56113
rect 145715 56085 145749 56113
rect 145777 56085 145811 56113
rect 145839 56085 145887 56113
rect 145577 56051 145887 56085
rect 145577 56023 145625 56051
rect 145653 56023 145687 56051
rect 145715 56023 145749 56051
rect 145777 56023 145811 56051
rect 145839 56023 145887 56051
rect 145577 55989 145887 56023
rect 145577 55961 145625 55989
rect 145653 55961 145687 55989
rect 145715 55961 145749 55989
rect 145777 55961 145811 55989
rect 145839 55961 145887 55989
rect 145577 47175 145887 55961
rect 145577 47147 145625 47175
rect 145653 47147 145687 47175
rect 145715 47147 145749 47175
rect 145777 47147 145811 47175
rect 145839 47147 145887 47175
rect 145577 47113 145887 47147
rect 145577 47085 145625 47113
rect 145653 47085 145687 47113
rect 145715 47085 145749 47113
rect 145777 47085 145811 47113
rect 145839 47085 145887 47113
rect 145577 47051 145887 47085
rect 145577 47023 145625 47051
rect 145653 47023 145687 47051
rect 145715 47023 145749 47051
rect 145777 47023 145811 47051
rect 145839 47023 145887 47051
rect 145577 46989 145887 47023
rect 145577 46961 145625 46989
rect 145653 46961 145687 46989
rect 145715 46961 145749 46989
rect 145777 46961 145811 46989
rect 145839 46961 145887 46989
rect 145577 38175 145887 46961
rect 145577 38147 145625 38175
rect 145653 38147 145687 38175
rect 145715 38147 145749 38175
rect 145777 38147 145811 38175
rect 145839 38147 145887 38175
rect 145577 38113 145887 38147
rect 145577 38085 145625 38113
rect 145653 38085 145687 38113
rect 145715 38085 145749 38113
rect 145777 38085 145811 38113
rect 145839 38085 145887 38113
rect 145577 38051 145887 38085
rect 145577 38023 145625 38051
rect 145653 38023 145687 38051
rect 145715 38023 145749 38051
rect 145777 38023 145811 38051
rect 145839 38023 145887 38051
rect 145577 37989 145887 38023
rect 145577 37961 145625 37989
rect 145653 37961 145687 37989
rect 145715 37961 145749 37989
rect 145777 37961 145811 37989
rect 145839 37961 145887 37989
rect 145577 29175 145887 37961
rect 145577 29147 145625 29175
rect 145653 29147 145687 29175
rect 145715 29147 145749 29175
rect 145777 29147 145811 29175
rect 145839 29147 145887 29175
rect 145577 29113 145887 29147
rect 145577 29085 145625 29113
rect 145653 29085 145687 29113
rect 145715 29085 145749 29113
rect 145777 29085 145811 29113
rect 145839 29085 145887 29113
rect 145577 29051 145887 29085
rect 145577 29023 145625 29051
rect 145653 29023 145687 29051
rect 145715 29023 145749 29051
rect 145777 29023 145811 29051
rect 145839 29023 145887 29051
rect 145577 28989 145887 29023
rect 145577 28961 145625 28989
rect 145653 28961 145687 28989
rect 145715 28961 145749 28989
rect 145777 28961 145811 28989
rect 145839 28961 145887 28989
rect 145577 20175 145887 28961
rect 145577 20147 145625 20175
rect 145653 20147 145687 20175
rect 145715 20147 145749 20175
rect 145777 20147 145811 20175
rect 145839 20147 145887 20175
rect 145577 20113 145887 20147
rect 145577 20085 145625 20113
rect 145653 20085 145687 20113
rect 145715 20085 145749 20113
rect 145777 20085 145811 20113
rect 145839 20085 145887 20113
rect 145577 20051 145887 20085
rect 145577 20023 145625 20051
rect 145653 20023 145687 20051
rect 145715 20023 145749 20051
rect 145777 20023 145811 20051
rect 145839 20023 145887 20051
rect 145577 19989 145887 20023
rect 145577 19961 145625 19989
rect 145653 19961 145687 19989
rect 145715 19961 145749 19989
rect 145777 19961 145811 19989
rect 145839 19961 145887 19989
rect 145577 11175 145887 19961
rect 145577 11147 145625 11175
rect 145653 11147 145687 11175
rect 145715 11147 145749 11175
rect 145777 11147 145811 11175
rect 145839 11147 145887 11175
rect 145577 11113 145887 11147
rect 145577 11085 145625 11113
rect 145653 11085 145687 11113
rect 145715 11085 145749 11113
rect 145777 11085 145811 11113
rect 145839 11085 145887 11113
rect 145577 11051 145887 11085
rect 145577 11023 145625 11051
rect 145653 11023 145687 11051
rect 145715 11023 145749 11051
rect 145777 11023 145811 11051
rect 145839 11023 145887 11051
rect 145577 10989 145887 11023
rect 145577 10961 145625 10989
rect 145653 10961 145687 10989
rect 145715 10961 145749 10989
rect 145777 10961 145811 10989
rect 145839 10961 145887 10989
rect 145577 2175 145887 10961
rect 145577 2147 145625 2175
rect 145653 2147 145687 2175
rect 145715 2147 145749 2175
rect 145777 2147 145811 2175
rect 145839 2147 145887 2175
rect 145577 2113 145887 2147
rect 145577 2085 145625 2113
rect 145653 2085 145687 2113
rect 145715 2085 145749 2113
rect 145777 2085 145811 2113
rect 145839 2085 145887 2113
rect 145577 2051 145887 2085
rect 145577 2023 145625 2051
rect 145653 2023 145687 2051
rect 145715 2023 145749 2051
rect 145777 2023 145811 2051
rect 145839 2023 145887 2051
rect 145577 1989 145887 2023
rect 145577 1961 145625 1989
rect 145653 1961 145687 1989
rect 145715 1961 145749 1989
rect 145777 1961 145811 1989
rect 145839 1961 145887 1989
rect 145577 -80 145887 1961
rect 145577 -108 145625 -80
rect 145653 -108 145687 -80
rect 145715 -108 145749 -80
rect 145777 -108 145811 -80
rect 145839 -108 145887 -80
rect 145577 -142 145887 -108
rect 145577 -170 145625 -142
rect 145653 -170 145687 -142
rect 145715 -170 145749 -142
rect 145777 -170 145811 -142
rect 145839 -170 145887 -142
rect 145577 -204 145887 -170
rect 145577 -232 145625 -204
rect 145653 -232 145687 -204
rect 145715 -232 145749 -204
rect 145777 -232 145811 -204
rect 145839 -232 145887 -204
rect 145577 -266 145887 -232
rect 145577 -294 145625 -266
rect 145653 -294 145687 -266
rect 145715 -294 145749 -266
rect 145777 -294 145811 -266
rect 145839 -294 145887 -266
rect 145577 -822 145887 -294
rect 147437 122175 147747 124261
rect 147437 122147 147485 122175
rect 147513 122147 147547 122175
rect 147575 122147 147609 122175
rect 147637 122147 147671 122175
rect 147699 122147 147747 122175
rect 147437 122113 147747 122147
rect 147437 122085 147485 122113
rect 147513 122085 147547 122113
rect 147575 122085 147609 122113
rect 147637 122085 147671 122113
rect 147699 122085 147747 122113
rect 147437 122051 147747 122085
rect 147437 122023 147485 122051
rect 147513 122023 147547 122051
rect 147575 122023 147609 122051
rect 147637 122023 147671 122051
rect 147699 122023 147747 122051
rect 147437 121989 147747 122023
rect 147437 121961 147485 121989
rect 147513 121961 147547 121989
rect 147575 121961 147609 121989
rect 147637 121961 147671 121989
rect 147699 121961 147747 121989
rect 147437 113175 147747 121961
rect 147437 113147 147485 113175
rect 147513 113147 147547 113175
rect 147575 113147 147609 113175
rect 147637 113147 147671 113175
rect 147699 113147 147747 113175
rect 147437 113113 147747 113147
rect 147437 113085 147485 113113
rect 147513 113085 147547 113113
rect 147575 113085 147609 113113
rect 147637 113085 147671 113113
rect 147699 113085 147747 113113
rect 147437 113051 147747 113085
rect 147437 113023 147485 113051
rect 147513 113023 147547 113051
rect 147575 113023 147609 113051
rect 147637 113023 147671 113051
rect 147699 113023 147747 113051
rect 147437 112989 147747 113023
rect 147437 112961 147485 112989
rect 147513 112961 147547 112989
rect 147575 112961 147609 112989
rect 147637 112961 147671 112989
rect 147699 112961 147747 112989
rect 147437 104175 147747 112961
rect 147437 104147 147485 104175
rect 147513 104147 147547 104175
rect 147575 104147 147609 104175
rect 147637 104147 147671 104175
rect 147699 104147 147747 104175
rect 147437 104113 147747 104147
rect 147437 104085 147485 104113
rect 147513 104085 147547 104113
rect 147575 104085 147609 104113
rect 147637 104085 147671 104113
rect 147699 104085 147747 104113
rect 147437 104051 147747 104085
rect 147437 104023 147485 104051
rect 147513 104023 147547 104051
rect 147575 104023 147609 104051
rect 147637 104023 147671 104051
rect 147699 104023 147747 104051
rect 147437 103989 147747 104023
rect 147437 103961 147485 103989
rect 147513 103961 147547 103989
rect 147575 103961 147609 103989
rect 147637 103961 147671 103989
rect 147699 103961 147747 103989
rect 147437 95175 147747 103961
rect 147437 95147 147485 95175
rect 147513 95147 147547 95175
rect 147575 95147 147609 95175
rect 147637 95147 147671 95175
rect 147699 95147 147747 95175
rect 147437 95113 147747 95147
rect 147437 95085 147485 95113
rect 147513 95085 147547 95113
rect 147575 95085 147609 95113
rect 147637 95085 147671 95113
rect 147699 95085 147747 95113
rect 147437 95051 147747 95085
rect 147437 95023 147485 95051
rect 147513 95023 147547 95051
rect 147575 95023 147609 95051
rect 147637 95023 147671 95051
rect 147699 95023 147747 95051
rect 147437 94989 147747 95023
rect 147437 94961 147485 94989
rect 147513 94961 147547 94989
rect 147575 94961 147609 94989
rect 147637 94961 147671 94989
rect 147699 94961 147747 94989
rect 147437 86175 147747 94961
rect 147437 86147 147485 86175
rect 147513 86147 147547 86175
rect 147575 86147 147609 86175
rect 147637 86147 147671 86175
rect 147699 86147 147747 86175
rect 147437 86113 147747 86147
rect 147437 86085 147485 86113
rect 147513 86085 147547 86113
rect 147575 86085 147609 86113
rect 147637 86085 147671 86113
rect 147699 86085 147747 86113
rect 147437 86051 147747 86085
rect 147437 86023 147485 86051
rect 147513 86023 147547 86051
rect 147575 86023 147609 86051
rect 147637 86023 147671 86051
rect 147699 86023 147747 86051
rect 147437 85989 147747 86023
rect 147437 85961 147485 85989
rect 147513 85961 147547 85989
rect 147575 85961 147609 85989
rect 147637 85961 147671 85989
rect 147699 85961 147747 85989
rect 147437 77175 147747 85961
rect 147437 77147 147485 77175
rect 147513 77147 147547 77175
rect 147575 77147 147609 77175
rect 147637 77147 147671 77175
rect 147699 77147 147747 77175
rect 147437 77113 147747 77147
rect 147437 77085 147485 77113
rect 147513 77085 147547 77113
rect 147575 77085 147609 77113
rect 147637 77085 147671 77113
rect 147699 77085 147747 77113
rect 147437 77051 147747 77085
rect 147437 77023 147485 77051
rect 147513 77023 147547 77051
rect 147575 77023 147609 77051
rect 147637 77023 147671 77051
rect 147699 77023 147747 77051
rect 147437 76989 147747 77023
rect 147437 76961 147485 76989
rect 147513 76961 147547 76989
rect 147575 76961 147609 76989
rect 147637 76961 147671 76989
rect 147699 76961 147747 76989
rect 147437 68175 147747 76961
rect 147437 68147 147485 68175
rect 147513 68147 147547 68175
rect 147575 68147 147609 68175
rect 147637 68147 147671 68175
rect 147699 68147 147747 68175
rect 147437 68113 147747 68147
rect 147437 68085 147485 68113
rect 147513 68085 147547 68113
rect 147575 68085 147609 68113
rect 147637 68085 147671 68113
rect 147699 68085 147747 68113
rect 147437 68051 147747 68085
rect 147437 68023 147485 68051
rect 147513 68023 147547 68051
rect 147575 68023 147609 68051
rect 147637 68023 147671 68051
rect 147699 68023 147747 68051
rect 147437 67989 147747 68023
rect 147437 67961 147485 67989
rect 147513 67961 147547 67989
rect 147575 67961 147609 67989
rect 147637 67961 147671 67989
rect 147699 67961 147747 67989
rect 147437 59175 147747 67961
rect 147437 59147 147485 59175
rect 147513 59147 147547 59175
rect 147575 59147 147609 59175
rect 147637 59147 147671 59175
rect 147699 59147 147747 59175
rect 147437 59113 147747 59147
rect 147437 59085 147485 59113
rect 147513 59085 147547 59113
rect 147575 59085 147609 59113
rect 147637 59085 147671 59113
rect 147699 59085 147747 59113
rect 147437 59051 147747 59085
rect 147437 59023 147485 59051
rect 147513 59023 147547 59051
rect 147575 59023 147609 59051
rect 147637 59023 147671 59051
rect 147699 59023 147747 59051
rect 147437 58989 147747 59023
rect 147437 58961 147485 58989
rect 147513 58961 147547 58989
rect 147575 58961 147609 58989
rect 147637 58961 147671 58989
rect 147699 58961 147747 58989
rect 147437 50175 147747 58961
rect 147437 50147 147485 50175
rect 147513 50147 147547 50175
rect 147575 50147 147609 50175
rect 147637 50147 147671 50175
rect 147699 50147 147747 50175
rect 147437 50113 147747 50147
rect 147437 50085 147485 50113
rect 147513 50085 147547 50113
rect 147575 50085 147609 50113
rect 147637 50085 147671 50113
rect 147699 50085 147747 50113
rect 147437 50051 147747 50085
rect 147437 50023 147485 50051
rect 147513 50023 147547 50051
rect 147575 50023 147609 50051
rect 147637 50023 147671 50051
rect 147699 50023 147747 50051
rect 147437 49989 147747 50023
rect 147437 49961 147485 49989
rect 147513 49961 147547 49989
rect 147575 49961 147609 49989
rect 147637 49961 147671 49989
rect 147699 49961 147747 49989
rect 147437 41175 147747 49961
rect 147437 41147 147485 41175
rect 147513 41147 147547 41175
rect 147575 41147 147609 41175
rect 147637 41147 147671 41175
rect 147699 41147 147747 41175
rect 147437 41113 147747 41147
rect 147437 41085 147485 41113
rect 147513 41085 147547 41113
rect 147575 41085 147609 41113
rect 147637 41085 147671 41113
rect 147699 41085 147747 41113
rect 147437 41051 147747 41085
rect 147437 41023 147485 41051
rect 147513 41023 147547 41051
rect 147575 41023 147609 41051
rect 147637 41023 147671 41051
rect 147699 41023 147747 41051
rect 147437 40989 147747 41023
rect 147437 40961 147485 40989
rect 147513 40961 147547 40989
rect 147575 40961 147609 40989
rect 147637 40961 147671 40989
rect 147699 40961 147747 40989
rect 147437 32175 147747 40961
rect 147437 32147 147485 32175
rect 147513 32147 147547 32175
rect 147575 32147 147609 32175
rect 147637 32147 147671 32175
rect 147699 32147 147747 32175
rect 147437 32113 147747 32147
rect 147437 32085 147485 32113
rect 147513 32085 147547 32113
rect 147575 32085 147609 32113
rect 147637 32085 147671 32113
rect 147699 32085 147747 32113
rect 147437 32051 147747 32085
rect 147437 32023 147485 32051
rect 147513 32023 147547 32051
rect 147575 32023 147609 32051
rect 147637 32023 147671 32051
rect 147699 32023 147747 32051
rect 147437 31989 147747 32023
rect 147437 31961 147485 31989
rect 147513 31961 147547 31989
rect 147575 31961 147609 31989
rect 147637 31961 147671 31989
rect 147699 31961 147747 31989
rect 147437 23175 147747 31961
rect 147437 23147 147485 23175
rect 147513 23147 147547 23175
rect 147575 23147 147609 23175
rect 147637 23147 147671 23175
rect 147699 23147 147747 23175
rect 147437 23113 147747 23147
rect 147437 23085 147485 23113
rect 147513 23085 147547 23113
rect 147575 23085 147609 23113
rect 147637 23085 147671 23113
rect 147699 23085 147747 23113
rect 147437 23051 147747 23085
rect 147437 23023 147485 23051
rect 147513 23023 147547 23051
rect 147575 23023 147609 23051
rect 147637 23023 147671 23051
rect 147699 23023 147747 23051
rect 147437 22989 147747 23023
rect 147437 22961 147485 22989
rect 147513 22961 147547 22989
rect 147575 22961 147609 22989
rect 147637 22961 147671 22989
rect 147699 22961 147747 22989
rect 147437 14175 147747 22961
rect 147437 14147 147485 14175
rect 147513 14147 147547 14175
rect 147575 14147 147609 14175
rect 147637 14147 147671 14175
rect 147699 14147 147747 14175
rect 147437 14113 147747 14147
rect 147437 14085 147485 14113
rect 147513 14085 147547 14113
rect 147575 14085 147609 14113
rect 147637 14085 147671 14113
rect 147699 14085 147747 14113
rect 147437 14051 147747 14085
rect 147437 14023 147485 14051
rect 147513 14023 147547 14051
rect 147575 14023 147609 14051
rect 147637 14023 147671 14051
rect 147699 14023 147747 14051
rect 147437 13989 147747 14023
rect 147437 13961 147485 13989
rect 147513 13961 147547 13989
rect 147575 13961 147609 13989
rect 147637 13961 147671 13989
rect 147699 13961 147747 13989
rect 147437 5175 147747 13961
rect 147437 5147 147485 5175
rect 147513 5147 147547 5175
rect 147575 5147 147609 5175
rect 147637 5147 147671 5175
rect 147699 5147 147747 5175
rect 147437 5113 147747 5147
rect 147437 5085 147485 5113
rect 147513 5085 147547 5113
rect 147575 5085 147609 5113
rect 147637 5085 147671 5113
rect 147699 5085 147747 5113
rect 147437 5051 147747 5085
rect 147437 5023 147485 5051
rect 147513 5023 147547 5051
rect 147575 5023 147609 5051
rect 147637 5023 147671 5051
rect 147699 5023 147747 5051
rect 147437 4989 147747 5023
rect 147437 4961 147485 4989
rect 147513 4961 147547 4989
rect 147575 4961 147609 4989
rect 147637 4961 147671 4989
rect 147699 4961 147747 4989
rect 147437 -560 147747 4961
rect 147437 -588 147485 -560
rect 147513 -588 147547 -560
rect 147575 -588 147609 -560
rect 147637 -588 147671 -560
rect 147699 -588 147747 -560
rect 147437 -622 147747 -588
rect 147437 -650 147485 -622
rect 147513 -650 147547 -622
rect 147575 -650 147609 -622
rect 147637 -650 147671 -622
rect 147699 -650 147747 -622
rect 147437 -684 147747 -650
rect 147437 -712 147485 -684
rect 147513 -712 147547 -684
rect 147575 -712 147609 -684
rect 147637 -712 147671 -684
rect 147699 -712 147747 -684
rect 147437 -746 147747 -712
rect 147437 -774 147485 -746
rect 147513 -774 147547 -746
rect 147575 -774 147609 -746
rect 147637 -774 147671 -746
rect 147699 -774 147747 -746
rect 147437 -822 147747 -774
rect 154577 119175 154887 127961
rect 154577 119147 154625 119175
rect 154653 119147 154687 119175
rect 154715 119147 154749 119175
rect 154777 119147 154811 119175
rect 154839 119147 154887 119175
rect 154577 119113 154887 119147
rect 154577 119085 154625 119113
rect 154653 119085 154687 119113
rect 154715 119085 154749 119113
rect 154777 119085 154811 119113
rect 154839 119085 154887 119113
rect 154577 119051 154887 119085
rect 154577 119023 154625 119051
rect 154653 119023 154687 119051
rect 154715 119023 154749 119051
rect 154777 119023 154811 119051
rect 154839 119023 154887 119051
rect 154577 118989 154887 119023
rect 154577 118961 154625 118989
rect 154653 118961 154687 118989
rect 154715 118961 154749 118989
rect 154777 118961 154811 118989
rect 154839 118961 154887 118989
rect 154577 110175 154887 118961
rect 154577 110147 154625 110175
rect 154653 110147 154687 110175
rect 154715 110147 154749 110175
rect 154777 110147 154811 110175
rect 154839 110147 154887 110175
rect 154577 110113 154887 110147
rect 154577 110085 154625 110113
rect 154653 110085 154687 110113
rect 154715 110085 154749 110113
rect 154777 110085 154811 110113
rect 154839 110085 154887 110113
rect 154577 110051 154887 110085
rect 154577 110023 154625 110051
rect 154653 110023 154687 110051
rect 154715 110023 154749 110051
rect 154777 110023 154811 110051
rect 154839 110023 154887 110051
rect 154577 109989 154887 110023
rect 154577 109961 154625 109989
rect 154653 109961 154687 109989
rect 154715 109961 154749 109989
rect 154777 109961 154811 109989
rect 154839 109961 154887 109989
rect 154577 101175 154887 109961
rect 154577 101147 154625 101175
rect 154653 101147 154687 101175
rect 154715 101147 154749 101175
rect 154777 101147 154811 101175
rect 154839 101147 154887 101175
rect 154577 101113 154887 101147
rect 154577 101085 154625 101113
rect 154653 101085 154687 101113
rect 154715 101085 154749 101113
rect 154777 101085 154811 101113
rect 154839 101085 154887 101113
rect 154577 101051 154887 101085
rect 154577 101023 154625 101051
rect 154653 101023 154687 101051
rect 154715 101023 154749 101051
rect 154777 101023 154811 101051
rect 154839 101023 154887 101051
rect 154577 100989 154887 101023
rect 154577 100961 154625 100989
rect 154653 100961 154687 100989
rect 154715 100961 154749 100989
rect 154777 100961 154811 100989
rect 154839 100961 154887 100989
rect 154577 92175 154887 100961
rect 154577 92147 154625 92175
rect 154653 92147 154687 92175
rect 154715 92147 154749 92175
rect 154777 92147 154811 92175
rect 154839 92147 154887 92175
rect 154577 92113 154887 92147
rect 154577 92085 154625 92113
rect 154653 92085 154687 92113
rect 154715 92085 154749 92113
rect 154777 92085 154811 92113
rect 154839 92085 154887 92113
rect 154577 92051 154887 92085
rect 154577 92023 154625 92051
rect 154653 92023 154687 92051
rect 154715 92023 154749 92051
rect 154777 92023 154811 92051
rect 154839 92023 154887 92051
rect 154577 91989 154887 92023
rect 154577 91961 154625 91989
rect 154653 91961 154687 91989
rect 154715 91961 154749 91989
rect 154777 91961 154811 91989
rect 154839 91961 154887 91989
rect 154577 83175 154887 91961
rect 154577 83147 154625 83175
rect 154653 83147 154687 83175
rect 154715 83147 154749 83175
rect 154777 83147 154811 83175
rect 154839 83147 154887 83175
rect 154577 83113 154887 83147
rect 154577 83085 154625 83113
rect 154653 83085 154687 83113
rect 154715 83085 154749 83113
rect 154777 83085 154811 83113
rect 154839 83085 154887 83113
rect 154577 83051 154887 83085
rect 154577 83023 154625 83051
rect 154653 83023 154687 83051
rect 154715 83023 154749 83051
rect 154777 83023 154811 83051
rect 154839 83023 154887 83051
rect 154577 82989 154887 83023
rect 154577 82961 154625 82989
rect 154653 82961 154687 82989
rect 154715 82961 154749 82989
rect 154777 82961 154811 82989
rect 154839 82961 154887 82989
rect 154577 74175 154887 82961
rect 154577 74147 154625 74175
rect 154653 74147 154687 74175
rect 154715 74147 154749 74175
rect 154777 74147 154811 74175
rect 154839 74147 154887 74175
rect 154577 74113 154887 74147
rect 154577 74085 154625 74113
rect 154653 74085 154687 74113
rect 154715 74085 154749 74113
rect 154777 74085 154811 74113
rect 154839 74085 154887 74113
rect 154577 74051 154887 74085
rect 154577 74023 154625 74051
rect 154653 74023 154687 74051
rect 154715 74023 154749 74051
rect 154777 74023 154811 74051
rect 154839 74023 154887 74051
rect 154577 73989 154887 74023
rect 154577 73961 154625 73989
rect 154653 73961 154687 73989
rect 154715 73961 154749 73989
rect 154777 73961 154811 73989
rect 154839 73961 154887 73989
rect 154577 65175 154887 73961
rect 154577 65147 154625 65175
rect 154653 65147 154687 65175
rect 154715 65147 154749 65175
rect 154777 65147 154811 65175
rect 154839 65147 154887 65175
rect 154577 65113 154887 65147
rect 154577 65085 154625 65113
rect 154653 65085 154687 65113
rect 154715 65085 154749 65113
rect 154777 65085 154811 65113
rect 154839 65085 154887 65113
rect 154577 65051 154887 65085
rect 154577 65023 154625 65051
rect 154653 65023 154687 65051
rect 154715 65023 154749 65051
rect 154777 65023 154811 65051
rect 154839 65023 154887 65051
rect 154577 64989 154887 65023
rect 154577 64961 154625 64989
rect 154653 64961 154687 64989
rect 154715 64961 154749 64989
rect 154777 64961 154811 64989
rect 154839 64961 154887 64989
rect 154577 56175 154887 64961
rect 154577 56147 154625 56175
rect 154653 56147 154687 56175
rect 154715 56147 154749 56175
rect 154777 56147 154811 56175
rect 154839 56147 154887 56175
rect 154577 56113 154887 56147
rect 154577 56085 154625 56113
rect 154653 56085 154687 56113
rect 154715 56085 154749 56113
rect 154777 56085 154811 56113
rect 154839 56085 154887 56113
rect 154577 56051 154887 56085
rect 154577 56023 154625 56051
rect 154653 56023 154687 56051
rect 154715 56023 154749 56051
rect 154777 56023 154811 56051
rect 154839 56023 154887 56051
rect 154577 55989 154887 56023
rect 154577 55961 154625 55989
rect 154653 55961 154687 55989
rect 154715 55961 154749 55989
rect 154777 55961 154811 55989
rect 154839 55961 154887 55989
rect 154577 47175 154887 55961
rect 154577 47147 154625 47175
rect 154653 47147 154687 47175
rect 154715 47147 154749 47175
rect 154777 47147 154811 47175
rect 154839 47147 154887 47175
rect 154577 47113 154887 47147
rect 154577 47085 154625 47113
rect 154653 47085 154687 47113
rect 154715 47085 154749 47113
rect 154777 47085 154811 47113
rect 154839 47085 154887 47113
rect 154577 47051 154887 47085
rect 154577 47023 154625 47051
rect 154653 47023 154687 47051
rect 154715 47023 154749 47051
rect 154777 47023 154811 47051
rect 154839 47023 154887 47051
rect 154577 46989 154887 47023
rect 154577 46961 154625 46989
rect 154653 46961 154687 46989
rect 154715 46961 154749 46989
rect 154777 46961 154811 46989
rect 154839 46961 154887 46989
rect 154577 38175 154887 46961
rect 154577 38147 154625 38175
rect 154653 38147 154687 38175
rect 154715 38147 154749 38175
rect 154777 38147 154811 38175
rect 154839 38147 154887 38175
rect 154577 38113 154887 38147
rect 154577 38085 154625 38113
rect 154653 38085 154687 38113
rect 154715 38085 154749 38113
rect 154777 38085 154811 38113
rect 154839 38085 154887 38113
rect 154577 38051 154887 38085
rect 154577 38023 154625 38051
rect 154653 38023 154687 38051
rect 154715 38023 154749 38051
rect 154777 38023 154811 38051
rect 154839 38023 154887 38051
rect 154577 37989 154887 38023
rect 154577 37961 154625 37989
rect 154653 37961 154687 37989
rect 154715 37961 154749 37989
rect 154777 37961 154811 37989
rect 154839 37961 154887 37989
rect 154577 29175 154887 37961
rect 154577 29147 154625 29175
rect 154653 29147 154687 29175
rect 154715 29147 154749 29175
rect 154777 29147 154811 29175
rect 154839 29147 154887 29175
rect 154577 29113 154887 29147
rect 154577 29085 154625 29113
rect 154653 29085 154687 29113
rect 154715 29085 154749 29113
rect 154777 29085 154811 29113
rect 154839 29085 154887 29113
rect 154577 29051 154887 29085
rect 154577 29023 154625 29051
rect 154653 29023 154687 29051
rect 154715 29023 154749 29051
rect 154777 29023 154811 29051
rect 154839 29023 154887 29051
rect 154577 28989 154887 29023
rect 154577 28961 154625 28989
rect 154653 28961 154687 28989
rect 154715 28961 154749 28989
rect 154777 28961 154811 28989
rect 154839 28961 154887 28989
rect 154577 20175 154887 28961
rect 154577 20147 154625 20175
rect 154653 20147 154687 20175
rect 154715 20147 154749 20175
rect 154777 20147 154811 20175
rect 154839 20147 154887 20175
rect 154577 20113 154887 20147
rect 154577 20085 154625 20113
rect 154653 20085 154687 20113
rect 154715 20085 154749 20113
rect 154777 20085 154811 20113
rect 154839 20085 154887 20113
rect 154577 20051 154887 20085
rect 154577 20023 154625 20051
rect 154653 20023 154687 20051
rect 154715 20023 154749 20051
rect 154777 20023 154811 20051
rect 154839 20023 154887 20051
rect 154577 19989 154887 20023
rect 154577 19961 154625 19989
rect 154653 19961 154687 19989
rect 154715 19961 154749 19989
rect 154777 19961 154811 19989
rect 154839 19961 154887 19989
rect 154577 11175 154887 19961
rect 154577 11147 154625 11175
rect 154653 11147 154687 11175
rect 154715 11147 154749 11175
rect 154777 11147 154811 11175
rect 154839 11147 154887 11175
rect 154577 11113 154887 11147
rect 154577 11085 154625 11113
rect 154653 11085 154687 11113
rect 154715 11085 154749 11113
rect 154777 11085 154811 11113
rect 154839 11085 154887 11113
rect 154577 11051 154887 11085
rect 154577 11023 154625 11051
rect 154653 11023 154687 11051
rect 154715 11023 154749 11051
rect 154777 11023 154811 11051
rect 154839 11023 154887 11051
rect 154577 10989 154887 11023
rect 154577 10961 154625 10989
rect 154653 10961 154687 10989
rect 154715 10961 154749 10989
rect 154777 10961 154811 10989
rect 154839 10961 154887 10989
rect 154577 2175 154887 10961
rect 154577 2147 154625 2175
rect 154653 2147 154687 2175
rect 154715 2147 154749 2175
rect 154777 2147 154811 2175
rect 154839 2147 154887 2175
rect 154577 2113 154887 2147
rect 154577 2085 154625 2113
rect 154653 2085 154687 2113
rect 154715 2085 154749 2113
rect 154777 2085 154811 2113
rect 154839 2085 154887 2113
rect 154577 2051 154887 2085
rect 154577 2023 154625 2051
rect 154653 2023 154687 2051
rect 154715 2023 154749 2051
rect 154777 2023 154811 2051
rect 154839 2023 154887 2051
rect 154577 1989 154887 2023
rect 154577 1961 154625 1989
rect 154653 1961 154687 1989
rect 154715 1961 154749 1989
rect 154777 1961 154811 1989
rect 154839 1961 154887 1989
rect 154577 -80 154887 1961
rect 154577 -108 154625 -80
rect 154653 -108 154687 -80
rect 154715 -108 154749 -80
rect 154777 -108 154811 -80
rect 154839 -108 154887 -80
rect 154577 -142 154887 -108
rect 154577 -170 154625 -142
rect 154653 -170 154687 -142
rect 154715 -170 154749 -142
rect 154777 -170 154811 -142
rect 154839 -170 154887 -142
rect 154577 -204 154887 -170
rect 154577 -232 154625 -204
rect 154653 -232 154687 -204
rect 154715 -232 154749 -204
rect 154777 -232 154811 -204
rect 154839 -232 154887 -204
rect 154577 -266 154887 -232
rect 154577 -294 154625 -266
rect 154653 -294 154687 -266
rect 154715 -294 154749 -266
rect 154777 -294 154811 -266
rect 154839 -294 154887 -266
rect 154577 -822 154887 -294
rect 156437 299086 156747 299134
rect 156437 299058 156485 299086
rect 156513 299058 156547 299086
rect 156575 299058 156609 299086
rect 156637 299058 156671 299086
rect 156699 299058 156747 299086
rect 156437 299024 156747 299058
rect 156437 298996 156485 299024
rect 156513 298996 156547 299024
rect 156575 298996 156609 299024
rect 156637 298996 156671 299024
rect 156699 298996 156747 299024
rect 156437 298962 156747 298996
rect 156437 298934 156485 298962
rect 156513 298934 156547 298962
rect 156575 298934 156609 298962
rect 156637 298934 156671 298962
rect 156699 298934 156747 298962
rect 156437 298900 156747 298934
rect 156437 298872 156485 298900
rect 156513 298872 156547 298900
rect 156575 298872 156609 298900
rect 156637 298872 156671 298900
rect 156699 298872 156747 298900
rect 156437 293175 156747 298872
rect 156437 293147 156485 293175
rect 156513 293147 156547 293175
rect 156575 293147 156609 293175
rect 156637 293147 156671 293175
rect 156699 293147 156747 293175
rect 156437 293113 156747 293147
rect 156437 293085 156485 293113
rect 156513 293085 156547 293113
rect 156575 293085 156609 293113
rect 156637 293085 156671 293113
rect 156699 293085 156747 293113
rect 156437 293051 156747 293085
rect 156437 293023 156485 293051
rect 156513 293023 156547 293051
rect 156575 293023 156609 293051
rect 156637 293023 156671 293051
rect 156699 293023 156747 293051
rect 156437 292989 156747 293023
rect 156437 292961 156485 292989
rect 156513 292961 156547 292989
rect 156575 292961 156609 292989
rect 156637 292961 156671 292989
rect 156699 292961 156747 292989
rect 156437 284175 156747 292961
rect 156437 284147 156485 284175
rect 156513 284147 156547 284175
rect 156575 284147 156609 284175
rect 156637 284147 156671 284175
rect 156699 284147 156747 284175
rect 156437 284113 156747 284147
rect 156437 284085 156485 284113
rect 156513 284085 156547 284113
rect 156575 284085 156609 284113
rect 156637 284085 156671 284113
rect 156699 284085 156747 284113
rect 156437 284051 156747 284085
rect 156437 284023 156485 284051
rect 156513 284023 156547 284051
rect 156575 284023 156609 284051
rect 156637 284023 156671 284051
rect 156699 284023 156747 284051
rect 156437 283989 156747 284023
rect 156437 283961 156485 283989
rect 156513 283961 156547 283989
rect 156575 283961 156609 283989
rect 156637 283961 156671 283989
rect 156699 283961 156747 283989
rect 156437 275175 156747 283961
rect 156437 275147 156485 275175
rect 156513 275147 156547 275175
rect 156575 275147 156609 275175
rect 156637 275147 156671 275175
rect 156699 275147 156747 275175
rect 156437 275113 156747 275147
rect 156437 275085 156485 275113
rect 156513 275085 156547 275113
rect 156575 275085 156609 275113
rect 156637 275085 156671 275113
rect 156699 275085 156747 275113
rect 156437 275051 156747 275085
rect 156437 275023 156485 275051
rect 156513 275023 156547 275051
rect 156575 275023 156609 275051
rect 156637 275023 156671 275051
rect 156699 275023 156747 275051
rect 156437 274989 156747 275023
rect 156437 274961 156485 274989
rect 156513 274961 156547 274989
rect 156575 274961 156609 274989
rect 156637 274961 156671 274989
rect 156699 274961 156747 274989
rect 156437 266175 156747 274961
rect 156437 266147 156485 266175
rect 156513 266147 156547 266175
rect 156575 266147 156609 266175
rect 156637 266147 156671 266175
rect 156699 266147 156747 266175
rect 156437 266113 156747 266147
rect 156437 266085 156485 266113
rect 156513 266085 156547 266113
rect 156575 266085 156609 266113
rect 156637 266085 156671 266113
rect 156699 266085 156747 266113
rect 156437 266051 156747 266085
rect 156437 266023 156485 266051
rect 156513 266023 156547 266051
rect 156575 266023 156609 266051
rect 156637 266023 156671 266051
rect 156699 266023 156747 266051
rect 156437 265989 156747 266023
rect 156437 265961 156485 265989
rect 156513 265961 156547 265989
rect 156575 265961 156609 265989
rect 156637 265961 156671 265989
rect 156699 265961 156747 265989
rect 156437 257175 156747 265961
rect 156437 257147 156485 257175
rect 156513 257147 156547 257175
rect 156575 257147 156609 257175
rect 156637 257147 156671 257175
rect 156699 257147 156747 257175
rect 156437 257113 156747 257147
rect 156437 257085 156485 257113
rect 156513 257085 156547 257113
rect 156575 257085 156609 257113
rect 156637 257085 156671 257113
rect 156699 257085 156747 257113
rect 156437 257051 156747 257085
rect 156437 257023 156485 257051
rect 156513 257023 156547 257051
rect 156575 257023 156609 257051
rect 156637 257023 156671 257051
rect 156699 257023 156747 257051
rect 156437 256989 156747 257023
rect 156437 256961 156485 256989
rect 156513 256961 156547 256989
rect 156575 256961 156609 256989
rect 156637 256961 156671 256989
rect 156699 256961 156747 256989
rect 156437 248175 156747 256961
rect 156437 248147 156485 248175
rect 156513 248147 156547 248175
rect 156575 248147 156609 248175
rect 156637 248147 156671 248175
rect 156699 248147 156747 248175
rect 156437 248113 156747 248147
rect 156437 248085 156485 248113
rect 156513 248085 156547 248113
rect 156575 248085 156609 248113
rect 156637 248085 156671 248113
rect 156699 248085 156747 248113
rect 156437 248051 156747 248085
rect 156437 248023 156485 248051
rect 156513 248023 156547 248051
rect 156575 248023 156609 248051
rect 156637 248023 156671 248051
rect 156699 248023 156747 248051
rect 156437 247989 156747 248023
rect 156437 247961 156485 247989
rect 156513 247961 156547 247989
rect 156575 247961 156609 247989
rect 156637 247961 156671 247989
rect 156699 247961 156747 247989
rect 156437 239175 156747 247961
rect 156437 239147 156485 239175
rect 156513 239147 156547 239175
rect 156575 239147 156609 239175
rect 156637 239147 156671 239175
rect 156699 239147 156747 239175
rect 156437 239113 156747 239147
rect 156437 239085 156485 239113
rect 156513 239085 156547 239113
rect 156575 239085 156609 239113
rect 156637 239085 156671 239113
rect 156699 239085 156747 239113
rect 156437 239051 156747 239085
rect 156437 239023 156485 239051
rect 156513 239023 156547 239051
rect 156575 239023 156609 239051
rect 156637 239023 156671 239051
rect 156699 239023 156747 239051
rect 156437 238989 156747 239023
rect 156437 238961 156485 238989
rect 156513 238961 156547 238989
rect 156575 238961 156609 238989
rect 156637 238961 156671 238989
rect 156699 238961 156747 238989
rect 156437 230175 156747 238961
rect 156437 230147 156485 230175
rect 156513 230147 156547 230175
rect 156575 230147 156609 230175
rect 156637 230147 156671 230175
rect 156699 230147 156747 230175
rect 156437 230113 156747 230147
rect 156437 230085 156485 230113
rect 156513 230085 156547 230113
rect 156575 230085 156609 230113
rect 156637 230085 156671 230113
rect 156699 230085 156747 230113
rect 156437 230051 156747 230085
rect 156437 230023 156485 230051
rect 156513 230023 156547 230051
rect 156575 230023 156609 230051
rect 156637 230023 156671 230051
rect 156699 230023 156747 230051
rect 156437 229989 156747 230023
rect 156437 229961 156485 229989
rect 156513 229961 156547 229989
rect 156575 229961 156609 229989
rect 156637 229961 156671 229989
rect 156699 229961 156747 229989
rect 156437 221175 156747 229961
rect 156437 221147 156485 221175
rect 156513 221147 156547 221175
rect 156575 221147 156609 221175
rect 156637 221147 156671 221175
rect 156699 221147 156747 221175
rect 156437 221113 156747 221147
rect 156437 221085 156485 221113
rect 156513 221085 156547 221113
rect 156575 221085 156609 221113
rect 156637 221085 156671 221113
rect 156699 221085 156747 221113
rect 156437 221051 156747 221085
rect 156437 221023 156485 221051
rect 156513 221023 156547 221051
rect 156575 221023 156609 221051
rect 156637 221023 156671 221051
rect 156699 221023 156747 221051
rect 156437 220989 156747 221023
rect 156437 220961 156485 220989
rect 156513 220961 156547 220989
rect 156575 220961 156609 220989
rect 156637 220961 156671 220989
rect 156699 220961 156747 220989
rect 156437 212175 156747 220961
rect 156437 212147 156485 212175
rect 156513 212147 156547 212175
rect 156575 212147 156609 212175
rect 156637 212147 156671 212175
rect 156699 212147 156747 212175
rect 156437 212113 156747 212147
rect 156437 212085 156485 212113
rect 156513 212085 156547 212113
rect 156575 212085 156609 212113
rect 156637 212085 156671 212113
rect 156699 212085 156747 212113
rect 156437 212051 156747 212085
rect 156437 212023 156485 212051
rect 156513 212023 156547 212051
rect 156575 212023 156609 212051
rect 156637 212023 156671 212051
rect 156699 212023 156747 212051
rect 156437 211989 156747 212023
rect 156437 211961 156485 211989
rect 156513 211961 156547 211989
rect 156575 211961 156609 211989
rect 156637 211961 156671 211989
rect 156699 211961 156747 211989
rect 156437 203175 156747 211961
rect 156437 203147 156485 203175
rect 156513 203147 156547 203175
rect 156575 203147 156609 203175
rect 156637 203147 156671 203175
rect 156699 203147 156747 203175
rect 156437 203113 156747 203147
rect 156437 203085 156485 203113
rect 156513 203085 156547 203113
rect 156575 203085 156609 203113
rect 156637 203085 156671 203113
rect 156699 203085 156747 203113
rect 156437 203051 156747 203085
rect 156437 203023 156485 203051
rect 156513 203023 156547 203051
rect 156575 203023 156609 203051
rect 156637 203023 156671 203051
rect 156699 203023 156747 203051
rect 156437 202989 156747 203023
rect 156437 202961 156485 202989
rect 156513 202961 156547 202989
rect 156575 202961 156609 202989
rect 156637 202961 156671 202989
rect 156699 202961 156747 202989
rect 156437 194175 156747 202961
rect 156437 194147 156485 194175
rect 156513 194147 156547 194175
rect 156575 194147 156609 194175
rect 156637 194147 156671 194175
rect 156699 194147 156747 194175
rect 156437 194113 156747 194147
rect 156437 194085 156485 194113
rect 156513 194085 156547 194113
rect 156575 194085 156609 194113
rect 156637 194085 156671 194113
rect 156699 194085 156747 194113
rect 156437 194051 156747 194085
rect 156437 194023 156485 194051
rect 156513 194023 156547 194051
rect 156575 194023 156609 194051
rect 156637 194023 156671 194051
rect 156699 194023 156747 194051
rect 156437 193989 156747 194023
rect 156437 193961 156485 193989
rect 156513 193961 156547 193989
rect 156575 193961 156609 193989
rect 156637 193961 156671 193989
rect 156699 193961 156747 193989
rect 156437 185175 156747 193961
rect 156437 185147 156485 185175
rect 156513 185147 156547 185175
rect 156575 185147 156609 185175
rect 156637 185147 156671 185175
rect 156699 185147 156747 185175
rect 156437 185113 156747 185147
rect 156437 185085 156485 185113
rect 156513 185085 156547 185113
rect 156575 185085 156609 185113
rect 156637 185085 156671 185113
rect 156699 185085 156747 185113
rect 156437 185051 156747 185085
rect 156437 185023 156485 185051
rect 156513 185023 156547 185051
rect 156575 185023 156609 185051
rect 156637 185023 156671 185051
rect 156699 185023 156747 185051
rect 156437 184989 156747 185023
rect 156437 184961 156485 184989
rect 156513 184961 156547 184989
rect 156575 184961 156609 184989
rect 156637 184961 156671 184989
rect 156699 184961 156747 184989
rect 156437 176175 156747 184961
rect 156437 176147 156485 176175
rect 156513 176147 156547 176175
rect 156575 176147 156609 176175
rect 156637 176147 156671 176175
rect 156699 176147 156747 176175
rect 156437 176113 156747 176147
rect 156437 176085 156485 176113
rect 156513 176085 156547 176113
rect 156575 176085 156609 176113
rect 156637 176085 156671 176113
rect 156699 176085 156747 176113
rect 156437 176051 156747 176085
rect 156437 176023 156485 176051
rect 156513 176023 156547 176051
rect 156575 176023 156609 176051
rect 156637 176023 156671 176051
rect 156699 176023 156747 176051
rect 156437 175989 156747 176023
rect 156437 175961 156485 175989
rect 156513 175961 156547 175989
rect 156575 175961 156609 175989
rect 156637 175961 156671 175989
rect 156699 175961 156747 175989
rect 156437 167175 156747 175961
rect 156437 167147 156485 167175
rect 156513 167147 156547 167175
rect 156575 167147 156609 167175
rect 156637 167147 156671 167175
rect 156699 167147 156747 167175
rect 156437 167113 156747 167147
rect 156437 167085 156485 167113
rect 156513 167085 156547 167113
rect 156575 167085 156609 167113
rect 156637 167085 156671 167113
rect 156699 167085 156747 167113
rect 156437 167051 156747 167085
rect 156437 167023 156485 167051
rect 156513 167023 156547 167051
rect 156575 167023 156609 167051
rect 156637 167023 156671 167051
rect 156699 167023 156747 167051
rect 156437 166989 156747 167023
rect 156437 166961 156485 166989
rect 156513 166961 156547 166989
rect 156575 166961 156609 166989
rect 156637 166961 156671 166989
rect 156699 166961 156747 166989
rect 156437 158175 156747 166961
rect 156437 158147 156485 158175
rect 156513 158147 156547 158175
rect 156575 158147 156609 158175
rect 156637 158147 156671 158175
rect 156699 158147 156747 158175
rect 156437 158113 156747 158147
rect 156437 158085 156485 158113
rect 156513 158085 156547 158113
rect 156575 158085 156609 158113
rect 156637 158085 156671 158113
rect 156699 158085 156747 158113
rect 156437 158051 156747 158085
rect 156437 158023 156485 158051
rect 156513 158023 156547 158051
rect 156575 158023 156609 158051
rect 156637 158023 156671 158051
rect 156699 158023 156747 158051
rect 156437 157989 156747 158023
rect 156437 157961 156485 157989
rect 156513 157961 156547 157989
rect 156575 157961 156609 157989
rect 156637 157961 156671 157989
rect 156699 157961 156747 157989
rect 156437 149175 156747 157961
rect 156437 149147 156485 149175
rect 156513 149147 156547 149175
rect 156575 149147 156609 149175
rect 156637 149147 156671 149175
rect 156699 149147 156747 149175
rect 156437 149113 156747 149147
rect 156437 149085 156485 149113
rect 156513 149085 156547 149113
rect 156575 149085 156609 149113
rect 156637 149085 156671 149113
rect 156699 149085 156747 149113
rect 156437 149051 156747 149085
rect 156437 149023 156485 149051
rect 156513 149023 156547 149051
rect 156575 149023 156609 149051
rect 156637 149023 156671 149051
rect 156699 149023 156747 149051
rect 156437 148989 156747 149023
rect 156437 148961 156485 148989
rect 156513 148961 156547 148989
rect 156575 148961 156609 148989
rect 156637 148961 156671 148989
rect 156699 148961 156747 148989
rect 156437 140175 156747 148961
rect 156437 140147 156485 140175
rect 156513 140147 156547 140175
rect 156575 140147 156609 140175
rect 156637 140147 156671 140175
rect 156699 140147 156747 140175
rect 156437 140113 156747 140147
rect 156437 140085 156485 140113
rect 156513 140085 156547 140113
rect 156575 140085 156609 140113
rect 156637 140085 156671 140113
rect 156699 140085 156747 140113
rect 156437 140051 156747 140085
rect 156437 140023 156485 140051
rect 156513 140023 156547 140051
rect 156575 140023 156609 140051
rect 156637 140023 156671 140051
rect 156699 140023 156747 140051
rect 156437 139989 156747 140023
rect 156437 139961 156485 139989
rect 156513 139961 156547 139989
rect 156575 139961 156609 139989
rect 156637 139961 156671 139989
rect 156699 139961 156747 139989
rect 156437 131175 156747 139961
rect 156437 131147 156485 131175
rect 156513 131147 156547 131175
rect 156575 131147 156609 131175
rect 156637 131147 156671 131175
rect 156699 131147 156747 131175
rect 156437 131113 156747 131147
rect 156437 131085 156485 131113
rect 156513 131085 156547 131113
rect 156575 131085 156609 131113
rect 156637 131085 156671 131113
rect 156699 131085 156747 131113
rect 156437 131051 156747 131085
rect 156437 131023 156485 131051
rect 156513 131023 156547 131051
rect 156575 131023 156609 131051
rect 156637 131023 156671 131051
rect 156699 131023 156747 131051
rect 156437 130989 156747 131023
rect 156437 130961 156485 130989
rect 156513 130961 156547 130989
rect 156575 130961 156609 130989
rect 156637 130961 156671 130989
rect 156699 130961 156747 130989
rect 156437 122175 156747 130961
rect 156437 122147 156485 122175
rect 156513 122147 156547 122175
rect 156575 122147 156609 122175
rect 156637 122147 156671 122175
rect 156699 122147 156747 122175
rect 156437 122113 156747 122147
rect 156437 122085 156485 122113
rect 156513 122085 156547 122113
rect 156575 122085 156609 122113
rect 156637 122085 156671 122113
rect 156699 122085 156747 122113
rect 156437 122051 156747 122085
rect 156437 122023 156485 122051
rect 156513 122023 156547 122051
rect 156575 122023 156609 122051
rect 156637 122023 156671 122051
rect 156699 122023 156747 122051
rect 156437 121989 156747 122023
rect 156437 121961 156485 121989
rect 156513 121961 156547 121989
rect 156575 121961 156609 121989
rect 156637 121961 156671 121989
rect 156699 121961 156747 121989
rect 156437 113175 156747 121961
rect 156437 113147 156485 113175
rect 156513 113147 156547 113175
rect 156575 113147 156609 113175
rect 156637 113147 156671 113175
rect 156699 113147 156747 113175
rect 156437 113113 156747 113147
rect 156437 113085 156485 113113
rect 156513 113085 156547 113113
rect 156575 113085 156609 113113
rect 156637 113085 156671 113113
rect 156699 113085 156747 113113
rect 156437 113051 156747 113085
rect 156437 113023 156485 113051
rect 156513 113023 156547 113051
rect 156575 113023 156609 113051
rect 156637 113023 156671 113051
rect 156699 113023 156747 113051
rect 156437 112989 156747 113023
rect 156437 112961 156485 112989
rect 156513 112961 156547 112989
rect 156575 112961 156609 112989
rect 156637 112961 156671 112989
rect 156699 112961 156747 112989
rect 156437 104175 156747 112961
rect 156437 104147 156485 104175
rect 156513 104147 156547 104175
rect 156575 104147 156609 104175
rect 156637 104147 156671 104175
rect 156699 104147 156747 104175
rect 156437 104113 156747 104147
rect 156437 104085 156485 104113
rect 156513 104085 156547 104113
rect 156575 104085 156609 104113
rect 156637 104085 156671 104113
rect 156699 104085 156747 104113
rect 156437 104051 156747 104085
rect 156437 104023 156485 104051
rect 156513 104023 156547 104051
rect 156575 104023 156609 104051
rect 156637 104023 156671 104051
rect 156699 104023 156747 104051
rect 156437 103989 156747 104023
rect 156437 103961 156485 103989
rect 156513 103961 156547 103989
rect 156575 103961 156609 103989
rect 156637 103961 156671 103989
rect 156699 103961 156747 103989
rect 156437 95175 156747 103961
rect 156437 95147 156485 95175
rect 156513 95147 156547 95175
rect 156575 95147 156609 95175
rect 156637 95147 156671 95175
rect 156699 95147 156747 95175
rect 156437 95113 156747 95147
rect 156437 95085 156485 95113
rect 156513 95085 156547 95113
rect 156575 95085 156609 95113
rect 156637 95085 156671 95113
rect 156699 95085 156747 95113
rect 156437 95051 156747 95085
rect 156437 95023 156485 95051
rect 156513 95023 156547 95051
rect 156575 95023 156609 95051
rect 156637 95023 156671 95051
rect 156699 95023 156747 95051
rect 156437 94989 156747 95023
rect 156437 94961 156485 94989
rect 156513 94961 156547 94989
rect 156575 94961 156609 94989
rect 156637 94961 156671 94989
rect 156699 94961 156747 94989
rect 156437 86175 156747 94961
rect 156437 86147 156485 86175
rect 156513 86147 156547 86175
rect 156575 86147 156609 86175
rect 156637 86147 156671 86175
rect 156699 86147 156747 86175
rect 156437 86113 156747 86147
rect 156437 86085 156485 86113
rect 156513 86085 156547 86113
rect 156575 86085 156609 86113
rect 156637 86085 156671 86113
rect 156699 86085 156747 86113
rect 156437 86051 156747 86085
rect 156437 86023 156485 86051
rect 156513 86023 156547 86051
rect 156575 86023 156609 86051
rect 156637 86023 156671 86051
rect 156699 86023 156747 86051
rect 156437 85989 156747 86023
rect 156437 85961 156485 85989
rect 156513 85961 156547 85989
rect 156575 85961 156609 85989
rect 156637 85961 156671 85989
rect 156699 85961 156747 85989
rect 156437 77175 156747 85961
rect 156437 77147 156485 77175
rect 156513 77147 156547 77175
rect 156575 77147 156609 77175
rect 156637 77147 156671 77175
rect 156699 77147 156747 77175
rect 156437 77113 156747 77147
rect 156437 77085 156485 77113
rect 156513 77085 156547 77113
rect 156575 77085 156609 77113
rect 156637 77085 156671 77113
rect 156699 77085 156747 77113
rect 156437 77051 156747 77085
rect 156437 77023 156485 77051
rect 156513 77023 156547 77051
rect 156575 77023 156609 77051
rect 156637 77023 156671 77051
rect 156699 77023 156747 77051
rect 156437 76989 156747 77023
rect 156437 76961 156485 76989
rect 156513 76961 156547 76989
rect 156575 76961 156609 76989
rect 156637 76961 156671 76989
rect 156699 76961 156747 76989
rect 156437 68175 156747 76961
rect 156437 68147 156485 68175
rect 156513 68147 156547 68175
rect 156575 68147 156609 68175
rect 156637 68147 156671 68175
rect 156699 68147 156747 68175
rect 156437 68113 156747 68147
rect 156437 68085 156485 68113
rect 156513 68085 156547 68113
rect 156575 68085 156609 68113
rect 156637 68085 156671 68113
rect 156699 68085 156747 68113
rect 156437 68051 156747 68085
rect 156437 68023 156485 68051
rect 156513 68023 156547 68051
rect 156575 68023 156609 68051
rect 156637 68023 156671 68051
rect 156699 68023 156747 68051
rect 156437 67989 156747 68023
rect 156437 67961 156485 67989
rect 156513 67961 156547 67989
rect 156575 67961 156609 67989
rect 156637 67961 156671 67989
rect 156699 67961 156747 67989
rect 156437 59175 156747 67961
rect 156437 59147 156485 59175
rect 156513 59147 156547 59175
rect 156575 59147 156609 59175
rect 156637 59147 156671 59175
rect 156699 59147 156747 59175
rect 156437 59113 156747 59147
rect 156437 59085 156485 59113
rect 156513 59085 156547 59113
rect 156575 59085 156609 59113
rect 156637 59085 156671 59113
rect 156699 59085 156747 59113
rect 156437 59051 156747 59085
rect 156437 59023 156485 59051
rect 156513 59023 156547 59051
rect 156575 59023 156609 59051
rect 156637 59023 156671 59051
rect 156699 59023 156747 59051
rect 156437 58989 156747 59023
rect 156437 58961 156485 58989
rect 156513 58961 156547 58989
rect 156575 58961 156609 58989
rect 156637 58961 156671 58989
rect 156699 58961 156747 58989
rect 156437 50175 156747 58961
rect 156437 50147 156485 50175
rect 156513 50147 156547 50175
rect 156575 50147 156609 50175
rect 156637 50147 156671 50175
rect 156699 50147 156747 50175
rect 156437 50113 156747 50147
rect 156437 50085 156485 50113
rect 156513 50085 156547 50113
rect 156575 50085 156609 50113
rect 156637 50085 156671 50113
rect 156699 50085 156747 50113
rect 156437 50051 156747 50085
rect 156437 50023 156485 50051
rect 156513 50023 156547 50051
rect 156575 50023 156609 50051
rect 156637 50023 156671 50051
rect 156699 50023 156747 50051
rect 156437 49989 156747 50023
rect 156437 49961 156485 49989
rect 156513 49961 156547 49989
rect 156575 49961 156609 49989
rect 156637 49961 156671 49989
rect 156699 49961 156747 49989
rect 156437 41175 156747 49961
rect 156437 41147 156485 41175
rect 156513 41147 156547 41175
rect 156575 41147 156609 41175
rect 156637 41147 156671 41175
rect 156699 41147 156747 41175
rect 156437 41113 156747 41147
rect 156437 41085 156485 41113
rect 156513 41085 156547 41113
rect 156575 41085 156609 41113
rect 156637 41085 156671 41113
rect 156699 41085 156747 41113
rect 156437 41051 156747 41085
rect 156437 41023 156485 41051
rect 156513 41023 156547 41051
rect 156575 41023 156609 41051
rect 156637 41023 156671 41051
rect 156699 41023 156747 41051
rect 156437 40989 156747 41023
rect 156437 40961 156485 40989
rect 156513 40961 156547 40989
rect 156575 40961 156609 40989
rect 156637 40961 156671 40989
rect 156699 40961 156747 40989
rect 156437 32175 156747 40961
rect 156437 32147 156485 32175
rect 156513 32147 156547 32175
rect 156575 32147 156609 32175
rect 156637 32147 156671 32175
rect 156699 32147 156747 32175
rect 156437 32113 156747 32147
rect 156437 32085 156485 32113
rect 156513 32085 156547 32113
rect 156575 32085 156609 32113
rect 156637 32085 156671 32113
rect 156699 32085 156747 32113
rect 156437 32051 156747 32085
rect 156437 32023 156485 32051
rect 156513 32023 156547 32051
rect 156575 32023 156609 32051
rect 156637 32023 156671 32051
rect 156699 32023 156747 32051
rect 156437 31989 156747 32023
rect 156437 31961 156485 31989
rect 156513 31961 156547 31989
rect 156575 31961 156609 31989
rect 156637 31961 156671 31989
rect 156699 31961 156747 31989
rect 156437 23175 156747 31961
rect 156437 23147 156485 23175
rect 156513 23147 156547 23175
rect 156575 23147 156609 23175
rect 156637 23147 156671 23175
rect 156699 23147 156747 23175
rect 156437 23113 156747 23147
rect 156437 23085 156485 23113
rect 156513 23085 156547 23113
rect 156575 23085 156609 23113
rect 156637 23085 156671 23113
rect 156699 23085 156747 23113
rect 156437 23051 156747 23085
rect 156437 23023 156485 23051
rect 156513 23023 156547 23051
rect 156575 23023 156609 23051
rect 156637 23023 156671 23051
rect 156699 23023 156747 23051
rect 156437 22989 156747 23023
rect 156437 22961 156485 22989
rect 156513 22961 156547 22989
rect 156575 22961 156609 22989
rect 156637 22961 156671 22989
rect 156699 22961 156747 22989
rect 156437 14175 156747 22961
rect 156437 14147 156485 14175
rect 156513 14147 156547 14175
rect 156575 14147 156609 14175
rect 156637 14147 156671 14175
rect 156699 14147 156747 14175
rect 156437 14113 156747 14147
rect 156437 14085 156485 14113
rect 156513 14085 156547 14113
rect 156575 14085 156609 14113
rect 156637 14085 156671 14113
rect 156699 14085 156747 14113
rect 156437 14051 156747 14085
rect 156437 14023 156485 14051
rect 156513 14023 156547 14051
rect 156575 14023 156609 14051
rect 156637 14023 156671 14051
rect 156699 14023 156747 14051
rect 156437 13989 156747 14023
rect 156437 13961 156485 13989
rect 156513 13961 156547 13989
rect 156575 13961 156609 13989
rect 156637 13961 156671 13989
rect 156699 13961 156747 13989
rect 156437 5175 156747 13961
rect 156437 5147 156485 5175
rect 156513 5147 156547 5175
rect 156575 5147 156609 5175
rect 156637 5147 156671 5175
rect 156699 5147 156747 5175
rect 156437 5113 156747 5147
rect 156437 5085 156485 5113
rect 156513 5085 156547 5113
rect 156575 5085 156609 5113
rect 156637 5085 156671 5113
rect 156699 5085 156747 5113
rect 156437 5051 156747 5085
rect 156437 5023 156485 5051
rect 156513 5023 156547 5051
rect 156575 5023 156609 5051
rect 156637 5023 156671 5051
rect 156699 5023 156747 5051
rect 156437 4989 156747 5023
rect 156437 4961 156485 4989
rect 156513 4961 156547 4989
rect 156575 4961 156609 4989
rect 156637 4961 156671 4989
rect 156699 4961 156747 4989
rect 156437 -560 156747 4961
rect 156437 -588 156485 -560
rect 156513 -588 156547 -560
rect 156575 -588 156609 -560
rect 156637 -588 156671 -560
rect 156699 -588 156747 -560
rect 156437 -622 156747 -588
rect 156437 -650 156485 -622
rect 156513 -650 156547 -622
rect 156575 -650 156609 -622
rect 156637 -650 156671 -622
rect 156699 -650 156747 -622
rect 156437 -684 156747 -650
rect 156437 -712 156485 -684
rect 156513 -712 156547 -684
rect 156575 -712 156609 -684
rect 156637 -712 156671 -684
rect 156699 -712 156747 -684
rect 156437 -746 156747 -712
rect 156437 -774 156485 -746
rect 156513 -774 156547 -746
rect 156575 -774 156609 -746
rect 156637 -774 156671 -746
rect 156699 -774 156747 -746
rect 156437 -822 156747 -774
rect 163577 298606 163887 299134
rect 163577 298578 163625 298606
rect 163653 298578 163687 298606
rect 163715 298578 163749 298606
rect 163777 298578 163811 298606
rect 163839 298578 163887 298606
rect 163577 298544 163887 298578
rect 163577 298516 163625 298544
rect 163653 298516 163687 298544
rect 163715 298516 163749 298544
rect 163777 298516 163811 298544
rect 163839 298516 163887 298544
rect 163577 298482 163887 298516
rect 163577 298454 163625 298482
rect 163653 298454 163687 298482
rect 163715 298454 163749 298482
rect 163777 298454 163811 298482
rect 163839 298454 163887 298482
rect 163577 298420 163887 298454
rect 163577 298392 163625 298420
rect 163653 298392 163687 298420
rect 163715 298392 163749 298420
rect 163777 298392 163811 298420
rect 163839 298392 163887 298420
rect 163577 290175 163887 298392
rect 163577 290147 163625 290175
rect 163653 290147 163687 290175
rect 163715 290147 163749 290175
rect 163777 290147 163811 290175
rect 163839 290147 163887 290175
rect 163577 290113 163887 290147
rect 163577 290085 163625 290113
rect 163653 290085 163687 290113
rect 163715 290085 163749 290113
rect 163777 290085 163811 290113
rect 163839 290085 163887 290113
rect 163577 290051 163887 290085
rect 163577 290023 163625 290051
rect 163653 290023 163687 290051
rect 163715 290023 163749 290051
rect 163777 290023 163811 290051
rect 163839 290023 163887 290051
rect 163577 289989 163887 290023
rect 163577 289961 163625 289989
rect 163653 289961 163687 289989
rect 163715 289961 163749 289989
rect 163777 289961 163811 289989
rect 163839 289961 163887 289989
rect 163577 281175 163887 289961
rect 163577 281147 163625 281175
rect 163653 281147 163687 281175
rect 163715 281147 163749 281175
rect 163777 281147 163811 281175
rect 163839 281147 163887 281175
rect 163577 281113 163887 281147
rect 163577 281085 163625 281113
rect 163653 281085 163687 281113
rect 163715 281085 163749 281113
rect 163777 281085 163811 281113
rect 163839 281085 163887 281113
rect 163577 281051 163887 281085
rect 163577 281023 163625 281051
rect 163653 281023 163687 281051
rect 163715 281023 163749 281051
rect 163777 281023 163811 281051
rect 163839 281023 163887 281051
rect 163577 280989 163887 281023
rect 163577 280961 163625 280989
rect 163653 280961 163687 280989
rect 163715 280961 163749 280989
rect 163777 280961 163811 280989
rect 163839 280961 163887 280989
rect 163577 272175 163887 280961
rect 163577 272147 163625 272175
rect 163653 272147 163687 272175
rect 163715 272147 163749 272175
rect 163777 272147 163811 272175
rect 163839 272147 163887 272175
rect 163577 272113 163887 272147
rect 163577 272085 163625 272113
rect 163653 272085 163687 272113
rect 163715 272085 163749 272113
rect 163777 272085 163811 272113
rect 163839 272085 163887 272113
rect 163577 272051 163887 272085
rect 163577 272023 163625 272051
rect 163653 272023 163687 272051
rect 163715 272023 163749 272051
rect 163777 272023 163811 272051
rect 163839 272023 163887 272051
rect 163577 271989 163887 272023
rect 163577 271961 163625 271989
rect 163653 271961 163687 271989
rect 163715 271961 163749 271989
rect 163777 271961 163811 271989
rect 163839 271961 163887 271989
rect 163577 263175 163887 271961
rect 163577 263147 163625 263175
rect 163653 263147 163687 263175
rect 163715 263147 163749 263175
rect 163777 263147 163811 263175
rect 163839 263147 163887 263175
rect 163577 263113 163887 263147
rect 163577 263085 163625 263113
rect 163653 263085 163687 263113
rect 163715 263085 163749 263113
rect 163777 263085 163811 263113
rect 163839 263085 163887 263113
rect 163577 263051 163887 263085
rect 163577 263023 163625 263051
rect 163653 263023 163687 263051
rect 163715 263023 163749 263051
rect 163777 263023 163811 263051
rect 163839 263023 163887 263051
rect 163577 262989 163887 263023
rect 163577 262961 163625 262989
rect 163653 262961 163687 262989
rect 163715 262961 163749 262989
rect 163777 262961 163811 262989
rect 163839 262961 163887 262989
rect 163577 254175 163887 262961
rect 163577 254147 163625 254175
rect 163653 254147 163687 254175
rect 163715 254147 163749 254175
rect 163777 254147 163811 254175
rect 163839 254147 163887 254175
rect 163577 254113 163887 254147
rect 163577 254085 163625 254113
rect 163653 254085 163687 254113
rect 163715 254085 163749 254113
rect 163777 254085 163811 254113
rect 163839 254085 163887 254113
rect 163577 254051 163887 254085
rect 163577 254023 163625 254051
rect 163653 254023 163687 254051
rect 163715 254023 163749 254051
rect 163777 254023 163811 254051
rect 163839 254023 163887 254051
rect 163577 253989 163887 254023
rect 163577 253961 163625 253989
rect 163653 253961 163687 253989
rect 163715 253961 163749 253989
rect 163777 253961 163811 253989
rect 163839 253961 163887 253989
rect 163577 245175 163887 253961
rect 163577 245147 163625 245175
rect 163653 245147 163687 245175
rect 163715 245147 163749 245175
rect 163777 245147 163811 245175
rect 163839 245147 163887 245175
rect 163577 245113 163887 245147
rect 163577 245085 163625 245113
rect 163653 245085 163687 245113
rect 163715 245085 163749 245113
rect 163777 245085 163811 245113
rect 163839 245085 163887 245113
rect 163577 245051 163887 245085
rect 163577 245023 163625 245051
rect 163653 245023 163687 245051
rect 163715 245023 163749 245051
rect 163777 245023 163811 245051
rect 163839 245023 163887 245051
rect 163577 244989 163887 245023
rect 163577 244961 163625 244989
rect 163653 244961 163687 244989
rect 163715 244961 163749 244989
rect 163777 244961 163811 244989
rect 163839 244961 163887 244989
rect 163577 236175 163887 244961
rect 163577 236147 163625 236175
rect 163653 236147 163687 236175
rect 163715 236147 163749 236175
rect 163777 236147 163811 236175
rect 163839 236147 163887 236175
rect 163577 236113 163887 236147
rect 163577 236085 163625 236113
rect 163653 236085 163687 236113
rect 163715 236085 163749 236113
rect 163777 236085 163811 236113
rect 163839 236085 163887 236113
rect 163577 236051 163887 236085
rect 163577 236023 163625 236051
rect 163653 236023 163687 236051
rect 163715 236023 163749 236051
rect 163777 236023 163811 236051
rect 163839 236023 163887 236051
rect 163577 235989 163887 236023
rect 163577 235961 163625 235989
rect 163653 235961 163687 235989
rect 163715 235961 163749 235989
rect 163777 235961 163811 235989
rect 163839 235961 163887 235989
rect 163577 227175 163887 235961
rect 163577 227147 163625 227175
rect 163653 227147 163687 227175
rect 163715 227147 163749 227175
rect 163777 227147 163811 227175
rect 163839 227147 163887 227175
rect 163577 227113 163887 227147
rect 163577 227085 163625 227113
rect 163653 227085 163687 227113
rect 163715 227085 163749 227113
rect 163777 227085 163811 227113
rect 163839 227085 163887 227113
rect 163577 227051 163887 227085
rect 163577 227023 163625 227051
rect 163653 227023 163687 227051
rect 163715 227023 163749 227051
rect 163777 227023 163811 227051
rect 163839 227023 163887 227051
rect 163577 226989 163887 227023
rect 163577 226961 163625 226989
rect 163653 226961 163687 226989
rect 163715 226961 163749 226989
rect 163777 226961 163811 226989
rect 163839 226961 163887 226989
rect 163577 218175 163887 226961
rect 163577 218147 163625 218175
rect 163653 218147 163687 218175
rect 163715 218147 163749 218175
rect 163777 218147 163811 218175
rect 163839 218147 163887 218175
rect 163577 218113 163887 218147
rect 163577 218085 163625 218113
rect 163653 218085 163687 218113
rect 163715 218085 163749 218113
rect 163777 218085 163811 218113
rect 163839 218085 163887 218113
rect 163577 218051 163887 218085
rect 163577 218023 163625 218051
rect 163653 218023 163687 218051
rect 163715 218023 163749 218051
rect 163777 218023 163811 218051
rect 163839 218023 163887 218051
rect 163577 217989 163887 218023
rect 163577 217961 163625 217989
rect 163653 217961 163687 217989
rect 163715 217961 163749 217989
rect 163777 217961 163811 217989
rect 163839 217961 163887 217989
rect 163577 209175 163887 217961
rect 163577 209147 163625 209175
rect 163653 209147 163687 209175
rect 163715 209147 163749 209175
rect 163777 209147 163811 209175
rect 163839 209147 163887 209175
rect 163577 209113 163887 209147
rect 163577 209085 163625 209113
rect 163653 209085 163687 209113
rect 163715 209085 163749 209113
rect 163777 209085 163811 209113
rect 163839 209085 163887 209113
rect 163577 209051 163887 209085
rect 163577 209023 163625 209051
rect 163653 209023 163687 209051
rect 163715 209023 163749 209051
rect 163777 209023 163811 209051
rect 163839 209023 163887 209051
rect 163577 208989 163887 209023
rect 163577 208961 163625 208989
rect 163653 208961 163687 208989
rect 163715 208961 163749 208989
rect 163777 208961 163811 208989
rect 163839 208961 163887 208989
rect 163577 200175 163887 208961
rect 163577 200147 163625 200175
rect 163653 200147 163687 200175
rect 163715 200147 163749 200175
rect 163777 200147 163811 200175
rect 163839 200147 163887 200175
rect 163577 200113 163887 200147
rect 163577 200085 163625 200113
rect 163653 200085 163687 200113
rect 163715 200085 163749 200113
rect 163777 200085 163811 200113
rect 163839 200085 163887 200113
rect 163577 200051 163887 200085
rect 163577 200023 163625 200051
rect 163653 200023 163687 200051
rect 163715 200023 163749 200051
rect 163777 200023 163811 200051
rect 163839 200023 163887 200051
rect 163577 199989 163887 200023
rect 163577 199961 163625 199989
rect 163653 199961 163687 199989
rect 163715 199961 163749 199989
rect 163777 199961 163811 199989
rect 163839 199961 163887 199989
rect 163577 191175 163887 199961
rect 163577 191147 163625 191175
rect 163653 191147 163687 191175
rect 163715 191147 163749 191175
rect 163777 191147 163811 191175
rect 163839 191147 163887 191175
rect 163577 191113 163887 191147
rect 163577 191085 163625 191113
rect 163653 191085 163687 191113
rect 163715 191085 163749 191113
rect 163777 191085 163811 191113
rect 163839 191085 163887 191113
rect 163577 191051 163887 191085
rect 163577 191023 163625 191051
rect 163653 191023 163687 191051
rect 163715 191023 163749 191051
rect 163777 191023 163811 191051
rect 163839 191023 163887 191051
rect 163577 190989 163887 191023
rect 163577 190961 163625 190989
rect 163653 190961 163687 190989
rect 163715 190961 163749 190989
rect 163777 190961 163811 190989
rect 163839 190961 163887 190989
rect 163577 182175 163887 190961
rect 163577 182147 163625 182175
rect 163653 182147 163687 182175
rect 163715 182147 163749 182175
rect 163777 182147 163811 182175
rect 163839 182147 163887 182175
rect 163577 182113 163887 182147
rect 163577 182085 163625 182113
rect 163653 182085 163687 182113
rect 163715 182085 163749 182113
rect 163777 182085 163811 182113
rect 163839 182085 163887 182113
rect 163577 182051 163887 182085
rect 163577 182023 163625 182051
rect 163653 182023 163687 182051
rect 163715 182023 163749 182051
rect 163777 182023 163811 182051
rect 163839 182023 163887 182051
rect 163577 181989 163887 182023
rect 163577 181961 163625 181989
rect 163653 181961 163687 181989
rect 163715 181961 163749 181989
rect 163777 181961 163811 181989
rect 163839 181961 163887 181989
rect 163577 173175 163887 181961
rect 163577 173147 163625 173175
rect 163653 173147 163687 173175
rect 163715 173147 163749 173175
rect 163777 173147 163811 173175
rect 163839 173147 163887 173175
rect 163577 173113 163887 173147
rect 163577 173085 163625 173113
rect 163653 173085 163687 173113
rect 163715 173085 163749 173113
rect 163777 173085 163811 173113
rect 163839 173085 163887 173113
rect 163577 173051 163887 173085
rect 163577 173023 163625 173051
rect 163653 173023 163687 173051
rect 163715 173023 163749 173051
rect 163777 173023 163811 173051
rect 163839 173023 163887 173051
rect 163577 172989 163887 173023
rect 163577 172961 163625 172989
rect 163653 172961 163687 172989
rect 163715 172961 163749 172989
rect 163777 172961 163811 172989
rect 163839 172961 163887 172989
rect 163577 164175 163887 172961
rect 163577 164147 163625 164175
rect 163653 164147 163687 164175
rect 163715 164147 163749 164175
rect 163777 164147 163811 164175
rect 163839 164147 163887 164175
rect 163577 164113 163887 164147
rect 163577 164085 163625 164113
rect 163653 164085 163687 164113
rect 163715 164085 163749 164113
rect 163777 164085 163811 164113
rect 163839 164085 163887 164113
rect 163577 164051 163887 164085
rect 163577 164023 163625 164051
rect 163653 164023 163687 164051
rect 163715 164023 163749 164051
rect 163777 164023 163811 164051
rect 163839 164023 163887 164051
rect 163577 163989 163887 164023
rect 163577 163961 163625 163989
rect 163653 163961 163687 163989
rect 163715 163961 163749 163989
rect 163777 163961 163811 163989
rect 163839 163961 163887 163989
rect 163577 155175 163887 163961
rect 163577 155147 163625 155175
rect 163653 155147 163687 155175
rect 163715 155147 163749 155175
rect 163777 155147 163811 155175
rect 163839 155147 163887 155175
rect 163577 155113 163887 155147
rect 163577 155085 163625 155113
rect 163653 155085 163687 155113
rect 163715 155085 163749 155113
rect 163777 155085 163811 155113
rect 163839 155085 163887 155113
rect 163577 155051 163887 155085
rect 163577 155023 163625 155051
rect 163653 155023 163687 155051
rect 163715 155023 163749 155051
rect 163777 155023 163811 155051
rect 163839 155023 163887 155051
rect 163577 154989 163887 155023
rect 163577 154961 163625 154989
rect 163653 154961 163687 154989
rect 163715 154961 163749 154989
rect 163777 154961 163811 154989
rect 163839 154961 163887 154989
rect 163577 146175 163887 154961
rect 163577 146147 163625 146175
rect 163653 146147 163687 146175
rect 163715 146147 163749 146175
rect 163777 146147 163811 146175
rect 163839 146147 163887 146175
rect 163577 146113 163887 146147
rect 163577 146085 163625 146113
rect 163653 146085 163687 146113
rect 163715 146085 163749 146113
rect 163777 146085 163811 146113
rect 163839 146085 163887 146113
rect 163577 146051 163887 146085
rect 163577 146023 163625 146051
rect 163653 146023 163687 146051
rect 163715 146023 163749 146051
rect 163777 146023 163811 146051
rect 163839 146023 163887 146051
rect 163577 145989 163887 146023
rect 163577 145961 163625 145989
rect 163653 145961 163687 145989
rect 163715 145961 163749 145989
rect 163777 145961 163811 145989
rect 163839 145961 163887 145989
rect 163577 137175 163887 145961
rect 163577 137147 163625 137175
rect 163653 137147 163687 137175
rect 163715 137147 163749 137175
rect 163777 137147 163811 137175
rect 163839 137147 163887 137175
rect 163577 137113 163887 137147
rect 163577 137085 163625 137113
rect 163653 137085 163687 137113
rect 163715 137085 163749 137113
rect 163777 137085 163811 137113
rect 163839 137085 163887 137113
rect 163577 137051 163887 137085
rect 163577 137023 163625 137051
rect 163653 137023 163687 137051
rect 163715 137023 163749 137051
rect 163777 137023 163811 137051
rect 163839 137023 163887 137051
rect 163577 136989 163887 137023
rect 163577 136961 163625 136989
rect 163653 136961 163687 136989
rect 163715 136961 163749 136989
rect 163777 136961 163811 136989
rect 163839 136961 163887 136989
rect 163577 128175 163887 136961
rect 163577 128147 163625 128175
rect 163653 128147 163687 128175
rect 163715 128147 163749 128175
rect 163777 128147 163811 128175
rect 163839 128147 163887 128175
rect 163577 128113 163887 128147
rect 163577 128085 163625 128113
rect 163653 128085 163687 128113
rect 163715 128085 163749 128113
rect 163777 128085 163811 128113
rect 163839 128085 163887 128113
rect 163577 128051 163887 128085
rect 163577 128023 163625 128051
rect 163653 128023 163687 128051
rect 163715 128023 163749 128051
rect 163777 128023 163811 128051
rect 163839 128023 163887 128051
rect 163577 127989 163887 128023
rect 163577 127961 163625 127989
rect 163653 127961 163687 127989
rect 163715 127961 163749 127989
rect 163777 127961 163811 127989
rect 163839 127961 163887 127989
rect 163577 119175 163887 127961
rect 163577 119147 163625 119175
rect 163653 119147 163687 119175
rect 163715 119147 163749 119175
rect 163777 119147 163811 119175
rect 163839 119147 163887 119175
rect 163577 119113 163887 119147
rect 163577 119085 163625 119113
rect 163653 119085 163687 119113
rect 163715 119085 163749 119113
rect 163777 119085 163811 119113
rect 163839 119085 163887 119113
rect 163577 119051 163887 119085
rect 163577 119023 163625 119051
rect 163653 119023 163687 119051
rect 163715 119023 163749 119051
rect 163777 119023 163811 119051
rect 163839 119023 163887 119051
rect 163577 118989 163887 119023
rect 163577 118961 163625 118989
rect 163653 118961 163687 118989
rect 163715 118961 163749 118989
rect 163777 118961 163811 118989
rect 163839 118961 163887 118989
rect 163577 110175 163887 118961
rect 163577 110147 163625 110175
rect 163653 110147 163687 110175
rect 163715 110147 163749 110175
rect 163777 110147 163811 110175
rect 163839 110147 163887 110175
rect 163577 110113 163887 110147
rect 163577 110085 163625 110113
rect 163653 110085 163687 110113
rect 163715 110085 163749 110113
rect 163777 110085 163811 110113
rect 163839 110085 163887 110113
rect 163577 110051 163887 110085
rect 163577 110023 163625 110051
rect 163653 110023 163687 110051
rect 163715 110023 163749 110051
rect 163777 110023 163811 110051
rect 163839 110023 163887 110051
rect 163577 109989 163887 110023
rect 163577 109961 163625 109989
rect 163653 109961 163687 109989
rect 163715 109961 163749 109989
rect 163777 109961 163811 109989
rect 163839 109961 163887 109989
rect 163577 101175 163887 109961
rect 163577 101147 163625 101175
rect 163653 101147 163687 101175
rect 163715 101147 163749 101175
rect 163777 101147 163811 101175
rect 163839 101147 163887 101175
rect 163577 101113 163887 101147
rect 163577 101085 163625 101113
rect 163653 101085 163687 101113
rect 163715 101085 163749 101113
rect 163777 101085 163811 101113
rect 163839 101085 163887 101113
rect 163577 101051 163887 101085
rect 163577 101023 163625 101051
rect 163653 101023 163687 101051
rect 163715 101023 163749 101051
rect 163777 101023 163811 101051
rect 163839 101023 163887 101051
rect 163577 100989 163887 101023
rect 163577 100961 163625 100989
rect 163653 100961 163687 100989
rect 163715 100961 163749 100989
rect 163777 100961 163811 100989
rect 163839 100961 163887 100989
rect 163577 92175 163887 100961
rect 163577 92147 163625 92175
rect 163653 92147 163687 92175
rect 163715 92147 163749 92175
rect 163777 92147 163811 92175
rect 163839 92147 163887 92175
rect 163577 92113 163887 92147
rect 163577 92085 163625 92113
rect 163653 92085 163687 92113
rect 163715 92085 163749 92113
rect 163777 92085 163811 92113
rect 163839 92085 163887 92113
rect 163577 92051 163887 92085
rect 163577 92023 163625 92051
rect 163653 92023 163687 92051
rect 163715 92023 163749 92051
rect 163777 92023 163811 92051
rect 163839 92023 163887 92051
rect 163577 91989 163887 92023
rect 163577 91961 163625 91989
rect 163653 91961 163687 91989
rect 163715 91961 163749 91989
rect 163777 91961 163811 91989
rect 163839 91961 163887 91989
rect 163577 83175 163887 91961
rect 163577 83147 163625 83175
rect 163653 83147 163687 83175
rect 163715 83147 163749 83175
rect 163777 83147 163811 83175
rect 163839 83147 163887 83175
rect 163577 83113 163887 83147
rect 163577 83085 163625 83113
rect 163653 83085 163687 83113
rect 163715 83085 163749 83113
rect 163777 83085 163811 83113
rect 163839 83085 163887 83113
rect 163577 83051 163887 83085
rect 163577 83023 163625 83051
rect 163653 83023 163687 83051
rect 163715 83023 163749 83051
rect 163777 83023 163811 83051
rect 163839 83023 163887 83051
rect 163577 82989 163887 83023
rect 163577 82961 163625 82989
rect 163653 82961 163687 82989
rect 163715 82961 163749 82989
rect 163777 82961 163811 82989
rect 163839 82961 163887 82989
rect 163577 74175 163887 82961
rect 163577 74147 163625 74175
rect 163653 74147 163687 74175
rect 163715 74147 163749 74175
rect 163777 74147 163811 74175
rect 163839 74147 163887 74175
rect 163577 74113 163887 74147
rect 163577 74085 163625 74113
rect 163653 74085 163687 74113
rect 163715 74085 163749 74113
rect 163777 74085 163811 74113
rect 163839 74085 163887 74113
rect 163577 74051 163887 74085
rect 163577 74023 163625 74051
rect 163653 74023 163687 74051
rect 163715 74023 163749 74051
rect 163777 74023 163811 74051
rect 163839 74023 163887 74051
rect 163577 73989 163887 74023
rect 163577 73961 163625 73989
rect 163653 73961 163687 73989
rect 163715 73961 163749 73989
rect 163777 73961 163811 73989
rect 163839 73961 163887 73989
rect 163577 65175 163887 73961
rect 163577 65147 163625 65175
rect 163653 65147 163687 65175
rect 163715 65147 163749 65175
rect 163777 65147 163811 65175
rect 163839 65147 163887 65175
rect 163577 65113 163887 65147
rect 163577 65085 163625 65113
rect 163653 65085 163687 65113
rect 163715 65085 163749 65113
rect 163777 65085 163811 65113
rect 163839 65085 163887 65113
rect 163577 65051 163887 65085
rect 163577 65023 163625 65051
rect 163653 65023 163687 65051
rect 163715 65023 163749 65051
rect 163777 65023 163811 65051
rect 163839 65023 163887 65051
rect 163577 64989 163887 65023
rect 163577 64961 163625 64989
rect 163653 64961 163687 64989
rect 163715 64961 163749 64989
rect 163777 64961 163811 64989
rect 163839 64961 163887 64989
rect 163577 56175 163887 64961
rect 163577 56147 163625 56175
rect 163653 56147 163687 56175
rect 163715 56147 163749 56175
rect 163777 56147 163811 56175
rect 163839 56147 163887 56175
rect 163577 56113 163887 56147
rect 163577 56085 163625 56113
rect 163653 56085 163687 56113
rect 163715 56085 163749 56113
rect 163777 56085 163811 56113
rect 163839 56085 163887 56113
rect 163577 56051 163887 56085
rect 163577 56023 163625 56051
rect 163653 56023 163687 56051
rect 163715 56023 163749 56051
rect 163777 56023 163811 56051
rect 163839 56023 163887 56051
rect 163577 55989 163887 56023
rect 163577 55961 163625 55989
rect 163653 55961 163687 55989
rect 163715 55961 163749 55989
rect 163777 55961 163811 55989
rect 163839 55961 163887 55989
rect 163577 47175 163887 55961
rect 163577 47147 163625 47175
rect 163653 47147 163687 47175
rect 163715 47147 163749 47175
rect 163777 47147 163811 47175
rect 163839 47147 163887 47175
rect 163577 47113 163887 47147
rect 163577 47085 163625 47113
rect 163653 47085 163687 47113
rect 163715 47085 163749 47113
rect 163777 47085 163811 47113
rect 163839 47085 163887 47113
rect 163577 47051 163887 47085
rect 163577 47023 163625 47051
rect 163653 47023 163687 47051
rect 163715 47023 163749 47051
rect 163777 47023 163811 47051
rect 163839 47023 163887 47051
rect 163577 46989 163887 47023
rect 163577 46961 163625 46989
rect 163653 46961 163687 46989
rect 163715 46961 163749 46989
rect 163777 46961 163811 46989
rect 163839 46961 163887 46989
rect 163577 38175 163887 46961
rect 163577 38147 163625 38175
rect 163653 38147 163687 38175
rect 163715 38147 163749 38175
rect 163777 38147 163811 38175
rect 163839 38147 163887 38175
rect 163577 38113 163887 38147
rect 163577 38085 163625 38113
rect 163653 38085 163687 38113
rect 163715 38085 163749 38113
rect 163777 38085 163811 38113
rect 163839 38085 163887 38113
rect 163577 38051 163887 38085
rect 163577 38023 163625 38051
rect 163653 38023 163687 38051
rect 163715 38023 163749 38051
rect 163777 38023 163811 38051
rect 163839 38023 163887 38051
rect 163577 37989 163887 38023
rect 163577 37961 163625 37989
rect 163653 37961 163687 37989
rect 163715 37961 163749 37989
rect 163777 37961 163811 37989
rect 163839 37961 163887 37989
rect 163577 29175 163887 37961
rect 163577 29147 163625 29175
rect 163653 29147 163687 29175
rect 163715 29147 163749 29175
rect 163777 29147 163811 29175
rect 163839 29147 163887 29175
rect 163577 29113 163887 29147
rect 163577 29085 163625 29113
rect 163653 29085 163687 29113
rect 163715 29085 163749 29113
rect 163777 29085 163811 29113
rect 163839 29085 163887 29113
rect 163577 29051 163887 29085
rect 163577 29023 163625 29051
rect 163653 29023 163687 29051
rect 163715 29023 163749 29051
rect 163777 29023 163811 29051
rect 163839 29023 163887 29051
rect 163577 28989 163887 29023
rect 163577 28961 163625 28989
rect 163653 28961 163687 28989
rect 163715 28961 163749 28989
rect 163777 28961 163811 28989
rect 163839 28961 163887 28989
rect 163577 20175 163887 28961
rect 163577 20147 163625 20175
rect 163653 20147 163687 20175
rect 163715 20147 163749 20175
rect 163777 20147 163811 20175
rect 163839 20147 163887 20175
rect 163577 20113 163887 20147
rect 163577 20085 163625 20113
rect 163653 20085 163687 20113
rect 163715 20085 163749 20113
rect 163777 20085 163811 20113
rect 163839 20085 163887 20113
rect 163577 20051 163887 20085
rect 163577 20023 163625 20051
rect 163653 20023 163687 20051
rect 163715 20023 163749 20051
rect 163777 20023 163811 20051
rect 163839 20023 163887 20051
rect 163577 19989 163887 20023
rect 163577 19961 163625 19989
rect 163653 19961 163687 19989
rect 163715 19961 163749 19989
rect 163777 19961 163811 19989
rect 163839 19961 163887 19989
rect 163577 11175 163887 19961
rect 163577 11147 163625 11175
rect 163653 11147 163687 11175
rect 163715 11147 163749 11175
rect 163777 11147 163811 11175
rect 163839 11147 163887 11175
rect 163577 11113 163887 11147
rect 163577 11085 163625 11113
rect 163653 11085 163687 11113
rect 163715 11085 163749 11113
rect 163777 11085 163811 11113
rect 163839 11085 163887 11113
rect 163577 11051 163887 11085
rect 163577 11023 163625 11051
rect 163653 11023 163687 11051
rect 163715 11023 163749 11051
rect 163777 11023 163811 11051
rect 163839 11023 163887 11051
rect 163577 10989 163887 11023
rect 163577 10961 163625 10989
rect 163653 10961 163687 10989
rect 163715 10961 163749 10989
rect 163777 10961 163811 10989
rect 163839 10961 163887 10989
rect 163577 2175 163887 10961
rect 163577 2147 163625 2175
rect 163653 2147 163687 2175
rect 163715 2147 163749 2175
rect 163777 2147 163811 2175
rect 163839 2147 163887 2175
rect 163577 2113 163887 2147
rect 163577 2085 163625 2113
rect 163653 2085 163687 2113
rect 163715 2085 163749 2113
rect 163777 2085 163811 2113
rect 163839 2085 163887 2113
rect 163577 2051 163887 2085
rect 163577 2023 163625 2051
rect 163653 2023 163687 2051
rect 163715 2023 163749 2051
rect 163777 2023 163811 2051
rect 163839 2023 163887 2051
rect 163577 1989 163887 2023
rect 163577 1961 163625 1989
rect 163653 1961 163687 1989
rect 163715 1961 163749 1989
rect 163777 1961 163811 1989
rect 163839 1961 163887 1989
rect 163577 -80 163887 1961
rect 163577 -108 163625 -80
rect 163653 -108 163687 -80
rect 163715 -108 163749 -80
rect 163777 -108 163811 -80
rect 163839 -108 163887 -80
rect 163577 -142 163887 -108
rect 163577 -170 163625 -142
rect 163653 -170 163687 -142
rect 163715 -170 163749 -142
rect 163777 -170 163811 -142
rect 163839 -170 163887 -142
rect 163577 -204 163887 -170
rect 163577 -232 163625 -204
rect 163653 -232 163687 -204
rect 163715 -232 163749 -204
rect 163777 -232 163811 -204
rect 163839 -232 163887 -204
rect 163577 -266 163887 -232
rect 163577 -294 163625 -266
rect 163653 -294 163687 -266
rect 163715 -294 163749 -266
rect 163777 -294 163811 -266
rect 163839 -294 163887 -266
rect 163577 -822 163887 -294
rect 165437 299086 165747 299134
rect 165437 299058 165485 299086
rect 165513 299058 165547 299086
rect 165575 299058 165609 299086
rect 165637 299058 165671 299086
rect 165699 299058 165747 299086
rect 165437 299024 165747 299058
rect 165437 298996 165485 299024
rect 165513 298996 165547 299024
rect 165575 298996 165609 299024
rect 165637 298996 165671 299024
rect 165699 298996 165747 299024
rect 165437 298962 165747 298996
rect 165437 298934 165485 298962
rect 165513 298934 165547 298962
rect 165575 298934 165609 298962
rect 165637 298934 165671 298962
rect 165699 298934 165747 298962
rect 165437 298900 165747 298934
rect 165437 298872 165485 298900
rect 165513 298872 165547 298900
rect 165575 298872 165609 298900
rect 165637 298872 165671 298900
rect 165699 298872 165747 298900
rect 165437 293175 165747 298872
rect 165437 293147 165485 293175
rect 165513 293147 165547 293175
rect 165575 293147 165609 293175
rect 165637 293147 165671 293175
rect 165699 293147 165747 293175
rect 165437 293113 165747 293147
rect 165437 293085 165485 293113
rect 165513 293085 165547 293113
rect 165575 293085 165609 293113
rect 165637 293085 165671 293113
rect 165699 293085 165747 293113
rect 165437 293051 165747 293085
rect 165437 293023 165485 293051
rect 165513 293023 165547 293051
rect 165575 293023 165609 293051
rect 165637 293023 165671 293051
rect 165699 293023 165747 293051
rect 165437 292989 165747 293023
rect 165437 292961 165485 292989
rect 165513 292961 165547 292989
rect 165575 292961 165609 292989
rect 165637 292961 165671 292989
rect 165699 292961 165747 292989
rect 165437 284175 165747 292961
rect 165437 284147 165485 284175
rect 165513 284147 165547 284175
rect 165575 284147 165609 284175
rect 165637 284147 165671 284175
rect 165699 284147 165747 284175
rect 165437 284113 165747 284147
rect 165437 284085 165485 284113
rect 165513 284085 165547 284113
rect 165575 284085 165609 284113
rect 165637 284085 165671 284113
rect 165699 284085 165747 284113
rect 165437 284051 165747 284085
rect 165437 284023 165485 284051
rect 165513 284023 165547 284051
rect 165575 284023 165609 284051
rect 165637 284023 165671 284051
rect 165699 284023 165747 284051
rect 165437 283989 165747 284023
rect 165437 283961 165485 283989
rect 165513 283961 165547 283989
rect 165575 283961 165609 283989
rect 165637 283961 165671 283989
rect 165699 283961 165747 283989
rect 165437 275175 165747 283961
rect 165437 275147 165485 275175
rect 165513 275147 165547 275175
rect 165575 275147 165609 275175
rect 165637 275147 165671 275175
rect 165699 275147 165747 275175
rect 165437 275113 165747 275147
rect 165437 275085 165485 275113
rect 165513 275085 165547 275113
rect 165575 275085 165609 275113
rect 165637 275085 165671 275113
rect 165699 275085 165747 275113
rect 165437 275051 165747 275085
rect 165437 275023 165485 275051
rect 165513 275023 165547 275051
rect 165575 275023 165609 275051
rect 165637 275023 165671 275051
rect 165699 275023 165747 275051
rect 165437 274989 165747 275023
rect 165437 274961 165485 274989
rect 165513 274961 165547 274989
rect 165575 274961 165609 274989
rect 165637 274961 165671 274989
rect 165699 274961 165747 274989
rect 165437 266175 165747 274961
rect 165437 266147 165485 266175
rect 165513 266147 165547 266175
rect 165575 266147 165609 266175
rect 165637 266147 165671 266175
rect 165699 266147 165747 266175
rect 165437 266113 165747 266147
rect 165437 266085 165485 266113
rect 165513 266085 165547 266113
rect 165575 266085 165609 266113
rect 165637 266085 165671 266113
rect 165699 266085 165747 266113
rect 165437 266051 165747 266085
rect 165437 266023 165485 266051
rect 165513 266023 165547 266051
rect 165575 266023 165609 266051
rect 165637 266023 165671 266051
rect 165699 266023 165747 266051
rect 165437 265989 165747 266023
rect 165437 265961 165485 265989
rect 165513 265961 165547 265989
rect 165575 265961 165609 265989
rect 165637 265961 165671 265989
rect 165699 265961 165747 265989
rect 165437 257175 165747 265961
rect 165437 257147 165485 257175
rect 165513 257147 165547 257175
rect 165575 257147 165609 257175
rect 165637 257147 165671 257175
rect 165699 257147 165747 257175
rect 165437 257113 165747 257147
rect 165437 257085 165485 257113
rect 165513 257085 165547 257113
rect 165575 257085 165609 257113
rect 165637 257085 165671 257113
rect 165699 257085 165747 257113
rect 165437 257051 165747 257085
rect 165437 257023 165485 257051
rect 165513 257023 165547 257051
rect 165575 257023 165609 257051
rect 165637 257023 165671 257051
rect 165699 257023 165747 257051
rect 165437 256989 165747 257023
rect 165437 256961 165485 256989
rect 165513 256961 165547 256989
rect 165575 256961 165609 256989
rect 165637 256961 165671 256989
rect 165699 256961 165747 256989
rect 165437 248175 165747 256961
rect 165437 248147 165485 248175
rect 165513 248147 165547 248175
rect 165575 248147 165609 248175
rect 165637 248147 165671 248175
rect 165699 248147 165747 248175
rect 165437 248113 165747 248147
rect 165437 248085 165485 248113
rect 165513 248085 165547 248113
rect 165575 248085 165609 248113
rect 165637 248085 165671 248113
rect 165699 248085 165747 248113
rect 165437 248051 165747 248085
rect 165437 248023 165485 248051
rect 165513 248023 165547 248051
rect 165575 248023 165609 248051
rect 165637 248023 165671 248051
rect 165699 248023 165747 248051
rect 165437 247989 165747 248023
rect 165437 247961 165485 247989
rect 165513 247961 165547 247989
rect 165575 247961 165609 247989
rect 165637 247961 165671 247989
rect 165699 247961 165747 247989
rect 165437 239175 165747 247961
rect 165437 239147 165485 239175
rect 165513 239147 165547 239175
rect 165575 239147 165609 239175
rect 165637 239147 165671 239175
rect 165699 239147 165747 239175
rect 165437 239113 165747 239147
rect 165437 239085 165485 239113
rect 165513 239085 165547 239113
rect 165575 239085 165609 239113
rect 165637 239085 165671 239113
rect 165699 239085 165747 239113
rect 165437 239051 165747 239085
rect 165437 239023 165485 239051
rect 165513 239023 165547 239051
rect 165575 239023 165609 239051
rect 165637 239023 165671 239051
rect 165699 239023 165747 239051
rect 165437 238989 165747 239023
rect 165437 238961 165485 238989
rect 165513 238961 165547 238989
rect 165575 238961 165609 238989
rect 165637 238961 165671 238989
rect 165699 238961 165747 238989
rect 165437 230175 165747 238961
rect 165437 230147 165485 230175
rect 165513 230147 165547 230175
rect 165575 230147 165609 230175
rect 165637 230147 165671 230175
rect 165699 230147 165747 230175
rect 165437 230113 165747 230147
rect 165437 230085 165485 230113
rect 165513 230085 165547 230113
rect 165575 230085 165609 230113
rect 165637 230085 165671 230113
rect 165699 230085 165747 230113
rect 165437 230051 165747 230085
rect 165437 230023 165485 230051
rect 165513 230023 165547 230051
rect 165575 230023 165609 230051
rect 165637 230023 165671 230051
rect 165699 230023 165747 230051
rect 165437 229989 165747 230023
rect 165437 229961 165485 229989
rect 165513 229961 165547 229989
rect 165575 229961 165609 229989
rect 165637 229961 165671 229989
rect 165699 229961 165747 229989
rect 165437 221175 165747 229961
rect 165437 221147 165485 221175
rect 165513 221147 165547 221175
rect 165575 221147 165609 221175
rect 165637 221147 165671 221175
rect 165699 221147 165747 221175
rect 165437 221113 165747 221147
rect 165437 221085 165485 221113
rect 165513 221085 165547 221113
rect 165575 221085 165609 221113
rect 165637 221085 165671 221113
rect 165699 221085 165747 221113
rect 165437 221051 165747 221085
rect 165437 221023 165485 221051
rect 165513 221023 165547 221051
rect 165575 221023 165609 221051
rect 165637 221023 165671 221051
rect 165699 221023 165747 221051
rect 165437 220989 165747 221023
rect 165437 220961 165485 220989
rect 165513 220961 165547 220989
rect 165575 220961 165609 220989
rect 165637 220961 165671 220989
rect 165699 220961 165747 220989
rect 165437 212175 165747 220961
rect 165437 212147 165485 212175
rect 165513 212147 165547 212175
rect 165575 212147 165609 212175
rect 165637 212147 165671 212175
rect 165699 212147 165747 212175
rect 165437 212113 165747 212147
rect 165437 212085 165485 212113
rect 165513 212085 165547 212113
rect 165575 212085 165609 212113
rect 165637 212085 165671 212113
rect 165699 212085 165747 212113
rect 165437 212051 165747 212085
rect 165437 212023 165485 212051
rect 165513 212023 165547 212051
rect 165575 212023 165609 212051
rect 165637 212023 165671 212051
rect 165699 212023 165747 212051
rect 165437 211989 165747 212023
rect 165437 211961 165485 211989
rect 165513 211961 165547 211989
rect 165575 211961 165609 211989
rect 165637 211961 165671 211989
rect 165699 211961 165747 211989
rect 165437 203175 165747 211961
rect 165437 203147 165485 203175
rect 165513 203147 165547 203175
rect 165575 203147 165609 203175
rect 165637 203147 165671 203175
rect 165699 203147 165747 203175
rect 165437 203113 165747 203147
rect 165437 203085 165485 203113
rect 165513 203085 165547 203113
rect 165575 203085 165609 203113
rect 165637 203085 165671 203113
rect 165699 203085 165747 203113
rect 165437 203051 165747 203085
rect 165437 203023 165485 203051
rect 165513 203023 165547 203051
rect 165575 203023 165609 203051
rect 165637 203023 165671 203051
rect 165699 203023 165747 203051
rect 165437 202989 165747 203023
rect 165437 202961 165485 202989
rect 165513 202961 165547 202989
rect 165575 202961 165609 202989
rect 165637 202961 165671 202989
rect 165699 202961 165747 202989
rect 165437 194175 165747 202961
rect 165437 194147 165485 194175
rect 165513 194147 165547 194175
rect 165575 194147 165609 194175
rect 165637 194147 165671 194175
rect 165699 194147 165747 194175
rect 165437 194113 165747 194147
rect 165437 194085 165485 194113
rect 165513 194085 165547 194113
rect 165575 194085 165609 194113
rect 165637 194085 165671 194113
rect 165699 194085 165747 194113
rect 165437 194051 165747 194085
rect 165437 194023 165485 194051
rect 165513 194023 165547 194051
rect 165575 194023 165609 194051
rect 165637 194023 165671 194051
rect 165699 194023 165747 194051
rect 165437 193989 165747 194023
rect 165437 193961 165485 193989
rect 165513 193961 165547 193989
rect 165575 193961 165609 193989
rect 165637 193961 165671 193989
rect 165699 193961 165747 193989
rect 165437 185175 165747 193961
rect 165437 185147 165485 185175
rect 165513 185147 165547 185175
rect 165575 185147 165609 185175
rect 165637 185147 165671 185175
rect 165699 185147 165747 185175
rect 165437 185113 165747 185147
rect 165437 185085 165485 185113
rect 165513 185085 165547 185113
rect 165575 185085 165609 185113
rect 165637 185085 165671 185113
rect 165699 185085 165747 185113
rect 165437 185051 165747 185085
rect 165437 185023 165485 185051
rect 165513 185023 165547 185051
rect 165575 185023 165609 185051
rect 165637 185023 165671 185051
rect 165699 185023 165747 185051
rect 165437 184989 165747 185023
rect 165437 184961 165485 184989
rect 165513 184961 165547 184989
rect 165575 184961 165609 184989
rect 165637 184961 165671 184989
rect 165699 184961 165747 184989
rect 165437 176175 165747 184961
rect 165437 176147 165485 176175
rect 165513 176147 165547 176175
rect 165575 176147 165609 176175
rect 165637 176147 165671 176175
rect 165699 176147 165747 176175
rect 165437 176113 165747 176147
rect 165437 176085 165485 176113
rect 165513 176085 165547 176113
rect 165575 176085 165609 176113
rect 165637 176085 165671 176113
rect 165699 176085 165747 176113
rect 165437 176051 165747 176085
rect 165437 176023 165485 176051
rect 165513 176023 165547 176051
rect 165575 176023 165609 176051
rect 165637 176023 165671 176051
rect 165699 176023 165747 176051
rect 165437 175989 165747 176023
rect 165437 175961 165485 175989
rect 165513 175961 165547 175989
rect 165575 175961 165609 175989
rect 165637 175961 165671 175989
rect 165699 175961 165747 175989
rect 165437 167175 165747 175961
rect 165437 167147 165485 167175
rect 165513 167147 165547 167175
rect 165575 167147 165609 167175
rect 165637 167147 165671 167175
rect 165699 167147 165747 167175
rect 165437 167113 165747 167147
rect 165437 167085 165485 167113
rect 165513 167085 165547 167113
rect 165575 167085 165609 167113
rect 165637 167085 165671 167113
rect 165699 167085 165747 167113
rect 165437 167051 165747 167085
rect 165437 167023 165485 167051
rect 165513 167023 165547 167051
rect 165575 167023 165609 167051
rect 165637 167023 165671 167051
rect 165699 167023 165747 167051
rect 165437 166989 165747 167023
rect 165437 166961 165485 166989
rect 165513 166961 165547 166989
rect 165575 166961 165609 166989
rect 165637 166961 165671 166989
rect 165699 166961 165747 166989
rect 165437 158175 165747 166961
rect 165437 158147 165485 158175
rect 165513 158147 165547 158175
rect 165575 158147 165609 158175
rect 165637 158147 165671 158175
rect 165699 158147 165747 158175
rect 165437 158113 165747 158147
rect 165437 158085 165485 158113
rect 165513 158085 165547 158113
rect 165575 158085 165609 158113
rect 165637 158085 165671 158113
rect 165699 158085 165747 158113
rect 165437 158051 165747 158085
rect 165437 158023 165485 158051
rect 165513 158023 165547 158051
rect 165575 158023 165609 158051
rect 165637 158023 165671 158051
rect 165699 158023 165747 158051
rect 165437 157989 165747 158023
rect 165437 157961 165485 157989
rect 165513 157961 165547 157989
rect 165575 157961 165609 157989
rect 165637 157961 165671 157989
rect 165699 157961 165747 157989
rect 165437 149175 165747 157961
rect 165437 149147 165485 149175
rect 165513 149147 165547 149175
rect 165575 149147 165609 149175
rect 165637 149147 165671 149175
rect 165699 149147 165747 149175
rect 165437 149113 165747 149147
rect 165437 149085 165485 149113
rect 165513 149085 165547 149113
rect 165575 149085 165609 149113
rect 165637 149085 165671 149113
rect 165699 149085 165747 149113
rect 165437 149051 165747 149085
rect 165437 149023 165485 149051
rect 165513 149023 165547 149051
rect 165575 149023 165609 149051
rect 165637 149023 165671 149051
rect 165699 149023 165747 149051
rect 165437 148989 165747 149023
rect 165437 148961 165485 148989
rect 165513 148961 165547 148989
rect 165575 148961 165609 148989
rect 165637 148961 165671 148989
rect 165699 148961 165747 148989
rect 165437 140175 165747 148961
rect 165437 140147 165485 140175
rect 165513 140147 165547 140175
rect 165575 140147 165609 140175
rect 165637 140147 165671 140175
rect 165699 140147 165747 140175
rect 165437 140113 165747 140147
rect 165437 140085 165485 140113
rect 165513 140085 165547 140113
rect 165575 140085 165609 140113
rect 165637 140085 165671 140113
rect 165699 140085 165747 140113
rect 165437 140051 165747 140085
rect 165437 140023 165485 140051
rect 165513 140023 165547 140051
rect 165575 140023 165609 140051
rect 165637 140023 165671 140051
rect 165699 140023 165747 140051
rect 165437 139989 165747 140023
rect 165437 139961 165485 139989
rect 165513 139961 165547 139989
rect 165575 139961 165609 139989
rect 165637 139961 165671 139989
rect 165699 139961 165747 139989
rect 165437 131175 165747 139961
rect 165437 131147 165485 131175
rect 165513 131147 165547 131175
rect 165575 131147 165609 131175
rect 165637 131147 165671 131175
rect 165699 131147 165747 131175
rect 165437 131113 165747 131147
rect 165437 131085 165485 131113
rect 165513 131085 165547 131113
rect 165575 131085 165609 131113
rect 165637 131085 165671 131113
rect 165699 131085 165747 131113
rect 165437 131051 165747 131085
rect 165437 131023 165485 131051
rect 165513 131023 165547 131051
rect 165575 131023 165609 131051
rect 165637 131023 165671 131051
rect 165699 131023 165747 131051
rect 165437 130989 165747 131023
rect 165437 130961 165485 130989
rect 165513 130961 165547 130989
rect 165575 130961 165609 130989
rect 165637 130961 165671 130989
rect 165699 130961 165747 130989
rect 165437 122175 165747 130961
rect 165437 122147 165485 122175
rect 165513 122147 165547 122175
rect 165575 122147 165609 122175
rect 165637 122147 165671 122175
rect 165699 122147 165747 122175
rect 165437 122113 165747 122147
rect 165437 122085 165485 122113
rect 165513 122085 165547 122113
rect 165575 122085 165609 122113
rect 165637 122085 165671 122113
rect 165699 122085 165747 122113
rect 165437 122051 165747 122085
rect 165437 122023 165485 122051
rect 165513 122023 165547 122051
rect 165575 122023 165609 122051
rect 165637 122023 165671 122051
rect 165699 122023 165747 122051
rect 165437 121989 165747 122023
rect 165437 121961 165485 121989
rect 165513 121961 165547 121989
rect 165575 121961 165609 121989
rect 165637 121961 165671 121989
rect 165699 121961 165747 121989
rect 165437 113175 165747 121961
rect 165437 113147 165485 113175
rect 165513 113147 165547 113175
rect 165575 113147 165609 113175
rect 165637 113147 165671 113175
rect 165699 113147 165747 113175
rect 165437 113113 165747 113147
rect 165437 113085 165485 113113
rect 165513 113085 165547 113113
rect 165575 113085 165609 113113
rect 165637 113085 165671 113113
rect 165699 113085 165747 113113
rect 165437 113051 165747 113085
rect 165437 113023 165485 113051
rect 165513 113023 165547 113051
rect 165575 113023 165609 113051
rect 165637 113023 165671 113051
rect 165699 113023 165747 113051
rect 165437 112989 165747 113023
rect 165437 112961 165485 112989
rect 165513 112961 165547 112989
rect 165575 112961 165609 112989
rect 165637 112961 165671 112989
rect 165699 112961 165747 112989
rect 165437 104175 165747 112961
rect 165437 104147 165485 104175
rect 165513 104147 165547 104175
rect 165575 104147 165609 104175
rect 165637 104147 165671 104175
rect 165699 104147 165747 104175
rect 165437 104113 165747 104147
rect 165437 104085 165485 104113
rect 165513 104085 165547 104113
rect 165575 104085 165609 104113
rect 165637 104085 165671 104113
rect 165699 104085 165747 104113
rect 165437 104051 165747 104085
rect 165437 104023 165485 104051
rect 165513 104023 165547 104051
rect 165575 104023 165609 104051
rect 165637 104023 165671 104051
rect 165699 104023 165747 104051
rect 165437 103989 165747 104023
rect 165437 103961 165485 103989
rect 165513 103961 165547 103989
rect 165575 103961 165609 103989
rect 165637 103961 165671 103989
rect 165699 103961 165747 103989
rect 165437 95175 165747 103961
rect 165437 95147 165485 95175
rect 165513 95147 165547 95175
rect 165575 95147 165609 95175
rect 165637 95147 165671 95175
rect 165699 95147 165747 95175
rect 165437 95113 165747 95147
rect 165437 95085 165485 95113
rect 165513 95085 165547 95113
rect 165575 95085 165609 95113
rect 165637 95085 165671 95113
rect 165699 95085 165747 95113
rect 165437 95051 165747 95085
rect 165437 95023 165485 95051
rect 165513 95023 165547 95051
rect 165575 95023 165609 95051
rect 165637 95023 165671 95051
rect 165699 95023 165747 95051
rect 165437 94989 165747 95023
rect 165437 94961 165485 94989
rect 165513 94961 165547 94989
rect 165575 94961 165609 94989
rect 165637 94961 165671 94989
rect 165699 94961 165747 94989
rect 165437 86175 165747 94961
rect 165437 86147 165485 86175
rect 165513 86147 165547 86175
rect 165575 86147 165609 86175
rect 165637 86147 165671 86175
rect 165699 86147 165747 86175
rect 165437 86113 165747 86147
rect 165437 86085 165485 86113
rect 165513 86085 165547 86113
rect 165575 86085 165609 86113
rect 165637 86085 165671 86113
rect 165699 86085 165747 86113
rect 165437 86051 165747 86085
rect 165437 86023 165485 86051
rect 165513 86023 165547 86051
rect 165575 86023 165609 86051
rect 165637 86023 165671 86051
rect 165699 86023 165747 86051
rect 165437 85989 165747 86023
rect 165437 85961 165485 85989
rect 165513 85961 165547 85989
rect 165575 85961 165609 85989
rect 165637 85961 165671 85989
rect 165699 85961 165747 85989
rect 165437 77175 165747 85961
rect 165437 77147 165485 77175
rect 165513 77147 165547 77175
rect 165575 77147 165609 77175
rect 165637 77147 165671 77175
rect 165699 77147 165747 77175
rect 165437 77113 165747 77147
rect 165437 77085 165485 77113
rect 165513 77085 165547 77113
rect 165575 77085 165609 77113
rect 165637 77085 165671 77113
rect 165699 77085 165747 77113
rect 165437 77051 165747 77085
rect 165437 77023 165485 77051
rect 165513 77023 165547 77051
rect 165575 77023 165609 77051
rect 165637 77023 165671 77051
rect 165699 77023 165747 77051
rect 165437 76989 165747 77023
rect 165437 76961 165485 76989
rect 165513 76961 165547 76989
rect 165575 76961 165609 76989
rect 165637 76961 165671 76989
rect 165699 76961 165747 76989
rect 165437 68175 165747 76961
rect 165437 68147 165485 68175
rect 165513 68147 165547 68175
rect 165575 68147 165609 68175
rect 165637 68147 165671 68175
rect 165699 68147 165747 68175
rect 165437 68113 165747 68147
rect 165437 68085 165485 68113
rect 165513 68085 165547 68113
rect 165575 68085 165609 68113
rect 165637 68085 165671 68113
rect 165699 68085 165747 68113
rect 165437 68051 165747 68085
rect 165437 68023 165485 68051
rect 165513 68023 165547 68051
rect 165575 68023 165609 68051
rect 165637 68023 165671 68051
rect 165699 68023 165747 68051
rect 165437 67989 165747 68023
rect 165437 67961 165485 67989
rect 165513 67961 165547 67989
rect 165575 67961 165609 67989
rect 165637 67961 165671 67989
rect 165699 67961 165747 67989
rect 165437 59175 165747 67961
rect 165437 59147 165485 59175
rect 165513 59147 165547 59175
rect 165575 59147 165609 59175
rect 165637 59147 165671 59175
rect 165699 59147 165747 59175
rect 165437 59113 165747 59147
rect 165437 59085 165485 59113
rect 165513 59085 165547 59113
rect 165575 59085 165609 59113
rect 165637 59085 165671 59113
rect 165699 59085 165747 59113
rect 165437 59051 165747 59085
rect 165437 59023 165485 59051
rect 165513 59023 165547 59051
rect 165575 59023 165609 59051
rect 165637 59023 165671 59051
rect 165699 59023 165747 59051
rect 165437 58989 165747 59023
rect 165437 58961 165485 58989
rect 165513 58961 165547 58989
rect 165575 58961 165609 58989
rect 165637 58961 165671 58989
rect 165699 58961 165747 58989
rect 165437 50175 165747 58961
rect 165437 50147 165485 50175
rect 165513 50147 165547 50175
rect 165575 50147 165609 50175
rect 165637 50147 165671 50175
rect 165699 50147 165747 50175
rect 165437 50113 165747 50147
rect 165437 50085 165485 50113
rect 165513 50085 165547 50113
rect 165575 50085 165609 50113
rect 165637 50085 165671 50113
rect 165699 50085 165747 50113
rect 165437 50051 165747 50085
rect 165437 50023 165485 50051
rect 165513 50023 165547 50051
rect 165575 50023 165609 50051
rect 165637 50023 165671 50051
rect 165699 50023 165747 50051
rect 165437 49989 165747 50023
rect 165437 49961 165485 49989
rect 165513 49961 165547 49989
rect 165575 49961 165609 49989
rect 165637 49961 165671 49989
rect 165699 49961 165747 49989
rect 165437 41175 165747 49961
rect 165437 41147 165485 41175
rect 165513 41147 165547 41175
rect 165575 41147 165609 41175
rect 165637 41147 165671 41175
rect 165699 41147 165747 41175
rect 165437 41113 165747 41147
rect 165437 41085 165485 41113
rect 165513 41085 165547 41113
rect 165575 41085 165609 41113
rect 165637 41085 165671 41113
rect 165699 41085 165747 41113
rect 165437 41051 165747 41085
rect 165437 41023 165485 41051
rect 165513 41023 165547 41051
rect 165575 41023 165609 41051
rect 165637 41023 165671 41051
rect 165699 41023 165747 41051
rect 165437 40989 165747 41023
rect 165437 40961 165485 40989
rect 165513 40961 165547 40989
rect 165575 40961 165609 40989
rect 165637 40961 165671 40989
rect 165699 40961 165747 40989
rect 165437 32175 165747 40961
rect 165437 32147 165485 32175
rect 165513 32147 165547 32175
rect 165575 32147 165609 32175
rect 165637 32147 165671 32175
rect 165699 32147 165747 32175
rect 165437 32113 165747 32147
rect 165437 32085 165485 32113
rect 165513 32085 165547 32113
rect 165575 32085 165609 32113
rect 165637 32085 165671 32113
rect 165699 32085 165747 32113
rect 165437 32051 165747 32085
rect 165437 32023 165485 32051
rect 165513 32023 165547 32051
rect 165575 32023 165609 32051
rect 165637 32023 165671 32051
rect 165699 32023 165747 32051
rect 165437 31989 165747 32023
rect 165437 31961 165485 31989
rect 165513 31961 165547 31989
rect 165575 31961 165609 31989
rect 165637 31961 165671 31989
rect 165699 31961 165747 31989
rect 165437 23175 165747 31961
rect 165437 23147 165485 23175
rect 165513 23147 165547 23175
rect 165575 23147 165609 23175
rect 165637 23147 165671 23175
rect 165699 23147 165747 23175
rect 165437 23113 165747 23147
rect 165437 23085 165485 23113
rect 165513 23085 165547 23113
rect 165575 23085 165609 23113
rect 165637 23085 165671 23113
rect 165699 23085 165747 23113
rect 165437 23051 165747 23085
rect 165437 23023 165485 23051
rect 165513 23023 165547 23051
rect 165575 23023 165609 23051
rect 165637 23023 165671 23051
rect 165699 23023 165747 23051
rect 165437 22989 165747 23023
rect 165437 22961 165485 22989
rect 165513 22961 165547 22989
rect 165575 22961 165609 22989
rect 165637 22961 165671 22989
rect 165699 22961 165747 22989
rect 165437 14175 165747 22961
rect 165437 14147 165485 14175
rect 165513 14147 165547 14175
rect 165575 14147 165609 14175
rect 165637 14147 165671 14175
rect 165699 14147 165747 14175
rect 165437 14113 165747 14147
rect 165437 14085 165485 14113
rect 165513 14085 165547 14113
rect 165575 14085 165609 14113
rect 165637 14085 165671 14113
rect 165699 14085 165747 14113
rect 165437 14051 165747 14085
rect 165437 14023 165485 14051
rect 165513 14023 165547 14051
rect 165575 14023 165609 14051
rect 165637 14023 165671 14051
rect 165699 14023 165747 14051
rect 165437 13989 165747 14023
rect 165437 13961 165485 13989
rect 165513 13961 165547 13989
rect 165575 13961 165609 13989
rect 165637 13961 165671 13989
rect 165699 13961 165747 13989
rect 165437 5175 165747 13961
rect 165437 5147 165485 5175
rect 165513 5147 165547 5175
rect 165575 5147 165609 5175
rect 165637 5147 165671 5175
rect 165699 5147 165747 5175
rect 165437 5113 165747 5147
rect 165437 5085 165485 5113
rect 165513 5085 165547 5113
rect 165575 5085 165609 5113
rect 165637 5085 165671 5113
rect 165699 5085 165747 5113
rect 165437 5051 165747 5085
rect 165437 5023 165485 5051
rect 165513 5023 165547 5051
rect 165575 5023 165609 5051
rect 165637 5023 165671 5051
rect 165699 5023 165747 5051
rect 165437 4989 165747 5023
rect 165437 4961 165485 4989
rect 165513 4961 165547 4989
rect 165575 4961 165609 4989
rect 165637 4961 165671 4989
rect 165699 4961 165747 4989
rect 165437 -560 165747 4961
rect 165437 -588 165485 -560
rect 165513 -588 165547 -560
rect 165575 -588 165609 -560
rect 165637 -588 165671 -560
rect 165699 -588 165747 -560
rect 165437 -622 165747 -588
rect 165437 -650 165485 -622
rect 165513 -650 165547 -622
rect 165575 -650 165609 -622
rect 165637 -650 165671 -622
rect 165699 -650 165747 -622
rect 165437 -684 165747 -650
rect 165437 -712 165485 -684
rect 165513 -712 165547 -684
rect 165575 -712 165609 -684
rect 165637 -712 165671 -684
rect 165699 -712 165747 -684
rect 165437 -746 165747 -712
rect 165437 -774 165485 -746
rect 165513 -774 165547 -746
rect 165575 -774 165609 -746
rect 165637 -774 165671 -746
rect 165699 -774 165747 -746
rect 165437 -822 165747 -774
rect 172577 298606 172887 299134
rect 172577 298578 172625 298606
rect 172653 298578 172687 298606
rect 172715 298578 172749 298606
rect 172777 298578 172811 298606
rect 172839 298578 172887 298606
rect 172577 298544 172887 298578
rect 172577 298516 172625 298544
rect 172653 298516 172687 298544
rect 172715 298516 172749 298544
rect 172777 298516 172811 298544
rect 172839 298516 172887 298544
rect 172577 298482 172887 298516
rect 172577 298454 172625 298482
rect 172653 298454 172687 298482
rect 172715 298454 172749 298482
rect 172777 298454 172811 298482
rect 172839 298454 172887 298482
rect 172577 298420 172887 298454
rect 172577 298392 172625 298420
rect 172653 298392 172687 298420
rect 172715 298392 172749 298420
rect 172777 298392 172811 298420
rect 172839 298392 172887 298420
rect 172577 290175 172887 298392
rect 172577 290147 172625 290175
rect 172653 290147 172687 290175
rect 172715 290147 172749 290175
rect 172777 290147 172811 290175
rect 172839 290147 172887 290175
rect 172577 290113 172887 290147
rect 172577 290085 172625 290113
rect 172653 290085 172687 290113
rect 172715 290085 172749 290113
rect 172777 290085 172811 290113
rect 172839 290085 172887 290113
rect 172577 290051 172887 290085
rect 172577 290023 172625 290051
rect 172653 290023 172687 290051
rect 172715 290023 172749 290051
rect 172777 290023 172811 290051
rect 172839 290023 172887 290051
rect 172577 289989 172887 290023
rect 172577 289961 172625 289989
rect 172653 289961 172687 289989
rect 172715 289961 172749 289989
rect 172777 289961 172811 289989
rect 172839 289961 172887 289989
rect 172577 281175 172887 289961
rect 172577 281147 172625 281175
rect 172653 281147 172687 281175
rect 172715 281147 172749 281175
rect 172777 281147 172811 281175
rect 172839 281147 172887 281175
rect 172577 281113 172887 281147
rect 172577 281085 172625 281113
rect 172653 281085 172687 281113
rect 172715 281085 172749 281113
rect 172777 281085 172811 281113
rect 172839 281085 172887 281113
rect 172577 281051 172887 281085
rect 172577 281023 172625 281051
rect 172653 281023 172687 281051
rect 172715 281023 172749 281051
rect 172777 281023 172811 281051
rect 172839 281023 172887 281051
rect 172577 280989 172887 281023
rect 172577 280961 172625 280989
rect 172653 280961 172687 280989
rect 172715 280961 172749 280989
rect 172777 280961 172811 280989
rect 172839 280961 172887 280989
rect 172577 272175 172887 280961
rect 172577 272147 172625 272175
rect 172653 272147 172687 272175
rect 172715 272147 172749 272175
rect 172777 272147 172811 272175
rect 172839 272147 172887 272175
rect 172577 272113 172887 272147
rect 172577 272085 172625 272113
rect 172653 272085 172687 272113
rect 172715 272085 172749 272113
rect 172777 272085 172811 272113
rect 172839 272085 172887 272113
rect 172577 272051 172887 272085
rect 172577 272023 172625 272051
rect 172653 272023 172687 272051
rect 172715 272023 172749 272051
rect 172777 272023 172811 272051
rect 172839 272023 172887 272051
rect 172577 271989 172887 272023
rect 172577 271961 172625 271989
rect 172653 271961 172687 271989
rect 172715 271961 172749 271989
rect 172777 271961 172811 271989
rect 172839 271961 172887 271989
rect 172577 263175 172887 271961
rect 172577 263147 172625 263175
rect 172653 263147 172687 263175
rect 172715 263147 172749 263175
rect 172777 263147 172811 263175
rect 172839 263147 172887 263175
rect 172577 263113 172887 263147
rect 172577 263085 172625 263113
rect 172653 263085 172687 263113
rect 172715 263085 172749 263113
rect 172777 263085 172811 263113
rect 172839 263085 172887 263113
rect 172577 263051 172887 263085
rect 172577 263023 172625 263051
rect 172653 263023 172687 263051
rect 172715 263023 172749 263051
rect 172777 263023 172811 263051
rect 172839 263023 172887 263051
rect 172577 262989 172887 263023
rect 172577 262961 172625 262989
rect 172653 262961 172687 262989
rect 172715 262961 172749 262989
rect 172777 262961 172811 262989
rect 172839 262961 172887 262989
rect 172577 254175 172887 262961
rect 172577 254147 172625 254175
rect 172653 254147 172687 254175
rect 172715 254147 172749 254175
rect 172777 254147 172811 254175
rect 172839 254147 172887 254175
rect 172577 254113 172887 254147
rect 172577 254085 172625 254113
rect 172653 254085 172687 254113
rect 172715 254085 172749 254113
rect 172777 254085 172811 254113
rect 172839 254085 172887 254113
rect 172577 254051 172887 254085
rect 172577 254023 172625 254051
rect 172653 254023 172687 254051
rect 172715 254023 172749 254051
rect 172777 254023 172811 254051
rect 172839 254023 172887 254051
rect 172577 253989 172887 254023
rect 172577 253961 172625 253989
rect 172653 253961 172687 253989
rect 172715 253961 172749 253989
rect 172777 253961 172811 253989
rect 172839 253961 172887 253989
rect 172577 245175 172887 253961
rect 172577 245147 172625 245175
rect 172653 245147 172687 245175
rect 172715 245147 172749 245175
rect 172777 245147 172811 245175
rect 172839 245147 172887 245175
rect 172577 245113 172887 245147
rect 172577 245085 172625 245113
rect 172653 245085 172687 245113
rect 172715 245085 172749 245113
rect 172777 245085 172811 245113
rect 172839 245085 172887 245113
rect 172577 245051 172887 245085
rect 172577 245023 172625 245051
rect 172653 245023 172687 245051
rect 172715 245023 172749 245051
rect 172777 245023 172811 245051
rect 172839 245023 172887 245051
rect 172577 244989 172887 245023
rect 172577 244961 172625 244989
rect 172653 244961 172687 244989
rect 172715 244961 172749 244989
rect 172777 244961 172811 244989
rect 172839 244961 172887 244989
rect 172577 236175 172887 244961
rect 172577 236147 172625 236175
rect 172653 236147 172687 236175
rect 172715 236147 172749 236175
rect 172777 236147 172811 236175
rect 172839 236147 172887 236175
rect 172577 236113 172887 236147
rect 172577 236085 172625 236113
rect 172653 236085 172687 236113
rect 172715 236085 172749 236113
rect 172777 236085 172811 236113
rect 172839 236085 172887 236113
rect 172577 236051 172887 236085
rect 172577 236023 172625 236051
rect 172653 236023 172687 236051
rect 172715 236023 172749 236051
rect 172777 236023 172811 236051
rect 172839 236023 172887 236051
rect 172577 235989 172887 236023
rect 172577 235961 172625 235989
rect 172653 235961 172687 235989
rect 172715 235961 172749 235989
rect 172777 235961 172811 235989
rect 172839 235961 172887 235989
rect 172577 227175 172887 235961
rect 172577 227147 172625 227175
rect 172653 227147 172687 227175
rect 172715 227147 172749 227175
rect 172777 227147 172811 227175
rect 172839 227147 172887 227175
rect 172577 227113 172887 227147
rect 172577 227085 172625 227113
rect 172653 227085 172687 227113
rect 172715 227085 172749 227113
rect 172777 227085 172811 227113
rect 172839 227085 172887 227113
rect 172577 227051 172887 227085
rect 172577 227023 172625 227051
rect 172653 227023 172687 227051
rect 172715 227023 172749 227051
rect 172777 227023 172811 227051
rect 172839 227023 172887 227051
rect 172577 226989 172887 227023
rect 172577 226961 172625 226989
rect 172653 226961 172687 226989
rect 172715 226961 172749 226989
rect 172777 226961 172811 226989
rect 172839 226961 172887 226989
rect 172577 218175 172887 226961
rect 172577 218147 172625 218175
rect 172653 218147 172687 218175
rect 172715 218147 172749 218175
rect 172777 218147 172811 218175
rect 172839 218147 172887 218175
rect 172577 218113 172887 218147
rect 172577 218085 172625 218113
rect 172653 218085 172687 218113
rect 172715 218085 172749 218113
rect 172777 218085 172811 218113
rect 172839 218085 172887 218113
rect 172577 218051 172887 218085
rect 172577 218023 172625 218051
rect 172653 218023 172687 218051
rect 172715 218023 172749 218051
rect 172777 218023 172811 218051
rect 172839 218023 172887 218051
rect 172577 217989 172887 218023
rect 172577 217961 172625 217989
rect 172653 217961 172687 217989
rect 172715 217961 172749 217989
rect 172777 217961 172811 217989
rect 172839 217961 172887 217989
rect 172577 209175 172887 217961
rect 172577 209147 172625 209175
rect 172653 209147 172687 209175
rect 172715 209147 172749 209175
rect 172777 209147 172811 209175
rect 172839 209147 172887 209175
rect 172577 209113 172887 209147
rect 172577 209085 172625 209113
rect 172653 209085 172687 209113
rect 172715 209085 172749 209113
rect 172777 209085 172811 209113
rect 172839 209085 172887 209113
rect 172577 209051 172887 209085
rect 172577 209023 172625 209051
rect 172653 209023 172687 209051
rect 172715 209023 172749 209051
rect 172777 209023 172811 209051
rect 172839 209023 172887 209051
rect 172577 208989 172887 209023
rect 172577 208961 172625 208989
rect 172653 208961 172687 208989
rect 172715 208961 172749 208989
rect 172777 208961 172811 208989
rect 172839 208961 172887 208989
rect 172577 200175 172887 208961
rect 172577 200147 172625 200175
rect 172653 200147 172687 200175
rect 172715 200147 172749 200175
rect 172777 200147 172811 200175
rect 172839 200147 172887 200175
rect 172577 200113 172887 200147
rect 172577 200085 172625 200113
rect 172653 200085 172687 200113
rect 172715 200085 172749 200113
rect 172777 200085 172811 200113
rect 172839 200085 172887 200113
rect 172577 200051 172887 200085
rect 172577 200023 172625 200051
rect 172653 200023 172687 200051
rect 172715 200023 172749 200051
rect 172777 200023 172811 200051
rect 172839 200023 172887 200051
rect 172577 199989 172887 200023
rect 172577 199961 172625 199989
rect 172653 199961 172687 199989
rect 172715 199961 172749 199989
rect 172777 199961 172811 199989
rect 172839 199961 172887 199989
rect 172577 191175 172887 199961
rect 172577 191147 172625 191175
rect 172653 191147 172687 191175
rect 172715 191147 172749 191175
rect 172777 191147 172811 191175
rect 172839 191147 172887 191175
rect 172577 191113 172887 191147
rect 172577 191085 172625 191113
rect 172653 191085 172687 191113
rect 172715 191085 172749 191113
rect 172777 191085 172811 191113
rect 172839 191085 172887 191113
rect 172577 191051 172887 191085
rect 172577 191023 172625 191051
rect 172653 191023 172687 191051
rect 172715 191023 172749 191051
rect 172777 191023 172811 191051
rect 172839 191023 172887 191051
rect 172577 190989 172887 191023
rect 172577 190961 172625 190989
rect 172653 190961 172687 190989
rect 172715 190961 172749 190989
rect 172777 190961 172811 190989
rect 172839 190961 172887 190989
rect 172577 182175 172887 190961
rect 172577 182147 172625 182175
rect 172653 182147 172687 182175
rect 172715 182147 172749 182175
rect 172777 182147 172811 182175
rect 172839 182147 172887 182175
rect 172577 182113 172887 182147
rect 172577 182085 172625 182113
rect 172653 182085 172687 182113
rect 172715 182085 172749 182113
rect 172777 182085 172811 182113
rect 172839 182085 172887 182113
rect 172577 182051 172887 182085
rect 172577 182023 172625 182051
rect 172653 182023 172687 182051
rect 172715 182023 172749 182051
rect 172777 182023 172811 182051
rect 172839 182023 172887 182051
rect 172577 181989 172887 182023
rect 172577 181961 172625 181989
rect 172653 181961 172687 181989
rect 172715 181961 172749 181989
rect 172777 181961 172811 181989
rect 172839 181961 172887 181989
rect 172577 173175 172887 181961
rect 172577 173147 172625 173175
rect 172653 173147 172687 173175
rect 172715 173147 172749 173175
rect 172777 173147 172811 173175
rect 172839 173147 172887 173175
rect 172577 173113 172887 173147
rect 172577 173085 172625 173113
rect 172653 173085 172687 173113
rect 172715 173085 172749 173113
rect 172777 173085 172811 173113
rect 172839 173085 172887 173113
rect 172577 173051 172887 173085
rect 172577 173023 172625 173051
rect 172653 173023 172687 173051
rect 172715 173023 172749 173051
rect 172777 173023 172811 173051
rect 172839 173023 172887 173051
rect 172577 172989 172887 173023
rect 172577 172961 172625 172989
rect 172653 172961 172687 172989
rect 172715 172961 172749 172989
rect 172777 172961 172811 172989
rect 172839 172961 172887 172989
rect 172577 164175 172887 172961
rect 172577 164147 172625 164175
rect 172653 164147 172687 164175
rect 172715 164147 172749 164175
rect 172777 164147 172811 164175
rect 172839 164147 172887 164175
rect 172577 164113 172887 164147
rect 172577 164085 172625 164113
rect 172653 164085 172687 164113
rect 172715 164085 172749 164113
rect 172777 164085 172811 164113
rect 172839 164085 172887 164113
rect 172577 164051 172887 164085
rect 172577 164023 172625 164051
rect 172653 164023 172687 164051
rect 172715 164023 172749 164051
rect 172777 164023 172811 164051
rect 172839 164023 172887 164051
rect 172577 163989 172887 164023
rect 172577 163961 172625 163989
rect 172653 163961 172687 163989
rect 172715 163961 172749 163989
rect 172777 163961 172811 163989
rect 172839 163961 172887 163989
rect 172577 155175 172887 163961
rect 172577 155147 172625 155175
rect 172653 155147 172687 155175
rect 172715 155147 172749 155175
rect 172777 155147 172811 155175
rect 172839 155147 172887 155175
rect 172577 155113 172887 155147
rect 172577 155085 172625 155113
rect 172653 155085 172687 155113
rect 172715 155085 172749 155113
rect 172777 155085 172811 155113
rect 172839 155085 172887 155113
rect 172577 155051 172887 155085
rect 172577 155023 172625 155051
rect 172653 155023 172687 155051
rect 172715 155023 172749 155051
rect 172777 155023 172811 155051
rect 172839 155023 172887 155051
rect 172577 154989 172887 155023
rect 172577 154961 172625 154989
rect 172653 154961 172687 154989
rect 172715 154961 172749 154989
rect 172777 154961 172811 154989
rect 172839 154961 172887 154989
rect 172577 146175 172887 154961
rect 172577 146147 172625 146175
rect 172653 146147 172687 146175
rect 172715 146147 172749 146175
rect 172777 146147 172811 146175
rect 172839 146147 172887 146175
rect 172577 146113 172887 146147
rect 172577 146085 172625 146113
rect 172653 146085 172687 146113
rect 172715 146085 172749 146113
rect 172777 146085 172811 146113
rect 172839 146085 172887 146113
rect 172577 146051 172887 146085
rect 172577 146023 172625 146051
rect 172653 146023 172687 146051
rect 172715 146023 172749 146051
rect 172777 146023 172811 146051
rect 172839 146023 172887 146051
rect 172577 145989 172887 146023
rect 172577 145961 172625 145989
rect 172653 145961 172687 145989
rect 172715 145961 172749 145989
rect 172777 145961 172811 145989
rect 172839 145961 172887 145989
rect 172577 137175 172887 145961
rect 172577 137147 172625 137175
rect 172653 137147 172687 137175
rect 172715 137147 172749 137175
rect 172777 137147 172811 137175
rect 172839 137147 172887 137175
rect 172577 137113 172887 137147
rect 172577 137085 172625 137113
rect 172653 137085 172687 137113
rect 172715 137085 172749 137113
rect 172777 137085 172811 137113
rect 172839 137085 172887 137113
rect 172577 137051 172887 137085
rect 172577 137023 172625 137051
rect 172653 137023 172687 137051
rect 172715 137023 172749 137051
rect 172777 137023 172811 137051
rect 172839 137023 172887 137051
rect 172577 136989 172887 137023
rect 172577 136961 172625 136989
rect 172653 136961 172687 136989
rect 172715 136961 172749 136989
rect 172777 136961 172811 136989
rect 172839 136961 172887 136989
rect 172577 128175 172887 136961
rect 172577 128147 172625 128175
rect 172653 128147 172687 128175
rect 172715 128147 172749 128175
rect 172777 128147 172811 128175
rect 172839 128147 172887 128175
rect 172577 128113 172887 128147
rect 172577 128085 172625 128113
rect 172653 128085 172687 128113
rect 172715 128085 172749 128113
rect 172777 128085 172811 128113
rect 172839 128085 172887 128113
rect 172577 128051 172887 128085
rect 172577 128023 172625 128051
rect 172653 128023 172687 128051
rect 172715 128023 172749 128051
rect 172777 128023 172811 128051
rect 172839 128023 172887 128051
rect 172577 127989 172887 128023
rect 172577 127961 172625 127989
rect 172653 127961 172687 127989
rect 172715 127961 172749 127989
rect 172777 127961 172811 127989
rect 172839 127961 172887 127989
rect 172577 119175 172887 127961
rect 172577 119147 172625 119175
rect 172653 119147 172687 119175
rect 172715 119147 172749 119175
rect 172777 119147 172811 119175
rect 172839 119147 172887 119175
rect 172577 119113 172887 119147
rect 172577 119085 172625 119113
rect 172653 119085 172687 119113
rect 172715 119085 172749 119113
rect 172777 119085 172811 119113
rect 172839 119085 172887 119113
rect 172577 119051 172887 119085
rect 172577 119023 172625 119051
rect 172653 119023 172687 119051
rect 172715 119023 172749 119051
rect 172777 119023 172811 119051
rect 172839 119023 172887 119051
rect 172577 118989 172887 119023
rect 172577 118961 172625 118989
rect 172653 118961 172687 118989
rect 172715 118961 172749 118989
rect 172777 118961 172811 118989
rect 172839 118961 172887 118989
rect 172577 110175 172887 118961
rect 172577 110147 172625 110175
rect 172653 110147 172687 110175
rect 172715 110147 172749 110175
rect 172777 110147 172811 110175
rect 172839 110147 172887 110175
rect 172577 110113 172887 110147
rect 172577 110085 172625 110113
rect 172653 110085 172687 110113
rect 172715 110085 172749 110113
rect 172777 110085 172811 110113
rect 172839 110085 172887 110113
rect 172577 110051 172887 110085
rect 172577 110023 172625 110051
rect 172653 110023 172687 110051
rect 172715 110023 172749 110051
rect 172777 110023 172811 110051
rect 172839 110023 172887 110051
rect 172577 109989 172887 110023
rect 172577 109961 172625 109989
rect 172653 109961 172687 109989
rect 172715 109961 172749 109989
rect 172777 109961 172811 109989
rect 172839 109961 172887 109989
rect 172577 101175 172887 109961
rect 172577 101147 172625 101175
rect 172653 101147 172687 101175
rect 172715 101147 172749 101175
rect 172777 101147 172811 101175
rect 172839 101147 172887 101175
rect 172577 101113 172887 101147
rect 172577 101085 172625 101113
rect 172653 101085 172687 101113
rect 172715 101085 172749 101113
rect 172777 101085 172811 101113
rect 172839 101085 172887 101113
rect 172577 101051 172887 101085
rect 172577 101023 172625 101051
rect 172653 101023 172687 101051
rect 172715 101023 172749 101051
rect 172777 101023 172811 101051
rect 172839 101023 172887 101051
rect 172577 100989 172887 101023
rect 172577 100961 172625 100989
rect 172653 100961 172687 100989
rect 172715 100961 172749 100989
rect 172777 100961 172811 100989
rect 172839 100961 172887 100989
rect 172577 92175 172887 100961
rect 172577 92147 172625 92175
rect 172653 92147 172687 92175
rect 172715 92147 172749 92175
rect 172777 92147 172811 92175
rect 172839 92147 172887 92175
rect 172577 92113 172887 92147
rect 172577 92085 172625 92113
rect 172653 92085 172687 92113
rect 172715 92085 172749 92113
rect 172777 92085 172811 92113
rect 172839 92085 172887 92113
rect 172577 92051 172887 92085
rect 172577 92023 172625 92051
rect 172653 92023 172687 92051
rect 172715 92023 172749 92051
rect 172777 92023 172811 92051
rect 172839 92023 172887 92051
rect 172577 91989 172887 92023
rect 172577 91961 172625 91989
rect 172653 91961 172687 91989
rect 172715 91961 172749 91989
rect 172777 91961 172811 91989
rect 172839 91961 172887 91989
rect 172577 83175 172887 91961
rect 172577 83147 172625 83175
rect 172653 83147 172687 83175
rect 172715 83147 172749 83175
rect 172777 83147 172811 83175
rect 172839 83147 172887 83175
rect 172577 83113 172887 83147
rect 172577 83085 172625 83113
rect 172653 83085 172687 83113
rect 172715 83085 172749 83113
rect 172777 83085 172811 83113
rect 172839 83085 172887 83113
rect 172577 83051 172887 83085
rect 172577 83023 172625 83051
rect 172653 83023 172687 83051
rect 172715 83023 172749 83051
rect 172777 83023 172811 83051
rect 172839 83023 172887 83051
rect 172577 82989 172887 83023
rect 172577 82961 172625 82989
rect 172653 82961 172687 82989
rect 172715 82961 172749 82989
rect 172777 82961 172811 82989
rect 172839 82961 172887 82989
rect 172577 74175 172887 82961
rect 172577 74147 172625 74175
rect 172653 74147 172687 74175
rect 172715 74147 172749 74175
rect 172777 74147 172811 74175
rect 172839 74147 172887 74175
rect 172577 74113 172887 74147
rect 172577 74085 172625 74113
rect 172653 74085 172687 74113
rect 172715 74085 172749 74113
rect 172777 74085 172811 74113
rect 172839 74085 172887 74113
rect 172577 74051 172887 74085
rect 172577 74023 172625 74051
rect 172653 74023 172687 74051
rect 172715 74023 172749 74051
rect 172777 74023 172811 74051
rect 172839 74023 172887 74051
rect 172577 73989 172887 74023
rect 172577 73961 172625 73989
rect 172653 73961 172687 73989
rect 172715 73961 172749 73989
rect 172777 73961 172811 73989
rect 172839 73961 172887 73989
rect 172577 65175 172887 73961
rect 172577 65147 172625 65175
rect 172653 65147 172687 65175
rect 172715 65147 172749 65175
rect 172777 65147 172811 65175
rect 172839 65147 172887 65175
rect 172577 65113 172887 65147
rect 172577 65085 172625 65113
rect 172653 65085 172687 65113
rect 172715 65085 172749 65113
rect 172777 65085 172811 65113
rect 172839 65085 172887 65113
rect 172577 65051 172887 65085
rect 172577 65023 172625 65051
rect 172653 65023 172687 65051
rect 172715 65023 172749 65051
rect 172777 65023 172811 65051
rect 172839 65023 172887 65051
rect 172577 64989 172887 65023
rect 172577 64961 172625 64989
rect 172653 64961 172687 64989
rect 172715 64961 172749 64989
rect 172777 64961 172811 64989
rect 172839 64961 172887 64989
rect 172577 56175 172887 64961
rect 172577 56147 172625 56175
rect 172653 56147 172687 56175
rect 172715 56147 172749 56175
rect 172777 56147 172811 56175
rect 172839 56147 172887 56175
rect 172577 56113 172887 56147
rect 172577 56085 172625 56113
rect 172653 56085 172687 56113
rect 172715 56085 172749 56113
rect 172777 56085 172811 56113
rect 172839 56085 172887 56113
rect 172577 56051 172887 56085
rect 172577 56023 172625 56051
rect 172653 56023 172687 56051
rect 172715 56023 172749 56051
rect 172777 56023 172811 56051
rect 172839 56023 172887 56051
rect 172577 55989 172887 56023
rect 172577 55961 172625 55989
rect 172653 55961 172687 55989
rect 172715 55961 172749 55989
rect 172777 55961 172811 55989
rect 172839 55961 172887 55989
rect 172577 47175 172887 55961
rect 172577 47147 172625 47175
rect 172653 47147 172687 47175
rect 172715 47147 172749 47175
rect 172777 47147 172811 47175
rect 172839 47147 172887 47175
rect 172577 47113 172887 47147
rect 172577 47085 172625 47113
rect 172653 47085 172687 47113
rect 172715 47085 172749 47113
rect 172777 47085 172811 47113
rect 172839 47085 172887 47113
rect 172577 47051 172887 47085
rect 172577 47023 172625 47051
rect 172653 47023 172687 47051
rect 172715 47023 172749 47051
rect 172777 47023 172811 47051
rect 172839 47023 172887 47051
rect 172577 46989 172887 47023
rect 172577 46961 172625 46989
rect 172653 46961 172687 46989
rect 172715 46961 172749 46989
rect 172777 46961 172811 46989
rect 172839 46961 172887 46989
rect 172577 38175 172887 46961
rect 172577 38147 172625 38175
rect 172653 38147 172687 38175
rect 172715 38147 172749 38175
rect 172777 38147 172811 38175
rect 172839 38147 172887 38175
rect 172577 38113 172887 38147
rect 172577 38085 172625 38113
rect 172653 38085 172687 38113
rect 172715 38085 172749 38113
rect 172777 38085 172811 38113
rect 172839 38085 172887 38113
rect 172577 38051 172887 38085
rect 172577 38023 172625 38051
rect 172653 38023 172687 38051
rect 172715 38023 172749 38051
rect 172777 38023 172811 38051
rect 172839 38023 172887 38051
rect 172577 37989 172887 38023
rect 172577 37961 172625 37989
rect 172653 37961 172687 37989
rect 172715 37961 172749 37989
rect 172777 37961 172811 37989
rect 172839 37961 172887 37989
rect 172577 29175 172887 37961
rect 172577 29147 172625 29175
rect 172653 29147 172687 29175
rect 172715 29147 172749 29175
rect 172777 29147 172811 29175
rect 172839 29147 172887 29175
rect 172577 29113 172887 29147
rect 172577 29085 172625 29113
rect 172653 29085 172687 29113
rect 172715 29085 172749 29113
rect 172777 29085 172811 29113
rect 172839 29085 172887 29113
rect 172577 29051 172887 29085
rect 172577 29023 172625 29051
rect 172653 29023 172687 29051
rect 172715 29023 172749 29051
rect 172777 29023 172811 29051
rect 172839 29023 172887 29051
rect 172577 28989 172887 29023
rect 172577 28961 172625 28989
rect 172653 28961 172687 28989
rect 172715 28961 172749 28989
rect 172777 28961 172811 28989
rect 172839 28961 172887 28989
rect 172577 20175 172887 28961
rect 172577 20147 172625 20175
rect 172653 20147 172687 20175
rect 172715 20147 172749 20175
rect 172777 20147 172811 20175
rect 172839 20147 172887 20175
rect 172577 20113 172887 20147
rect 172577 20085 172625 20113
rect 172653 20085 172687 20113
rect 172715 20085 172749 20113
rect 172777 20085 172811 20113
rect 172839 20085 172887 20113
rect 172577 20051 172887 20085
rect 172577 20023 172625 20051
rect 172653 20023 172687 20051
rect 172715 20023 172749 20051
rect 172777 20023 172811 20051
rect 172839 20023 172887 20051
rect 172577 19989 172887 20023
rect 172577 19961 172625 19989
rect 172653 19961 172687 19989
rect 172715 19961 172749 19989
rect 172777 19961 172811 19989
rect 172839 19961 172887 19989
rect 172577 11175 172887 19961
rect 172577 11147 172625 11175
rect 172653 11147 172687 11175
rect 172715 11147 172749 11175
rect 172777 11147 172811 11175
rect 172839 11147 172887 11175
rect 172577 11113 172887 11147
rect 172577 11085 172625 11113
rect 172653 11085 172687 11113
rect 172715 11085 172749 11113
rect 172777 11085 172811 11113
rect 172839 11085 172887 11113
rect 172577 11051 172887 11085
rect 172577 11023 172625 11051
rect 172653 11023 172687 11051
rect 172715 11023 172749 11051
rect 172777 11023 172811 11051
rect 172839 11023 172887 11051
rect 172577 10989 172887 11023
rect 172577 10961 172625 10989
rect 172653 10961 172687 10989
rect 172715 10961 172749 10989
rect 172777 10961 172811 10989
rect 172839 10961 172887 10989
rect 172577 2175 172887 10961
rect 172577 2147 172625 2175
rect 172653 2147 172687 2175
rect 172715 2147 172749 2175
rect 172777 2147 172811 2175
rect 172839 2147 172887 2175
rect 172577 2113 172887 2147
rect 172577 2085 172625 2113
rect 172653 2085 172687 2113
rect 172715 2085 172749 2113
rect 172777 2085 172811 2113
rect 172839 2085 172887 2113
rect 172577 2051 172887 2085
rect 172577 2023 172625 2051
rect 172653 2023 172687 2051
rect 172715 2023 172749 2051
rect 172777 2023 172811 2051
rect 172839 2023 172887 2051
rect 172577 1989 172887 2023
rect 172577 1961 172625 1989
rect 172653 1961 172687 1989
rect 172715 1961 172749 1989
rect 172777 1961 172811 1989
rect 172839 1961 172887 1989
rect 172577 -80 172887 1961
rect 172577 -108 172625 -80
rect 172653 -108 172687 -80
rect 172715 -108 172749 -80
rect 172777 -108 172811 -80
rect 172839 -108 172887 -80
rect 172577 -142 172887 -108
rect 172577 -170 172625 -142
rect 172653 -170 172687 -142
rect 172715 -170 172749 -142
rect 172777 -170 172811 -142
rect 172839 -170 172887 -142
rect 172577 -204 172887 -170
rect 172577 -232 172625 -204
rect 172653 -232 172687 -204
rect 172715 -232 172749 -204
rect 172777 -232 172811 -204
rect 172839 -232 172887 -204
rect 172577 -266 172887 -232
rect 172577 -294 172625 -266
rect 172653 -294 172687 -266
rect 172715 -294 172749 -266
rect 172777 -294 172811 -266
rect 172839 -294 172887 -266
rect 172577 -822 172887 -294
rect 174437 299086 174747 299134
rect 174437 299058 174485 299086
rect 174513 299058 174547 299086
rect 174575 299058 174609 299086
rect 174637 299058 174671 299086
rect 174699 299058 174747 299086
rect 174437 299024 174747 299058
rect 174437 298996 174485 299024
rect 174513 298996 174547 299024
rect 174575 298996 174609 299024
rect 174637 298996 174671 299024
rect 174699 298996 174747 299024
rect 174437 298962 174747 298996
rect 174437 298934 174485 298962
rect 174513 298934 174547 298962
rect 174575 298934 174609 298962
rect 174637 298934 174671 298962
rect 174699 298934 174747 298962
rect 174437 298900 174747 298934
rect 174437 298872 174485 298900
rect 174513 298872 174547 298900
rect 174575 298872 174609 298900
rect 174637 298872 174671 298900
rect 174699 298872 174747 298900
rect 174437 293175 174747 298872
rect 174437 293147 174485 293175
rect 174513 293147 174547 293175
rect 174575 293147 174609 293175
rect 174637 293147 174671 293175
rect 174699 293147 174747 293175
rect 174437 293113 174747 293147
rect 174437 293085 174485 293113
rect 174513 293085 174547 293113
rect 174575 293085 174609 293113
rect 174637 293085 174671 293113
rect 174699 293085 174747 293113
rect 174437 293051 174747 293085
rect 174437 293023 174485 293051
rect 174513 293023 174547 293051
rect 174575 293023 174609 293051
rect 174637 293023 174671 293051
rect 174699 293023 174747 293051
rect 174437 292989 174747 293023
rect 174437 292961 174485 292989
rect 174513 292961 174547 292989
rect 174575 292961 174609 292989
rect 174637 292961 174671 292989
rect 174699 292961 174747 292989
rect 174437 284175 174747 292961
rect 174437 284147 174485 284175
rect 174513 284147 174547 284175
rect 174575 284147 174609 284175
rect 174637 284147 174671 284175
rect 174699 284147 174747 284175
rect 174437 284113 174747 284147
rect 174437 284085 174485 284113
rect 174513 284085 174547 284113
rect 174575 284085 174609 284113
rect 174637 284085 174671 284113
rect 174699 284085 174747 284113
rect 174437 284051 174747 284085
rect 174437 284023 174485 284051
rect 174513 284023 174547 284051
rect 174575 284023 174609 284051
rect 174637 284023 174671 284051
rect 174699 284023 174747 284051
rect 174437 283989 174747 284023
rect 174437 283961 174485 283989
rect 174513 283961 174547 283989
rect 174575 283961 174609 283989
rect 174637 283961 174671 283989
rect 174699 283961 174747 283989
rect 174437 275175 174747 283961
rect 174437 275147 174485 275175
rect 174513 275147 174547 275175
rect 174575 275147 174609 275175
rect 174637 275147 174671 275175
rect 174699 275147 174747 275175
rect 174437 275113 174747 275147
rect 174437 275085 174485 275113
rect 174513 275085 174547 275113
rect 174575 275085 174609 275113
rect 174637 275085 174671 275113
rect 174699 275085 174747 275113
rect 174437 275051 174747 275085
rect 174437 275023 174485 275051
rect 174513 275023 174547 275051
rect 174575 275023 174609 275051
rect 174637 275023 174671 275051
rect 174699 275023 174747 275051
rect 174437 274989 174747 275023
rect 174437 274961 174485 274989
rect 174513 274961 174547 274989
rect 174575 274961 174609 274989
rect 174637 274961 174671 274989
rect 174699 274961 174747 274989
rect 174437 266175 174747 274961
rect 174437 266147 174485 266175
rect 174513 266147 174547 266175
rect 174575 266147 174609 266175
rect 174637 266147 174671 266175
rect 174699 266147 174747 266175
rect 174437 266113 174747 266147
rect 174437 266085 174485 266113
rect 174513 266085 174547 266113
rect 174575 266085 174609 266113
rect 174637 266085 174671 266113
rect 174699 266085 174747 266113
rect 174437 266051 174747 266085
rect 174437 266023 174485 266051
rect 174513 266023 174547 266051
rect 174575 266023 174609 266051
rect 174637 266023 174671 266051
rect 174699 266023 174747 266051
rect 174437 265989 174747 266023
rect 174437 265961 174485 265989
rect 174513 265961 174547 265989
rect 174575 265961 174609 265989
rect 174637 265961 174671 265989
rect 174699 265961 174747 265989
rect 174437 257175 174747 265961
rect 174437 257147 174485 257175
rect 174513 257147 174547 257175
rect 174575 257147 174609 257175
rect 174637 257147 174671 257175
rect 174699 257147 174747 257175
rect 174437 257113 174747 257147
rect 174437 257085 174485 257113
rect 174513 257085 174547 257113
rect 174575 257085 174609 257113
rect 174637 257085 174671 257113
rect 174699 257085 174747 257113
rect 174437 257051 174747 257085
rect 174437 257023 174485 257051
rect 174513 257023 174547 257051
rect 174575 257023 174609 257051
rect 174637 257023 174671 257051
rect 174699 257023 174747 257051
rect 174437 256989 174747 257023
rect 174437 256961 174485 256989
rect 174513 256961 174547 256989
rect 174575 256961 174609 256989
rect 174637 256961 174671 256989
rect 174699 256961 174747 256989
rect 174437 248175 174747 256961
rect 174437 248147 174485 248175
rect 174513 248147 174547 248175
rect 174575 248147 174609 248175
rect 174637 248147 174671 248175
rect 174699 248147 174747 248175
rect 174437 248113 174747 248147
rect 174437 248085 174485 248113
rect 174513 248085 174547 248113
rect 174575 248085 174609 248113
rect 174637 248085 174671 248113
rect 174699 248085 174747 248113
rect 174437 248051 174747 248085
rect 174437 248023 174485 248051
rect 174513 248023 174547 248051
rect 174575 248023 174609 248051
rect 174637 248023 174671 248051
rect 174699 248023 174747 248051
rect 174437 247989 174747 248023
rect 174437 247961 174485 247989
rect 174513 247961 174547 247989
rect 174575 247961 174609 247989
rect 174637 247961 174671 247989
rect 174699 247961 174747 247989
rect 174437 239175 174747 247961
rect 174437 239147 174485 239175
rect 174513 239147 174547 239175
rect 174575 239147 174609 239175
rect 174637 239147 174671 239175
rect 174699 239147 174747 239175
rect 174437 239113 174747 239147
rect 174437 239085 174485 239113
rect 174513 239085 174547 239113
rect 174575 239085 174609 239113
rect 174637 239085 174671 239113
rect 174699 239085 174747 239113
rect 174437 239051 174747 239085
rect 174437 239023 174485 239051
rect 174513 239023 174547 239051
rect 174575 239023 174609 239051
rect 174637 239023 174671 239051
rect 174699 239023 174747 239051
rect 174437 238989 174747 239023
rect 174437 238961 174485 238989
rect 174513 238961 174547 238989
rect 174575 238961 174609 238989
rect 174637 238961 174671 238989
rect 174699 238961 174747 238989
rect 174437 230175 174747 238961
rect 174437 230147 174485 230175
rect 174513 230147 174547 230175
rect 174575 230147 174609 230175
rect 174637 230147 174671 230175
rect 174699 230147 174747 230175
rect 174437 230113 174747 230147
rect 174437 230085 174485 230113
rect 174513 230085 174547 230113
rect 174575 230085 174609 230113
rect 174637 230085 174671 230113
rect 174699 230085 174747 230113
rect 174437 230051 174747 230085
rect 174437 230023 174485 230051
rect 174513 230023 174547 230051
rect 174575 230023 174609 230051
rect 174637 230023 174671 230051
rect 174699 230023 174747 230051
rect 174437 229989 174747 230023
rect 174437 229961 174485 229989
rect 174513 229961 174547 229989
rect 174575 229961 174609 229989
rect 174637 229961 174671 229989
rect 174699 229961 174747 229989
rect 174437 221175 174747 229961
rect 174437 221147 174485 221175
rect 174513 221147 174547 221175
rect 174575 221147 174609 221175
rect 174637 221147 174671 221175
rect 174699 221147 174747 221175
rect 174437 221113 174747 221147
rect 174437 221085 174485 221113
rect 174513 221085 174547 221113
rect 174575 221085 174609 221113
rect 174637 221085 174671 221113
rect 174699 221085 174747 221113
rect 174437 221051 174747 221085
rect 174437 221023 174485 221051
rect 174513 221023 174547 221051
rect 174575 221023 174609 221051
rect 174637 221023 174671 221051
rect 174699 221023 174747 221051
rect 174437 220989 174747 221023
rect 174437 220961 174485 220989
rect 174513 220961 174547 220989
rect 174575 220961 174609 220989
rect 174637 220961 174671 220989
rect 174699 220961 174747 220989
rect 174437 212175 174747 220961
rect 174437 212147 174485 212175
rect 174513 212147 174547 212175
rect 174575 212147 174609 212175
rect 174637 212147 174671 212175
rect 174699 212147 174747 212175
rect 174437 212113 174747 212147
rect 174437 212085 174485 212113
rect 174513 212085 174547 212113
rect 174575 212085 174609 212113
rect 174637 212085 174671 212113
rect 174699 212085 174747 212113
rect 174437 212051 174747 212085
rect 174437 212023 174485 212051
rect 174513 212023 174547 212051
rect 174575 212023 174609 212051
rect 174637 212023 174671 212051
rect 174699 212023 174747 212051
rect 174437 211989 174747 212023
rect 174437 211961 174485 211989
rect 174513 211961 174547 211989
rect 174575 211961 174609 211989
rect 174637 211961 174671 211989
rect 174699 211961 174747 211989
rect 174437 203175 174747 211961
rect 174437 203147 174485 203175
rect 174513 203147 174547 203175
rect 174575 203147 174609 203175
rect 174637 203147 174671 203175
rect 174699 203147 174747 203175
rect 174437 203113 174747 203147
rect 174437 203085 174485 203113
rect 174513 203085 174547 203113
rect 174575 203085 174609 203113
rect 174637 203085 174671 203113
rect 174699 203085 174747 203113
rect 174437 203051 174747 203085
rect 174437 203023 174485 203051
rect 174513 203023 174547 203051
rect 174575 203023 174609 203051
rect 174637 203023 174671 203051
rect 174699 203023 174747 203051
rect 174437 202989 174747 203023
rect 174437 202961 174485 202989
rect 174513 202961 174547 202989
rect 174575 202961 174609 202989
rect 174637 202961 174671 202989
rect 174699 202961 174747 202989
rect 174437 194175 174747 202961
rect 174437 194147 174485 194175
rect 174513 194147 174547 194175
rect 174575 194147 174609 194175
rect 174637 194147 174671 194175
rect 174699 194147 174747 194175
rect 174437 194113 174747 194147
rect 174437 194085 174485 194113
rect 174513 194085 174547 194113
rect 174575 194085 174609 194113
rect 174637 194085 174671 194113
rect 174699 194085 174747 194113
rect 174437 194051 174747 194085
rect 174437 194023 174485 194051
rect 174513 194023 174547 194051
rect 174575 194023 174609 194051
rect 174637 194023 174671 194051
rect 174699 194023 174747 194051
rect 174437 193989 174747 194023
rect 174437 193961 174485 193989
rect 174513 193961 174547 193989
rect 174575 193961 174609 193989
rect 174637 193961 174671 193989
rect 174699 193961 174747 193989
rect 174437 185175 174747 193961
rect 174437 185147 174485 185175
rect 174513 185147 174547 185175
rect 174575 185147 174609 185175
rect 174637 185147 174671 185175
rect 174699 185147 174747 185175
rect 174437 185113 174747 185147
rect 174437 185085 174485 185113
rect 174513 185085 174547 185113
rect 174575 185085 174609 185113
rect 174637 185085 174671 185113
rect 174699 185085 174747 185113
rect 174437 185051 174747 185085
rect 174437 185023 174485 185051
rect 174513 185023 174547 185051
rect 174575 185023 174609 185051
rect 174637 185023 174671 185051
rect 174699 185023 174747 185051
rect 174437 184989 174747 185023
rect 174437 184961 174485 184989
rect 174513 184961 174547 184989
rect 174575 184961 174609 184989
rect 174637 184961 174671 184989
rect 174699 184961 174747 184989
rect 174437 176175 174747 184961
rect 174437 176147 174485 176175
rect 174513 176147 174547 176175
rect 174575 176147 174609 176175
rect 174637 176147 174671 176175
rect 174699 176147 174747 176175
rect 174437 176113 174747 176147
rect 174437 176085 174485 176113
rect 174513 176085 174547 176113
rect 174575 176085 174609 176113
rect 174637 176085 174671 176113
rect 174699 176085 174747 176113
rect 174437 176051 174747 176085
rect 174437 176023 174485 176051
rect 174513 176023 174547 176051
rect 174575 176023 174609 176051
rect 174637 176023 174671 176051
rect 174699 176023 174747 176051
rect 174437 175989 174747 176023
rect 174437 175961 174485 175989
rect 174513 175961 174547 175989
rect 174575 175961 174609 175989
rect 174637 175961 174671 175989
rect 174699 175961 174747 175989
rect 174437 167175 174747 175961
rect 174437 167147 174485 167175
rect 174513 167147 174547 167175
rect 174575 167147 174609 167175
rect 174637 167147 174671 167175
rect 174699 167147 174747 167175
rect 174437 167113 174747 167147
rect 174437 167085 174485 167113
rect 174513 167085 174547 167113
rect 174575 167085 174609 167113
rect 174637 167085 174671 167113
rect 174699 167085 174747 167113
rect 174437 167051 174747 167085
rect 174437 167023 174485 167051
rect 174513 167023 174547 167051
rect 174575 167023 174609 167051
rect 174637 167023 174671 167051
rect 174699 167023 174747 167051
rect 174437 166989 174747 167023
rect 174437 166961 174485 166989
rect 174513 166961 174547 166989
rect 174575 166961 174609 166989
rect 174637 166961 174671 166989
rect 174699 166961 174747 166989
rect 174437 158175 174747 166961
rect 174437 158147 174485 158175
rect 174513 158147 174547 158175
rect 174575 158147 174609 158175
rect 174637 158147 174671 158175
rect 174699 158147 174747 158175
rect 174437 158113 174747 158147
rect 174437 158085 174485 158113
rect 174513 158085 174547 158113
rect 174575 158085 174609 158113
rect 174637 158085 174671 158113
rect 174699 158085 174747 158113
rect 174437 158051 174747 158085
rect 174437 158023 174485 158051
rect 174513 158023 174547 158051
rect 174575 158023 174609 158051
rect 174637 158023 174671 158051
rect 174699 158023 174747 158051
rect 174437 157989 174747 158023
rect 174437 157961 174485 157989
rect 174513 157961 174547 157989
rect 174575 157961 174609 157989
rect 174637 157961 174671 157989
rect 174699 157961 174747 157989
rect 174437 149175 174747 157961
rect 174437 149147 174485 149175
rect 174513 149147 174547 149175
rect 174575 149147 174609 149175
rect 174637 149147 174671 149175
rect 174699 149147 174747 149175
rect 174437 149113 174747 149147
rect 174437 149085 174485 149113
rect 174513 149085 174547 149113
rect 174575 149085 174609 149113
rect 174637 149085 174671 149113
rect 174699 149085 174747 149113
rect 174437 149051 174747 149085
rect 174437 149023 174485 149051
rect 174513 149023 174547 149051
rect 174575 149023 174609 149051
rect 174637 149023 174671 149051
rect 174699 149023 174747 149051
rect 174437 148989 174747 149023
rect 174437 148961 174485 148989
rect 174513 148961 174547 148989
rect 174575 148961 174609 148989
rect 174637 148961 174671 148989
rect 174699 148961 174747 148989
rect 174437 140175 174747 148961
rect 174437 140147 174485 140175
rect 174513 140147 174547 140175
rect 174575 140147 174609 140175
rect 174637 140147 174671 140175
rect 174699 140147 174747 140175
rect 174437 140113 174747 140147
rect 174437 140085 174485 140113
rect 174513 140085 174547 140113
rect 174575 140085 174609 140113
rect 174637 140085 174671 140113
rect 174699 140085 174747 140113
rect 174437 140051 174747 140085
rect 174437 140023 174485 140051
rect 174513 140023 174547 140051
rect 174575 140023 174609 140051
rect 174637 140023 174671 140051
rect 174699 140023 174747 140051
rect 174437 139989 174747 140023
rect 174437 139961 174485 139989
rect 174513 139961 174547 139989
rect 174575 139961 174609 139989
rect 174637 139961 174671 139989
rect 174699 139961 174747 139989
rect 174437 131175 174747 139961
rect 174437 131147 174485 131175
rect 174513 131147 174547 131175
rect 174575 131147 174609 131175
rect 174637 131147 174671 131175
rect 174699 131147 174747 131175
rect 174437 131113 174747 131147
rect 174437 131085 174485 131113
rect 174513 131085 174547 131113
rect 174575 131085 174609 131113
rect 174637 131085 174671 131113
rect 174699 131085 174747 131113
rect 174437 131051 174747 131085
rect 174437 131023 174485 131051
rect 174513 131023 174547 131051
rect 174575 131023 174609 131051
rect 174637 131023 174671 131051
rect 174699 131023 174747 131051
rect 174437 130989 174747 131023
rect 174437 130961 174485 130989
rect 174513 130961 174547 130989
rect 174575 130961 174609 130989
rect 174637 130961 174671 130989
rect 174699 130961 174747 130989
rect 174437 122175 174747 130961
rect 174437 122147 174485 122175
rect 174513 122147 174547 122175
rect 174575 122147 174609 122175
rect 174637 122147 174671 122175
rect 174699 122147 174747 122175
rect 174437 122113 174747 122147
rect 174437 122085 174485 122113
rect 174513 122085 174547 122113
rect 174575 122085 174609 122113
rect 174637 122085 174671 122113
rect 174699 122085 174747 122113
rect 174437 122051 174747 122085
rect 174437 122023 174485 122051
rect 174513 122023 174547 122051
rect 174575 122023 174609 122051
rect 174637 122023 174671 122051
rect 174699 122023 174747 122051
rect 174437 121989 174747 122023
rect 174437 121961 174485 121989
rect 174513 121961 174547 121989
rect 174575 121961 174609 121989
rect 174637 121961 174671 121989
rect 174699 121961 174747 121989
rect 174437 113175 174747 121961
rect 174437 113147 174485 113175
rect 174513 113147 174547 113175
rect 174575 113147 174609 113175
rect 174637 113147 174671 113175
rect 174699 113147 174747 113175
rect 174437 113113 174747 113147
rect 174437 113085 174485 113113
rect 174513 113085 174547 113113
rect 174575 113085 174609 113113
rect 174637 113085 174671 113113
rect 174699 113085 174747 113113
rect 174437 113051 174747 113085
rect 174437 113023 174485 113051
rect 174513 113023 174547 113051
rect 174575 113023 174609 113051
rect 174637 113023 174671 113051
rect 174699 113023 174747 113051
rect 174437 112989 174747 113023
rect 174437 112961 174485 112989
rect 174513 112961 174547 112989
rect 174575 112961 174609 112989
rect 174637 112961 174671 112989
rect 174699 112961 174747 112989
rect 174437 104175 174747 112961
rect 174437 104147 174485 104175
rect 174513 104147 174547 104175
rect 174575 104147 174609 104175
rect 174637 104147 174671 104175
rect 174699 104147 174747 104175
rect 174437 104113 174747 104147
rect 174437 104085 174485 104113
rect 174513 104085 174547 104113
rect 174575 104085 174609 104113
rect 174637 104085 174671 104113
rect 174699 104085 174747 104113
rect 174437 104051 174747 104085
rect 174437 104023 174485 104051
rect 174513 104023 174547 104051
rect 174575 104023 174609 104051
rect 174637 104023 174671 104051
rect 174699 104023 174747 104051
rect 174437 103989 174747 104023
rect 174437 103961 174485 103989
rect 174513 103961 174547 103989
rect 174575 103961 174609 103989
rect 174637 103961 174671 103989
rect 174699 103961 174747 103989
rect 174437 95175 174747 103961
rect 174437 95147 174485 95175
rect 174513 95147 174547 95175
rect 174575 95147 174609 95175
rect 174637 95147 174671 95175
rect 174699 95147 174747 95175
rect 174437 95113 174747 95147
rect 174437 95085 174485 95113
rect 174513 95085 174547 95113
rect 174575 95085 174609 95113
rect 174637 95085 174671 95113
rect 174699 95085 174747 95113
rect 174437 95051 174747 95085
rect 174437 95023 174485 95051
rect 174513 95023 174547 95051
rect 174575 95023 174609 95051
rect 174637 95023 174671 95051
rect 174699 95023 174747 95051
rect 174437 94989 174747 95023
rect 174437 94961 174485 94989
rect 174513 94961 174547 94989
rect 174575 94961 174609 94989
rect 174637 94961 174671 94989
rect 174699 94961 174747 94989
rect 174437 86175 174747 94961
rect 174437 86147 174485 86175
rect 174513 86147 174547 86175
rect 174575 86147 174609 86175
rect 174637 86147 174671 86175
rect 174699 86147 174747 86175
rect 174437 86113 174747 86147
rect 174437 86085 174485 86113
rect 174513 86085 174547 86113
rect 174575 86085 174609 86113
rect 174637 86085 174671 86113
rect 174699 86085 174747 86113
rect 174437 86051 174747 86085
rect 174437 86023 174485 86051
rect 174513 86023 174547 86051
rect 174575 86023 174609 86051
rect 174637 86023 174671 86051
rect 174699 86023 174747 86051
rect 174437 85989 174747 86023
rect 174437 85961 174485 85989
rect 174513 85961 174547 85989
rect 174575 85961 174609 85989
rect 174637 85961 174671 85989
rect 174699 85961 174747 85989
rect 174437 77175 174747 85961
rect 174437 77147 174485 77175
rect 174513 77147 174547 77175
rect 174575 77147 174609 77175
rect 174637 77147 174671 77175
rect 174699 77147 174747 77175
rect 174437 77113 174747 77147
rect 174437 77085 174485 77113
rect 174513 77085 174547 77113
rect 174575 77085 174609 77113
rect 174637 77085 174671 77113
rect 174699 77085 174747 77113
rect 174437 77051 174747 77085
rect 174437 77023 174485 77051
rect 174513 77023 174547 77051
rect 174575 77023 174609 77051
rect 174637 77023 174671 77051
rect 174699 77023 174747 77051
rect 174437 76989 174747 77023
rect 174437 76961 174485 76989
rect 174513 76961 174547 76989
rect 174575 76961 174609 76989
rect 174637 76961 174671 76989
rect 174699 76961 174747 76989
rect 174437 68175 174747 76961
rect 174437 68147 174485 68175
rect 174513 68147 174547 68175
rect 174575 68147 174609 68175
rect 174637 68147 174671 68175
rect 174699 68147 174747 68175
rect 174437 68113 174747 68147
rect 174437 68085 174485 68113
rect 174513 68085 174547 68113
rect 174575 68085 174609 68113
rect 174637 68085 174671 68113
rect 174699 68085 174747 68113
rect 174437 68051 174747 68085
rect 174437 68023 174485 68051
rect 174513 68023 174547 68051
rect 174575 68023 174609 68051
rect 174637 68023 174671 68051
rect 174699 68023 174747 68051
rect 174437 67989 174747 68023
rect 174437 67961 174485 67989
rect 174513 67961 174547 67989
rect 174575 67961 174609 67989
rect 174637 67961 174671 67989
rect 174699 67961 174747 67989
rect 174437 59175 174747 67961
rect 174437 59147 174485 59175
rect 174513 59147 174547 59175
rect 174575 59147 174609 59175
rect 174637 59147 174671 59175
rect 174699 59147 174747 59175
rect 174437 59113 174747 59147
rect 174437 59085 174485 59113
rect 174513 59085 174547 59113
rect 174575 59085 174609 59113
rect 174637 59085 174671 59113
rect 174699 59085 174747 59113
rect 174437 59051 174747 59085
rect 174437 59023 174485 59051
rect 174513 59023 174547 59051
rect 174575 59023 174609 59051
rect 174637 59023 174671 59051
rect 174699 59023 174747 59051
rect 174437 58989 174747 59023
rect 174437 58961 174485 58989
rect 174513 58961 174547 58989
rect 174575 58961 174609 58989
rect 174637 58961 174671 58989
rect 174699 58961 174747 58989
rect 174437 50175 174747 58961
rect 174437 50147 174485 50175
rect 174513 50147 174547 50175
rect 174575 50147 174609 50175
rect 174637 50147 174671 50175
rect 174699 50147 174747 50175
rect 174437 50113 174747 50147
rect 174437 50085 174485 50113
rect 174513 50085 174547 50113
rect 174575 50085 174609 50113
rect 174637 50085 174671 50113
rect 174699 50085 174747 50113
rect 174437 50051 174747 50085
rect 174437 50023 174485 50051
rect 174513 50023 174547 50051
rect 174575 50023 174609 50051
rect 174637 50023 174671 50051
rect 174699 50023 174747 50051
rect 174437 49989 174747 50023
rect 174437 49961 174485 49989
rect 174513 49961 174547 49989
rect 174575 49961 174609 49989
rect 174637 49961 174671 49989
rect 174699 49961 174747 49989
rect 174437 41175 174747 49961
rect 174437 41147 174485 41175
rect 174513 41147 174547 41175
rect 174575 41147 174609 41175
rect 174637 41147 174671 41175
rect 174699 41147 174747 41175
rect 174437 41113 174747 41147
rect 174437 41085 174485 41113
rect 174513 41085 174547 41113
rect 174575 41085 174609 41113
rect 174637 41085 174671 41113
rect 174699 41085 174747 41113
rect 174437 41051 174747 41085
rect 174437 41023 174485 41051
rect 174513 41023 174547 41051
rect 174575 41023 174609 41051
rect 174637 41023 174671 41051
rect 174699 41023 174747 41051
rect 174437 40989 174747 41023
rect 174437 40961 174485 40989
rect 174513 40961 174547 40989
rect 174575 40961 174609 40989
rect 174637 40961 174671 40989
rect 174699 40961 174747 40989
rect 174437 32175 174747 40961
rect 174437 32147 174485 32175
rect 174513 32147 174547 32175
rect 174575 32147 174609 32175
rect 174637 32147 174671 32175
rect 174699 32147 174747 32175
rect 174437 32113 174747 32147
rect 174437 32085 174485 32113
rect 174513 32085 174547 32113
rect 174575 32085 174609 32113
rect 174637 32085 174671 32113
rect 174699 32085 174747 32113
rect 174437 32051 174747 32085
rect 174437 32023 174485 32051
rect 174513 32023 174547 32051
rect 174575 32023 174609 32051
rect 174637 32023 174671 32051
rect 174699 32023 174747 32051
rect 174437 31989 174747 32023
rect 174437 31961 174485 31989
rect 174513 31961 174547 31989
rect 174575 31961 174609 31989
rect 174637 31961 174671 31989
rect 174699 31961 174747 31989
rect 174437 23175 174747 31961
rect 174437 23147 174485 23175
rect 174513 23147 174547 23175
rect 174575 23147 174609 23175
rect 174637 23147 174671 23175
rect 174699 23147 174747 23175
rect 174437 23113 174747 23147
rect 174437 23085 174485 23113
rect 174513 23085 174547 23113
rect 174575 23085 174609 23113
rect 174637 23085 174671 23113
rect 174699 23085 174747 23113
rect 174437 23051 174747 23085
rect 174437 23023 174485 23051
rect 174513 23023 174547 23051
rect 174575 23023 174609 23051
rect 174637 23023 174671 23051
rect 174699 23023 174747 23051
rect 174437 22989 174747 23023
rect 174437 22961 174485 22989
rect 174513 22961 174547 22989
rect 174575 22961 174609 22989
rect 174637 22961 174671 22989
rect 174699 22961 174747 22989
rect 174437 14175 174747 22961
rect 174437 14147 174485 14175
rect 174513 14147 174547 14175
rect 174575 14147 174609 14175
rect 174637 14147 174671 14175
rect 174699 14147 174747 14175
rect 174437 14113 174747 14147
rect 174437 14085 174485 14113
rect 174513 14085 174547 14113
rect 174575 14085 174609 14113
rect 174637 14085 174671 14113
rect 174699 14085 174747 14113
rect 174437 14051 174747 14085
rect 174437 14023 174485 14051
rect 174513 14023 174547 14051
rect 174575 14023 174609 14051
rect 174637 14023 174671 14051
rect 174699 14023 174747 14051
rect 174437 13989 174747 14023
rect 174437 13961 174485 13989
rect 174513 13961 174547 13989
rect 174575 13961 174609 13989
rect 174637 13961 174671 13989
rect 174699 13961 174747 13989
rect 174437 5175 174747 13961
rect 174437 5147 174485 5175
rect 174513 5147 174547 5175
rect 174575 5147 174609 5175
rect 174637 5147 174671 5175
rect 174699 5147 174747 5175
rect 174437 5113 174747 5147
rect 174437 5085 174485 5113
rect 174513 5085 174547 5113
rect 174575 5085 174609 5113
rect 174637 5085 174671 5113
rect 174699 5085 174747 5113
rect 174437 5051 174747 5085
rect 174437 5023 174485 5051
rect 174513 5023 174547 5051
rect 174575 5023 174609 5051
rect 174637 5023 174671 5051
rect 174699 5023 174747 5051
rect 174437 4989 174747 5023
rect 174437 4961 174485 4989
rect 174513 4961 174547 4989
rect 174575 4961 174609 4989
rect 174637 4961 174671 4989
rect 174699 4961 174747 4989
rect 174437 -560 174747 4961
rect 174437 -588 174485 -560
rect 174513 -588 174547 -560
rect 174575 -588 174609 -560
rect 174637 -588 174671 -560
rect 174699 -588 174747 -560
rect 174437 -622 174747 -588
rect 174437 -650 174485 -622
rect 174513 -650 174547 -622
rect 174575 -650 174609 -622
rect 174637 -650 174671 -622
rect 174699 -650 174747 -622
rect 174437 -684 174747 -650
rect 174437 -712 174485 -684
rect 174513 -712 174547 -684
rect 174575 -712 174609 -684
rect 174637 -712 174671 -684
rect 174699 -712 174747 -684
rect 174437 -746 174747 -712
rect 174437 -774 174485 -746
rect 174513 -774 174547 -746
rect 174575 -774 174609 -746
rect 174637 -774 174671 -746
rect 174699 -774 174747 -746
rect 174437 -822 174747 -774
rect 181577 298606 181887 299134
rect 181577 298578 181625 298606
rect 181653 298578 181687 298606
rect 181715 298578 181749 298606
rect 181777 298578 181811 298606
rect 181839 298578 181887 298606
rect 181577 298544 181887 298578
rect 181577 298516 181625 298544
rect 181653 298516 181687 298544
rect 181715 298516 181749 298544
rect 181777 298516 181811 298544
rect 181839 298516 181887 298544
rect 181577 298482 181887 298516
rect 181577 298454 181625 298482
rect 181653 298454 181687 298482
rect 181715 298454 181749 298482
rect 181777 298454 181811 298482
rect 181839 298454 181887 298482
rect 181577 298420 181887 298454
rect 181577 298392 181625 298420
rect 181653 298392 181687 298420
rect 181715 298392 181749 298420
rect 181777 298392 181811 298420
rect 181839 298392 181887 298420
rect 181577 290175 181887 298392
rect 181577 290147 181625 290175
rect 181653 290147 181687 290175
rect 181715 290147 181749 290175
rect 181777 290147 181811 290175
rect 181839 290147 181887 290175
rect 181577 290113 181887 290147
rect 181577 290085 181625 290113
rect 181653 290085 181687 290113
rect 181715 290085 181749 290113
rect 181777 290085 181811 290113
rect 181839 290085 181887 290113
rect 181577 290051 181887 290085
rect 181577 290023 181625 290051
rect 181653 290023 181687 290051
rect 181715 290023 181749 290051
rect 181777 290023 181811 290051
rect 181839 290023 181887 290051
rect 181577 289989 181887 290023
rect 181577 289961 181625 289989
rect 181653 289961 181687 289989
rect 181715 289961 181749 289989
rect 181777 289961 181811 289989
rect 181839 289961 181887 289989
rect 181577 281175 181887 289961
rect 181577 281147 181625 281175
rect 181653 281147 181687 281175
rect 181715 281147 181749 281175
rect 181777 281147 181811 281175
rect 181839 281147 181887 281175
rect 181577 281113 181887 281147
rect 181577 281085 181625 281113
rect 181653 281085 181687 281113
rect 181715 281085 181749 281113
rect 181777 281085 181811 281113
rect 181839 281085 181887 281113
rect 181577 281051 181887 281085
rect 181577 281023 181625 281051
rect 181653 281023 181687 281051
rect 181715 281023 181749 281051
rect 181777 281023 181811 281051
rect 181839 281023 181887 281051
rect 181577 280989 181887 281023
rect 181577 280961 181625 280989
rect 181653 280961 181687 280989
rect 181715 280961 181749 280989
rect 181777 280961 181811 280989
rect 181839 280961 181887 280989
rect 181577 272175 181887 280961
rect 181577 272147 181625 272175
rect 181653 272147 181687 272175
rect 181715 272147 181749 272175
rect 181777 272147 181811 272175
rect 181839 272147 181887 272175
rect 181577 272113 181887 272147
rect 181577 272085 181625 272113
rect 181653 272085 181687 272113
rect 181715 272085 181749 272113
rect 181777 272085 181811 272113
rect 181839 272085 181887 272113
rect 181577 272051 181887 272085
rect 181577 272023 181625 272051
rect 181653 272023 181687 272051
rect 181715 272023 181749 272051
rect 181777 272023 181811 272051
rect 181839 272023 181887 272051
rect 181577 271989 181887 272023
rect 181577 271961 181625 271989
rect 181653 271961 181687 271989
rect 181715 271961 181749 271989
rect 181777 271961 181811 271989
rect 181839 271961 181887 271989
rect 181577 263175 181887 271961
rect 181577 263147 181625 263175
rect 181653 263147 181687 263175
rect 181715 263147 181749 263175
rect 181777 263147 181811 263175
rect 181839 263147 181887 263175
rect 181577 263113 181887 263147
rect 181577 263085 181625 263113
rect 181653 263085 181687 263113
rect 181715 263085 181749 263113
rect 181777 263085 181811 263113
rect 181839 263085 181887 263113
rect 181577 263051 181887 263085
rect 181577 263023 181625 263051
rect 181653 263023 181687 263051
rect 181715 263023 181749 263051
rect 181777 263023 181811 263051
rect 181839 263023 181887 263051
rect 181577 262989 181887 263023
rect 181577 262961 181625 262989
rect 181653 262961 181687 262989
rect 181715 262961 181749 262989
rect 181777 262961 181811 262989
rect 181839 262961 181887 262989
rect 181577 254175 181887 262961
rect 181577 254147 181625 254175
rect 181653 254147 181687 254175
rect 181715 254147 181749 254175
rect 181777 254147 181811 254175
rect 181839 254147 181887 254175
rect 181577 254113 181887 254147
rect 181577 254085 181625 254113
rect 181653 254085 181687 254113
rect 181715 254085 181749 254113
rect 181777 254085 181811 254113
rect 181839 254085 181887 254113
rect 181577 254051 181887 254085
rect 181577 254023 181625 254051
rect 181653 254023 181687 254051
rect 181715 254023 181749 254051
rect 181777 254023 181811 254051
rect 181839 254023 181887 254051
rect 181577 253989 181887 254023
rect 181577 253961 181625 253989
rect 181653 253961 181687 253989
rect 181715 253961 181749 253989
rect 181777 253961 181811 253989
rect 181839 253961 181887 253989
rect 181577 245175 181887 253961
rect 181577 245147 181625 245175
rect 181653 245147 181687 245175
rect 181715 245147 181749 245175
rect 181777 245147 181811 245175
rect 181839 245147 181887 245175
rect 181577 245113 181887 245147
rect 181577 245085 181625 245113
rect 181653 245085 181687 245113
rect 181715 245085 181749 245113
rect 181777 245085 181811 245113
rect 181839 245085 181887 245113
rect 181577 245051 181887 245085
rect 181577 245023 181625 245051
rect 181653 245023 181687 245051
rect 181715 245023 181749 245051
rect 181777 245023 181811 245051
rect 181839 245023 181887 245051
rect 181577 244989 181887 245023
rect 181577 244961 181625 244989
rect 181653 244961 181687 244989
rect 181715 244961 181749 244989
rect 181777 244961 181811 244989
rect 181839 244961 181887 244989
rect 181577 236175 181887 244961
rect 181577 236147 181625 236175
rect 181653 236147 181687 236175
rect 181715 236147 181749 236175
rect 181777 236147 181811 236175
rect 181839 236147 181887 236175
rect 181577 236113 181887 236147
rect 181577 236085 181625 236113
rect 181653 236085 181687 236113
rect 181715 236085 181749 236113
rect 181777 236085 181811 236113
rect 181839 236085 181887 236113
rect 181577 236051 181887 236085
rect 181577 236023 181625 236051
rect 181653 236023 181687 236051
rect 181715 236023 181749 236051
rect 181777 236023 181811 236051
rect 181839 236023 181887 236051
rect 181577 235989 181887 236023
rect 181577 235961 181625 235989
rect 181653 235961 181687 235989
rect 181715 235961 181749 235989
rect 181777 235961 181811 235989
rect 181839 235961 181887 235989
rect 181577 227175 181887 235961
rect 181577 227147 181625 227175
rect 181653 227147 181687 227175
rect 181715 227147 181749 227175
rect 181777 227147 181811 227175
rect 181839 227147 181887 227175
rect 181577 227113 181887 227147
rect 181577 227085 181625 227113
rect 181653 227085 181687 227113
rect 181715 227085 181749 227113
rect 181777 227085 181811 227113
rect 181839 227085 181887 227113
rect 181577 227051 181887 227085
rect 181577 227023 181625 227051
rect 181653 227023 181687 227051
rect 181715 227023 181749 227051
rect 181777 227023 181811 227051
rect 181839 227023 181887 227051
rect 181577 226989 181887 227023
rect 181577 226961 181625 226989
rect 181653 226961 181687 226989
rect 181715 226961 181749 226989
rect 181777 226961 181811 226989
rect 181839 226961 181887 226989
rect 181577 218175 181887 226961
rect 181577 218147 181625 218175
rect 181653 218147 181687 218175
rect 181715 218147 181749 218175
rect 181777 218147 181811 218175
rect 181839 218147 181887 218175
rect 181577 218113 181887 218147
rect 181577 218085 181625 218113
rect 181653 218085 181687 218113
rect 181715 218085 181749 218113
rect 181777 218085 181811 218113
rect 181839 218085 181887 218113
rect 181577 218051 181887 218085
rect 181577 218023 181625 218051
rect 181653 218023 181687 218051
rect 181715 218023 181749 218051
rect 181777 218023 181811 218051
rect 181839 218023 181887 218051
rect 181577 217989 181887 218023
rect 181577 217961 181625 217989
rect 181653 217961 181687 217989
rect 181715 217961 181749 217989
rect 181777 217961 181811 217989
rect 181839 217961 181887 217989
rect 181577 209175 181887 217961
rect 181577 209147 181625 209175
rect 181653 209147 181687 209175
rect 181715 209147 181749 209175
rect 181777 209147 181811 209175
rect 181839 209147 181887 209175
rect 181577 209113 181887 209147
rect 181577 209085 181625 209113
rect 181653 209085 181687 209113
rect 181715 209085 181749 209113
rect 181777 209085 181811 209113
rect 181839 209085 181887 209113
rect 181577 209051 181887 209085
rect 181577 209023 181625 209051
rect 181653 209023 181687 209051
rect 181715 209023 181749 209051
rect 181777 209023 181811 209051
rect 181839 209023 181887 209051
rect 181577 208989 181887 209023
rect 181577 208961 181625 208989
rect 181653 208961 181687 208989
rect 181715 208961 181749 208989
rect 181777 208961 181811 208989
rect 181839 208961 181887 208989
rect 181577 200175 181887 208961
rect 181577 200147 181625 200175
rect 181653 200147 181687 200175
rect 181715 200147 181749 200175
rect 181777 200147 181811 200175
rect 181839 200147 181887 200175
rect 181577 200113 181887 200147
rect 181577 200085 181625 200113
rect 181653 200085 181687 200113
rect 181715 200085 181749 200113
rect 181777 200085 181811 200113
rect 181839 200085 181887 200113
rect 181577 200051 181887 200085
rect 181577 200023 181625 200051
rect 181653 200023 181687 200051
rect 181715 200023 181749 200051
rect 181777 200023 181811 200051
rect 181839 200023 181887 200051
rect 181577 199989 181887 200023
rect 181577 199961 181625 199989
rect 181653 199961 181687 199989
rect 181715 199961 181749 199989
rect 181777 199961 181811 199989
rect 181839 199961 181887 199989
rect 181577 191175 181887 199961
rect 181577 191147 181625 191175
rect 181653 191147 181687 191175
rect 181715 191147 181749 191175
rect 181777 191147 181811 191175
rect 181839 191147 181887 191175
rect 181577 191113 181887 191147
rect 181577 191085 181625 191113
rect 181653 191085 181687 191113
rect 181715 191085 181749 191113
rect 181777 191085 181811 191113
rect 181839 191085 181887 191113
rect 181577 191051 181887 191085
rect 181577 191023 181625 191051
rect 181653 191023 181687 191051
rect 181715 191023 181749 191051
rect 181777 191023 181811 191051
rect 181839 191023 181887 191051
rect 181577 190989 181887 191023
rect 181577 190961 181625 190989
rect 181653 190961 181687 190989
rect 181715 190961 181749 190989
rect 181777 190961 181811 190989
rect 181839 190961 181887 190989
rect 181577 182175 181887 190961
rect 181577 182147 181625 182175
rect 181653 182147 181687 182175
rect 181715 182147 181749 182175
rect 181777 182147 181811 182175
rect 181839 182147 181887 182175
rect 181577 182113 181887 182147
rect 181577 182085 181625 182113
rect 181653 182085 181687 182113
rect 181715 182085 181749 182113
rect 181777 182085 181811 182113
rect 181839 182085 181887 182113
rect 181577 182051 181887 182085
rect 181577 182023 181625 182051
rect 181653 182023 181687 182051
rect 181715 182023 181749 182051
rect 181777 182023 181811 182051
rect 181839 182023 181887 182051
rect 181577 181989 181887 182023
rect 181577 181961 181625 181989
rect 181653 181961 181687 181989
rect 181715 181961 181749 181989
rect 181777 181961 181811 181989
rect 181839 181961 181887 181989
rect 181577 173175 181887 181961
rect 181577 173147 181625 173175
rect 181653 173147 181687 173175
rect 181715 173147 181749 173175
rect 181777 173147 181811 173175
rect 181839 173147 181887 173175
rect 181577 173113 181887 173147
rect 181577 173085 181625 173113
rect 181653 173085 181687 173113
rect 181715 173085 181749 173113
rect 181777 173085 181811 173113
rect 181839 173085 181887 173113
rect 181577 173051 181887 173085
rect 181577 173023 181625 173051
rect 181653 173023 181687 173051
rect 181715 173023 181749 173051
rect 181777 173023 181811 173051
rect 181839 173023 181887 173051
rect 181577 172989 181887 173023
rect 181577 172961 181625 172989
rect 181653 172961 181687 172989
rect 181715 172961 181749 172989
rect 181777 172961 181811 172989
rect 181839 172961 181887 172989
rect 181577 164175 181887 172961
rect 181577 164147 181625 164175
rect 181653 164147 181687 164175
rect 181715 164147 181749 164175
rect 181777 164147 181811 164175
rect 181839 164147 181887 164175
rect 181577 164113 181887 164147
rect 181577 164085 181625 164113
rect 181653 164085 181687 164113
rect 181715 164085 181749 164113
rect 181777 164085 181811 164113
rect 181839 164085 181887 164113
rect 181577 164051 181887 164085
rect 181577 164023 181625 164051
rect 181653 164023 181687 164051
rect 181715 164023 181749 164051
rect 181777 164023 181811 164051
rect 181839 164023 181887 164051
rect 181577 163989 181887 164023
rect 181577 163961 181625 163989
rect 181653 163961 181687 163989
rect 181715 163961 181749 163989
rect 181777 163961 181811 163989
rect 181839 163961 181887 163989
rect 181577 155175 181887 163961
rect 181577 155147 181625 155175
rect 181653 155147 181687 155175
rect 181715 155147 181749 155175
rect 181777 155147 181811 155175
rect 181839 155147 181887 155175
rect 181577 155113 181887 155147
rect 181577 155085 181625 155113
rect 181653 155085 181687 155113
rect 181715 155085 181749 155113
rect 181777 155085 181811 155113
rect 181839 155085 181887 155113
rect 181577 155051 181887 155085
rect 181577 155023 181625 155051
rect 181653 155023 181687 155051
rect 181715 155023 181749 155051
rect 181777 155023 181811 155051
rect 181839 155023 181887 155051
rect 181577 154989 181887 155023
rect 181577 154961 181625 154989
rect 181653 154961 181687 154989
rect 181715 154961 181749 154989
rect 181777 154961 181811 154989
rect 181839 154961 181887 154989
rect 181577 146175 181887 154961
rect 181577 146147 181625 146175
rect 181653 146147 181687 146175
rect 181715 146147 181749 146175
rect 181777 146147 181811 146175
rect 181839 146147 181887 146175
rect 181577 146113 181887 146147
rect 181577 146085 181625 146113
rect 181653 146085 181687 146113
rect 181715 146085 181749 146113
rect 181777 146085 181811 146113
rect 181839 146085 181887 146113
rect 181577 146051 181887 146085
rect 181577 146023 181625 146051
rect 181653 146023 181687 146051
rect 181715 146023 181749 146051
rect 181777 146023 181811 146051
rect 181839 146023 181887 146051
rect 181577 145989 181887 146023
rect 181577 145961 181625 145989
rect 181653 145961 181687 145989
rect 181715 145961 181749 145989
rect 181777 145961 181811 145989
rect 181839 145961 181887 145989
rect 181577 137175 181887 145961
rect 181577 137147 181625 137175
rect 181653 137147 181687 137175
rect 181715 137147 181749 137175
rect 181777 137147 181811 137175
rect 181839 137147 181887 137175
rect 181577 137113 181887 137147
rect 181577 137085 181625 137113
rect 181653 137085 181687 137113
rect 181715 137085 181749 137113
rect 181777 137085 181811 137113
rect 181839 137085 181887 137113
rect 181577 137051 181887 137085
rect 181577 137023 181625 137051
rect 181653 137023 181687 137051
rect 181715 137023 181749 137051
rect 181777 137023 181811 137051
rect 181839 137023 181887 137051
rect 181577 136989 181887 137023
rect 181577 136961 181625 136989
rect 181653 136961 181687 136989
rect 181715 136961 181749 136989
rect 181777 136961 181811 136989
rect 181839 136961 181887 136989
rect 181577 128175 181887 136961
rect 181577 128147 181625 128175
rect 181653 128147 181687 128175
rect 181715 128147 181749 128175
rect 181777 128147 181811 128175
rect 181839 128147 181887 128175
rect 181577 128113 181887 128147
rect 181577 128085 181625 128113
rect 181653 128085 181687 128113
rect 181715 128085 181749 128113
rect 181777 128085 181811 128113
rect 181839 128085 181887 128113
rect 181577 128051 181887 128085
rect 181577 128023 181625 128051
rect 181653 128023 181687 128051
rect 181715 128023 181749 128051
rect 181777 128023 181811 128051
rect 181839 128023 181887 128051
rect 181577 127989 181887 128023
rect 181577 127961 181625 127989
rect 181653 127961 181687 127989
rect 181715 127961 181749 127989
rect 181777 127961 181811 127989
rect 181839 127961 181887 127989
rect 181577 119175 181887 127961
rect 181577 119147 181625 119175
rect 181653 119147 181687 119175
rect 181715 119147 181749 119175
rect 181777 119147 181811 119175
rect 181839 119147 181887 119175
rect 181577 119113 181887 119147
rect 181577 119085 181625 119113
rect 181653 119085 181687 119113
rect 181715 119085 181749 119113
rect 181777 119085 181811 119113
rect 181839 119085 181887 119113
rect 181577 119051 181887 119085
rect 181577 119023 181625 119051
rect 181653 119023 181687 119051
rect 181715 119023 181749 119051
rect 181777 119023 181811 119051
rect 181839 119023 181887 119051
rect 181577 118989 181887 119023
rect 181577 118961 181625 118989
rect 181653 118961 181687 118989
rect 181715 118961 181749 118989
rect 181777 118961 181811 118989
rect 181839 118961 181887 118989
rect 181577 110175 181887 118961
rect 181577 110147 181625 110175
rect 181653 110147 181687 110175
rect 181715 110147 181749 110175
rect 181777 110147 181811 110175
rect 181839 110147 181887 110175
rect 181577 110113 181887 110147
rect 181577 110085 181625 110113
rect 181653 110085 181687 110113
rect 181715 110085 181749 110113
rect 181777 110085 181811 110113
rect 181839 110085 181887 110113
rect 181577 110051 181887 110085
rect 181577 110023 181625 110051
rect 181653 110023 181687 110051
rect 181715 110023 181749 110051
rect 181777 110023 181811 110051
rect 181839 110023 181887 110051
rect 181577 109989 181887 110023
rect 181577 109961 181625 109989
rect 181653 109961 181687 109989
rect 181715 109961 181749 109989
rect 181777 109961 181811 109989
rect 181839 109961 181887 109989
rect 181577 101175 181887 109961
rect 181577 101147 181625 101175
rect 181653 101147 181687 101175
rect 181715 101147 181749 101175
rect 181777 101147 181811 101175
rect 181839 101147 181887 101175
rect 181577 101113 181887 101147
rect 181577 101085 181625 101113
rect 181653 101085 181687 101113
rect 181715 101085 181749 101113
rect 181777 101085 181811 101113
rect 181839 101085 181887 101113
rect 181577 101051 181887 101085
rect 181577 101023 181625 101051
rect 181653 101023 181687 101051
rect 181715 101023 181749 101051
rect 181777 101023 181811 101051
rect 181839 101023 181887 101051
rect 181577 100989 181887 101023
rect 181577 100961 181625 100989
rect 181653 100961 181687 100989
rect 181715 100961 181749 100989
rect 181777 100961 181811 100989
rect 181839 100961 181887 100989
rect 181577 92175 181887 100961
rect 181577 92147 181625 92175
rect 181653 92147 181687 92175
rect 181715 92147 181749 92175
rect 181777 92147 181811 92175
rect 181839 92147 181887 92175
rect 181577 92113 181887 92147
rect 181577 92085 181625 92113
rect 181653 92085 181687 92113
rect 181715 92085 181749 92113
rect 181777 92085 181811 92113
rect 181839 92085 181887 92113
rect 181577 92051 181887 92085
rect 181577 92023 181625 92051
rect 181653 92023 181687 92051
rect 181715 92023 181749 92051
rect 181777 92023 181811 92051
rect 181839 92023 181887 92051
rect 181577 91989 181887 92023
rect 181577 91961 181625 91989
rect 181653 91961 181687 91989
rect 181715 91961 181749 91989
rect 181777 91961 181811 91989
rect 181839 91961 181887 91989
rect 181577 83175 181887 91961
rect 181577 83147 181625 83175
rect 181653 83147 181687 83175
rect 181715 83147 181749 83175
rect 181777 83147 181811 83175
rect 181839 83147 181887 83175
rect 181577 83113 181887 83147
rect 181577 83085 181625 83113
rect 181653 83085 181687 83113
rect 181715 83085 181749 83113
rect 181777 83085 181811 83113
rect 181839 83085 181887 83113
rect 181577 83051 181887 83085
rect 181577 83023 181625 83051
rect 181653 83023 181687 83051
rect 181715 83023 181749 83051
rect 181777 83023 181811 83051
rect 181839 83023 181887 83051
rect 181577 82989 181887 83023
rect 181577 82961 181625 82989
rect 181653 82961 181687 82989
rect 181715 82961 181749 82989
rect 181777 82961 181811 82989
rect 181839 82961 181887 82989
rect 181577 74175 181887 82961
rect 181577 74147 181625 74175
rect 181653 74147 181687 74175
rect 181715 74147 181749 74175
rect 181777 74147 181811 74175
rect 181839 74147 181887 74175
rect 181577 74113 181887 74147
rect 181577 74085 181625 74113
rect 181653 74085 181687 74113
rect 181715 74085 181749 74113
rect 181777 74085 181811 74113
rect 181839 74085 181887 74113
rect 181577 74051 181887 74085
rect 181577 74023 181625 74051
rect 181653 74023 181687 74051
rect 181715 74023 181749 74051
rect 181777 74023 181811 74051
rect 181839 74023 181887 74051
rect 181577 73989 181887 74023
rect 181577 73961 181625 73989
rect 181653 73961 181687 73989
rect 181715 73961 181749 73989
rect 181777 73961 181811 73989
rect 181839 73961 181887 73989
rect 181577 65175 181887 73961
rect 181577 65147 181625 65175
rect 181653 65147 181687 65175
rect 181715 65147 181749 65175
rect 181777 65147 181811 65175
rect 181839 65147 181887 65175
rect 181577 65113 181887 65147
rect 181577 65085 181625 65113
rect 181653 65085 181687 65113
rect 181715 65085 181749 65113
rect 181777 65085 181811 65113
rect 181839 65085 181887 65113
rect 181577 65051 181887 65085
rect 181577 65023 181625 65051
rect 181653 65023 181687 65051
rect 181715 65023 181749 65051
rect 181777 65023 181811 65051
rect 181839 65023 181887 65051
rect 181577 64989 181887 65023
rect 181577 64961 181625 64989
rect 181653 64961 181687 64989
rect 181715 64961 181749 64989
rect 181777 64961 181811 64989
rect 181839 64961 181887 64989
rect 181577 56175 181887 64961
rect 181577 56147 181625 56175
rect 181653 56147 181687 56175
rect 181715 56147 181749 56175
rect 181777 56147 181811 56175
rect 181839 56147 181887 56175
rect 181577 56113 181887 56147
rect 181577 56085 181625 56113
rect 181653 56085 181687 56113
rect 181715 56085 181749 56113
rect 181777 56085 181811 56113
rect 181839 56085 181887 56113
rect 181577 56051 181887 56085
rect 181577 56023 181625 56051
rect 181653 56023 181687 56051
rect 181715 56023 181749 56051
rect 181777 56023 181811 56051
rect 181839 56023 181887 56051
rect 181577 55989 181887 56023
rect 181577 55961 181625 55989
rect 181653 55961 181687 55989
rect 181715 55961 181749 55989
rect 181777 55961 181811 55989
rect 181839 55961 181887 55989
rect 181577 47175 181887 55961
rect 181577 47147 181625 47175
rect 181653 47147 181687 47175
rect 181715 47147 181749 47175
rect 181777 47147 181811 47175
rect 181839 47147 181887 47175
rect 181577 47113 181887 47147
rect 181577 47085 181625 47113
rect 181653 47085 181687 47113
rect 181715 47085 181749 47113
rect 181777 47085 181811 47113
rect 181839 47085 181887 47113
rect 181577 47051 181887 47085
rect 181577 47023 181625 47051
rect 181653 47023 181687 47051
rect 181715 47023 181749 47051
rect 181777 47023 181811 47051
rect 181839 47023 181887 47051
rect 181577 46989 181887 47023
rect 181577 46961 181625 46989
rect 181653 46961 181687 46989
rect 181715 46961 181749 46989
rect 181777 46961 181811 46989
rect 181839 46961 181887 46989
rect 181577 38175 181887 46961
rect 181577 38147 181625 38175
rect 181653 38147 181687 38175
rect 181715 38147 181749 38175
rect 181777 38147 181811 38175
rect 181839 38147 181887 38175
rect 181577 38113 181887 38147
rect 181577 38085 181625 38113
rect 181653 38085 181687 38113
rect 181715 38085 181749 38113
rect 181777 38085 181811 38113
rect 181839 38085 181887 38113
rect 181577 38051 181887 38085
rect 181577 38023 181625 38051
rect 181653 38023 181687 38051
rect 181715 38023 181749 38051
rect 181777 38023 181811 38051
rect 181839 38023 181887 38051
rect 181577 37989 181887 38023
rect 181577 37961 181625 37989
rect 181653 37961 181687 37989
rect 181715 37961 181749 37989
rect 181777 37961 181811 37989
rect 181839 37961 181887 37989
rect 181577 29175 181887 37961
rect 181577 29147 181625 29175
rect 181653 29147 181687 29175
rect 181715 29147 181749 29175
rect 181777 29147 181811 29175
rect 181839 29147 181887 29175
rect 181577 29113 181887 29147
rect 181577 29085 181625 29113
rect 181653 29085 181687 29113
rect 181715 29085 181749 29113
rect 181777 29085 181811 29113
rect 181839 29085 181887 29113
rect 181577 29051 181887 29085
rect 181577 29023 181625 29051
rect 181653 29023 181687 29051
rect 181715 29023 181749 29051
rect 181777 29023 181811 29051
rect 181839 29023 181887 29051
rect 181577 28989 181887 29023
rect 181577 28961 181625 28989
rect 181653 28961 181687 28989
rect 181715 28961 181749 28989
rect 181777 28961 181811 28989
rect 181839 28961 181887 28989
rect 181577 20175 181887 28961
rect 181577 20147 181625 20175
rect 181653 20147 181687 20175
rect 181715 20147 181749 20175
rect 181777 20147 181811 20175
rect 181839 20147 181887 20175
rect 181577 20113 181887 20147
rect 181577 20085 181625 20113
rect 181653 20085 181687 20113
rect 181715 20085 181749 20113
rect 181777 20085 181811 20113
rect 181839 20085 181887 20113
rect 181577 20051 181887 20085
rect 181577 20023 181625 20051
rect 181653 20023 181687 20051
rect 181715 20023 181749 20051
rect 181777 20023 181811 20051
rect 181839 20023 181887 20051
rect 181577 19989 181887 20023
rect 181577 19961 181625 19989
rect 181653 19961 181687 19989
rect 181715 19961 181749 19989
rect 181777 19961 181811 19989
rect 181839 19961 181887 19989
rect 181577 11175 181887 19961
rect 181577 11147 181625 11175
rect 181653 11147 181687 11175
rect 181715 11147 181749 11175
rect 181777 11147 181811 11175
rect 181839 11147 181887 11175
rect 181577 11113 181887 11147
rect 181577 11085 181625 11113
rect 181653 11085 181687 11113
rect 181715 11085 181749 11113
rect 181777 11085 181811 11113
rect 181839 11085 181887 11113
rect 181577 11051 181887 11085
rect 181577 11023 181625 11051
rect 181653 11023 181687 11051
rect 181715 11023 181749 11051
rect 181777 11023 181811 11051
rect 181839 11023 181887 11051
rect 181577 10989 181887 11023
rect 181577 10961 181625 10989
rect 181653 10961 181687 10989
rect 181715 10961 181749 10989
rect 181777 10961 181811 10989
rect 181839 10961 181887 10989
rect 181577 2175 181887 10961
rect 181577 2147 181625 2175
rect 181653 2147 181687 2175
rect 181715 2147 181749 2175
rect 181777 2147 181811 2175
rect 181839 2147 181887 2175
rect 181577 2113 181887 2147
rect 181577 2085 181625 2113
rect 181653 2085 181687 2113
rect 181715 2085 181749 2113
rect 181777 2085 181811 2113
rect 181839 2085 181887 2113
rect 181577 2051 181887 2085
rect 181577 2023 181625 2051
rect 181653 2023 181687 2051
rect 181715 2023 181749 2051
rect 181777 2023 181811 2051
rect 181839 2023 181887 2051
rect 181577 1989 181887 2023
rect 181577 1961 181625 1989
rect 181653 1961 181687 1989
rect 181715 1961 181749 1989
rect 181777 1961 181811 1989
rect 181839 1961 181887 1989
rect 181577 -80 181887 1961
rect 181577 -108 181625 -80
rect 181653 -108 181687 -80
rect 181715 -108 181749 -80
rect 181777 -108 181811 -80
rect 181839 -108 181887 -80
rect 181577 -142 181887 -108
rect 181577 -170 181625 -142
rect 181653 -170 181687 -142
rect 181715 -170 181749 -142
rect 181777 -170 181811 -142
rect 181839 -170 181887 -142
rect 181577 -204 181887 -170
rect 181577 -232 181625 -204
rect 181653 -232 181687 -204
rect 181715 -232 181749 -204
rect 181777 -232 181811 -204
rect 181839 -232 181887 -204
rect 181577 -266 181887 -232
rect 181577 -294 181625 -266
rect 181653 -294 181687 -266
rect 181715 -294 181749 -266
rect 181777 -294 181811 -266
rect 181839 -294 181887 -266
rect 181577 -822 181887 -294
rect 183437 299086 183747 299134
rect 183437 299058 183485 299086
rect 183513 299058 183547 299086
rect 183575 299058 183609 299086
rect 183637 299058 183671 299086
rect 183699 299058 183747 299086
rect 183437 299024 183747 299058
rect 183437 298996 183485 299024
rect 183513 298996 183547 299024
rect 183575 298996 183609 299024
rect 183637 298996 183671 299024
rect 183699 298996 183747 299024
rect 183437 298962 183747 298996
rect 183437 298934 183485 298962
rect 183513 298934 183547 298962
rect 183575 298934 183609 298962
rect 183637 298934 183671 298962
rect 183699 298934 183747 298962
rect 183437 298900 183747 298934
rect 183437 298872 183485 298900
rect 183513 298872 183547 298900
rect 183575 298872 183609 298900
rect 183637 298872 183671 298900
rect 183699 298872 183747 298900
rect 183437 293175 183747 298872
rect 183437 293147 183485 293175
rect 183513 293147 183547 293175
rect 183575 293147 183609 293175
rect 183637 293147 183671 293175
rect 183699 293147 183747 293175
rect 183437 293113 183747 293147
rect 183437 293085 183485 293113
rect 183513 293085 183547 293113
rect 183575 293085 183609 293113
rect 183637 293085 183671 293113
rect 183699 293085 183747 293113
rect 183437 293051 183747 293085
rect 183437 293023 183485 293051
rect 183513 293023 183547 293051
rect 183575 293023 183609 293051
rect 183637 293023 183671 293051
rect 183699 293023 183747 293051
rect 183437 292989 183747 293023
rect 183437 292961 183485 292989
rect 183513 292961 183547 292989
rect 183575 292961 183609 292989
rect 183637 292961 183671 292989
rect 183699 292961 183747 292989
rect 183437 284175 183747 292961
rect 183437 284147 183485 284175
rect 183513 284147 183547 284175
rect 183575 284147 183609 284175
rect 183637 284147 183671 284175
rect 183699 284147 183747 284175
rect 183437 284113 183747 284147
rect 183437 284085 183485 284113
rect 183513 284085 183547 284113
rect 183575 284085 183609 284113
rect 183637 284085 183671 284113
rect 183699 284085 183747 284113
rect 183437 284051 183747 284085
rect 183437 284023 183485 284051
rect 183513 284023 183547 284051
rect 183575 284023 183609 284051
rect 183637 284023 183671 284051
rect 183699 284023 183747 284051
rect 183437 283989 183747 284023
rect 183437 283961 183485 283989
rect 183513 283961 183547 283989
rect 183575 283961 183609 283989
rect 183637 283961 183671 283989
rect 183699 283961 183747 283989
rect 183437 275175 183747 283961
rect 183437 275147 183485 275175
rect 183513 275147 183547 275175
rect 183575 275147 183609 275175
rect 183637 275147 183671 275175
rect 183699 275147 183747 275175
rect 183437 275113 183747 275147
rect 183437 275085 183485 275113
rect 183513 275085 183547 275113
rect 183575 275085 183609 275113
rect 183637 275085 183671 275113
rect 183699 275085 183747 275113
rect 183437 275051 183747 275085
rect 183437 275023 183485 275051
rect 183513 275023 183547 275051
rect 183575 275023 183609 275051
rect 183637 275023 183671 275051
rect 183699 275023 183747 275051
rect 183437 274989 183747 275023
rect 183437 274961 183485 274989
rect 183513 274961 183547 274989
rect 183575 274961 183609 274989
rect 183637 274961 183671 274989
rect 183699 274961 183747 274989
rect 183437 266175 183747 274961
rect 183437 266147 183485 266175
rect 183513 266147 183547 266175
rect 183575 266147 183609 266175
rect 183637 266147 183671 266175
rect 183699 266147 183747 266175
rect 183437 266113 183747 266147
rect 183437 266085 183485 266113
rect 183513 266085 183547 266113
rect 183575 266085 183609 266113
rect 183637 266085 183671 266113
rect 183699 266085 183747 266113
rect 183437 266051 183747 266085
rect 183437 266023 183485 266051
rect 183513 266023 183547 266051
rect 183575 266023 183609 266051
rect 183637 266023 183671 266051
rect 183699 266023 183747 266051
rect 183437 265989 183747 266023
rect 183437 265961 183485 265989
rect 183513 265961 183547 265989
rect 183575 265961 183609 265989
rect 183637 265961 183671 265989
rect 183699 265961 183747 265989
rect 183437 257175 183747 265961
rect 183437 257147 183485 257175
rect 183513 257147 183547 257175
rect 183575 257147 183609 257175
rect 183637 257147 183671 257175
rect 183699 257147 183747 257175
rect 183437 257113 183747 257147
rect 183437 257085 183485 257113
rect 183513 257085 183547 257113
rect 183575 257085 183609 257113
rect 183637 257085 183671 257113
rect 183699 257085 183747 257113
rect 183437 257051 183747 257085
rect 183437 257023 183485 257051
rect 183513 257023 183547 257051
rect 183575 257023 183609 257051
rect 183637 257023 183671 257051
rect 183699 257023 183747 257051
rect 183437 256989 183747 257023
rect 183437 256961 183485 256989
rect 183513 256961 183547 256989
rect 183575 256961 183609 256989
rect 183637 256961 183671 256989
rect 183699 256961 183747 256989
rect 183437 248175 183747 256961
rect 183437 248147 183485 248175
rect 183513 248147 183547 248175
rect 183575 248147 183609 248175
rect 183637 248147 183671 248175
rect 183699 248147 183747 248175
rect 183437 248113 183747 248147
rect 183437 248085 183485 248113
rect 183513 248085 183547 248113
rect 183575 248085 183609 248113
rect 183637 248085 183671 248113
rect 183699 248085 183747 248113
rect 183437 248051 183747 248085
rect 183437 248023 183485 248051
rect 183513 248023 183547 248051
rect 183575 248023 183609 248051
rect 183637 248023 183671 248051
rect 183699 248023 183747 248051
rect 183437 247989 183747 248023
rect 183437 247961 183485 247989
rect 183513 247961 183547 247989
rect 183575 247961 183609 247989
rect 183637 247961 183671 247989
rect 183699 247961 183747 247989
rect 183437 239175 183747 247961
rect 183437 239147 183485 239175
rect 183513 239147 183547 239175
rect 183575 239147 183609 239175
rect 183637 239147 183671 239175
rect 183699 239147 183747 239175
rect 183437 239113 183747 239147
rect 183437 239085 183485 239113
rect 183513 239085 183547 239113
rect 183575 239085 183609 239113
rect 183637 239085 183671 239113
rect 183699 239085 183747 239113
rect 183437 239051 183747 239085
rect 183437 239023 183485 239051
rect 183513 239023 183547 239051
rect 183575 239023 183609 239051
rect 183637 239023 183671 239051
rect 183699 239023 183747 239051
rect 183437 238989 183747 239023
rect 183437 238961 183485 238989
rect 183513 238961 183547 238989
rect 183575 238961 183609 238989
rect 183637 238961 183671 238989
rect 183699 238961 183747 238989
rect 183437 230175 183747 238961
rect 183437 230147 183485 230175
rect 183513 230147 183547 230175
rect 183575 230147 183609 230175
rect 183637 230147 183671 230175
rect 183699 230147 183747 230175
rect 183437 230113 183747 230147
rect 183437 230085 183485 230113
rect 183513 230085 183547 230113
rect 183575 230085 183609 230113
rect 183637 230085 183671 230113
rect 183699 230085 183747 230113
rect 183437 230051 183747 230085
rect 183437 230023 183485 230051
rect 183513 230023 183547 230051
rect 183575 230023 183609 230051
rect 183637 230023 183671 230051
rect 183699 230023 183747 230051
rect 183437 229989 183747 230023
rect 183437 229961 183485 229989
rect 183513 229961 183547 229989
rect 183575 229961 183609 229989
rect 183637 229961 183671 229989
rect 183699 229961 183747 229989
rect 183437 221175 183747 229961
rect 183437 221147 183485 221175
rect 183513 221147 183547 221175
rect 183575 221147 183609 221175
rect 183637 221147 183671 221175
rect 183699 221147 183747 221175
rect 183437 221113 183747 221147
rect 183437 221085 183485 221113
rect 183513 221085 183547 221113
rect 183575 221085 183609 221113
rect 183637 221085 183671 221113
rect 183699 221085 183747 221113
rect 183437 221051 183747 221085
rect 183437 221023 183485 221051
rect 183513 221023 183547 221051
rect 183575 221023 183609 221051
rect 183637 221023 183671 221051
rect 183699 221023 183747 221051
rect 183437 220989 183747 221023
rect 183437 220961 183485 220989
rect 183513 220961 183547 220989
rect 183575 220961 183609 220989
rect 183637 220961 183671 220989
rect 183699 220961 183747 220989
rect 183437 212175 183747 220961
rect 183437 212147 183485 212175
rect 183513 212147 183547 212175
rect 183575 212147 183609 212175
rect 183637 212147 183671 212175
rect 183699 212147 183747 212175
rect 183437 212113 183747 212147
rect 183437 212085 183485 212113
rect 183513 212085 183547 212113
rect 183575 212085 183609 212113
rect 183637 212085 183671 212113
rect 183699 212085 183747 212113
rect 183437 212051 183747 212085
rect 183437 212023 183485 212051
rect 183513 212023 183547 212051
rect 183575 212023 183609 212051
rect 183637 212023 183671 212051
rect 183699 212023 183747 212051
rect 183437 211989 183747 212023
rect 183437 211961 183485 211989
rect 183513 211961 183547 211989
rect 183575 211961 183609 211989
rect 183637 211961 183671 211989
rect 183699 211961 183747 211989
rect 183437 203175 183747 211961
rect 183437 203147 183485 203175
rect 183513 203147 183547 203175
rect 183575 203147 183609 203175
rect 183637 203147 183671 203175
rect 183699 203147 183747 203175
rect 183437 203113 183747 203147
rect 183437 203085 183485 203113
rect 183513 203085 183547 203113
rect 183575 203085 183609 203113
rect 183637 203085 183671 203113
rect 183699 203085 183747 203113
rect 183437 203051 183747 203085
rect 183437 203023 183485 203051
rect 183513 203023 183547 203051
rect 183575 203023 183609 203051
rect 183637 203023 183671 203051
rect 183699 203023 183747 203051
rect 183437 202989 183747 203023
rect 183437 202961 183485 202989
rect 183513 202961 183547 202989
rect 183575 202961 183609 202989
rect 183637 202961 183671 202989
rect 183699 202961 183747 202989
rect 183437 194175 183747 202961
rect 183437 194147 183485 194175
rect 183513 194147 183547 194175
rect 183575 194147 183609 194175
rect 183637 194147 183671 194175
rect 183699 194147 183747 194175
rect 183437 194113 183747 194147
rect 183437 194085 183485 194113
rect 183513 194085 183547 194113
rect 183575 194085 183609 194113
rect 183637 194085 183671 194113
rect 183699 194085 183747 194113
rect 183437 194051 183747 194085
rect 183437 194023 183485 194051
rect 183513 194023 183547 194051
rect 183575 194023 183609 194051
rect 183637 194023 183671 194051
rect 183699 194023 183747 194051
rect 183437 193989 183747 194023
rect 183437 193961 183485 193989
rect 183513 193961 183547 193989
rect 183575 193961 183609 193989
rect 183637 193961 183671 193989
rect 183699 193961 183747 193989
rect 183437 185175 183747 193961
rect 183437 185147 183485 185175
rect 183513 185147 183547 185175
rect 183575 185147 183609 185175
rect 183637 185147 183671 185175
rect 183699 185147 183747 185175
rect 183437 185113 183747 185147
rect 183437 185085 183485 185113
rect 183513 185085 183547 185113
rect 183575 185085 183609 185113
rect 183637 185085 183671 185113
rect 183699 185085 183747 185113
rect 183437 185051 183747 185085
rect 183437 185023 183485 185051
rect 183513 185023 183547 185051
rect 183575 185023 183609 185051
rect 183637 185023 183671 185051
rect 183699 185023 183747 185051
rect 183437 184989 183747 185023
rect 183437 184961 183485 184989
rect 183513 184961 183547 184989
rect 183575 184961 183609 184989
rect 183637 184961 183671 184989
rect 183699 184961 183747 184989
rect 183437 176175 183747 184961
rect 183437 176147 183485 176175
rect 183513 176147 183547 176175
rect 183575 176147 183609 176175
rect 183637 176147 183671 176175
rect 183699 176147 183747 176175
rect 183437 176113 183747 176147
rect 183437 176085 183485 176113
rect 183513 176085 183547 176113
rect 183575 176085 183609 176113
rect 183637 176085 183671 176113
rect 183699 176085 183747 176113
rect 183437 176051 183747 176085
rect 183437 176023 183485 176051
rect 183513 176023 183547 176051
rect 183575 176023 183609 176051
rect 183637 176023 183671 176051
rect 183699 176023 183747 176051
rect 183437 175989 183747 176023
rect 183437 175961 183485 175989
rect 183513 175961 183547 175989
rect 183575 175961 183609 175989
rect 183637 175961 183671 175989
rect 183699 175961 183747 175989
rect 183437 167175 183747 175961
rect 183437 167147 183485 167175
rect 183513 167147 183547 167175
rect 183575 167147 183609 167175
rect 183637 167147 183671 167175
rect 183699 167147 183747 167175
rect 183437 167113 183747 167147
rect 183437 167085 183485 167113
rect 183513 167085 183547 167113
rect 183575 167085 183609 167113
rect 183637 167085 183671 167113
rect 183699 167085 183747 167113
rect 183437 167051 183747 167085
rect 183437 167023 183485 167051
rect 183513 167023 183547 167051
rect 183575 167023 183609 167051
rect 183637 167023 183671 167051
rect 183699 167023 183747 167051
rect 183437 166989 183747 167023
rect 183437 166961 183485 166989
rect 183513 166961 183547 166989
rect 183575 166961 183609 166989
rect 183637 166961 183671 166989
rect 183699 166961 183747 166989
rect 183437 158175 183747 166961
rect 183437 158147 183485 158175
rect 183513 158147 183547 158175
rect 183575 158147 183609 158175
rect 183637 158147 183671 158175
rect 183699 158147 183747 158175
rect 183437 158113 183747 158147
rect 183437 158085 183485 158113
rect 183513 158085 183547 158113
rect 183575 158085 183609 158113
rect 183637 158085 183671 158113
rect 183699 158085 183747 158113
rect 183437 158051 183747 158085
rect 183437 158023 183485 158051
rect 183513 158023 183547 158051
rect 183575 158023 183609 158051
rect 183637 158023 183671 158051
rect 183699 158023 183747 158051
rect 183437 157989 183747 158023
rect 183437 157961 183485 157989
rect 183513 157961 183547 157989
rect 183575 157961 183609 157989
rect 183637 157961 183671 157989
rect 183699 157961 183747 157989
rect 183437 149175 183747 157961
rect 183437 149147 183485 149175
rect 183513 149147 183547 149175
rect 183575 149147 183609 149175
rect 183637 149147 183671 149175
rect 183699 149147 183747 149175
rect 183437 149113 183747 149147
rect 183437 149085 183485 149113
rect 183513 149085 183547 149113
rect 183575 149085 183609 149113
rect 183637 149085 183671 149113
rect 183699 149085 183747 149113
rect 183437 149051 183747 149085
rect 183437 149023 183485 149051
rect 183513 149023 183547 149051
rect 183575 149023 183609 149051
rect 183637 149023 183671 149051
rect 183699 149023 183747 149051
rect 183437 148989 183747 149023
rect 183437 148961 183485 148989
rect 183513 148961 183547 148989
rect 183575 148961 183609 148989
rect 183637 148961 183671 148989
rect 183699 148961 183747 148989
rect 183437 140175 183747 148961
rect 183437 140147 183485 140175
rect 183513 140147 183547 140175
rect 183575 140147 183609 140175
rect 183637 140147 183671 140175
rect 183699 140147 183747 140175
rect 183437 140113 183747 140147
rect 183437 140085 183485 140113
rect 183513 140085 183547 140113
rect 183575 140085 183609 140113
rect 183637 140085 183671 140113
rect 183699 140085 183747 140113
rect 183437 140051 183747 140085
rect 183437 140023 183485 140051
rect 183513 140023 183547 140051
rect 183575 140023 183609 140051
rect 183637 140023 183671 140051
rect 183699 140023 183747 140051
rect 183437 139989 183747 140023
rect 183437 139961 183485 139989
rect 183513 139961 183547 139989
rect 183575 139961 183609 139989
rect 183637 139961 183671 139989
rect 183699 139961 183747 139989
rect 183437 131175 183747 139961
rect 183437 131147 183485 131175
rect 183513 131147 183547 131175
rect 183575 131147 183609 131175
rect 183637 131147 183671 131175
rect 183699 131147 183747 131175
rect 183437 131113 183747 131147
rect 183437 131085 183485 131113
rect 183513 131085 183547 131113
rect 183575 131085 183609 131113
rect 183637 131085 183671 131113
rect 183699 131085 183747 131113
rect 183437 131051 183747 131085
rect 183437 131023 183485 131051
rect 183513 131023 183547 131051
rect 183575 131023 183609 131051
rect 183637 131023 183671 131051
rect 183699 131023 183747 131051
rect 183437 130989 183747 131023
rect 183437 130961 183485 130989
rect 183513 130961 183547 130989
rect 183575 130961 183609 130989
rect 183637 130961 183671 130989
rect 183699 130961 183747 130989
rect 183437 122175 183747 130961
rect 183437 122147 183485 122175
rect 183513 122147 183547 122175
rect 183575 122147 183609 122175
rect 183637 122147 183671 122175
rect 183699 122147 183747 122175
rect 183437 122113 183747 122147
rect 183437 122085 183485 122113
rect 183513 122085 183547 122113
rect 183575 122085 183609 122113
rect 183637 122085 183671 122113
rect 183699 122085 183747 122113
rect 183437 122051 183747 122085
rect 183437 122023 183485 122051
rect 183513 122023 183547 122051
rect 183575 122023 183609 122051
rect 183637 122023 183671 122051
rect 183699 122023 183747 122051
rect 183437 121989 183747 122023
rect 183437 121961 183485 121989
rect 183513 121961 183547 121989
rect 183575 121961 183609 121989
rect 183637 121961 183671 121989
rect 183699 121961 183747 121989
rect 183437 113175 183747 121961
rect 183437 113147 183485 113175
rect 183513 113147 183547 113175
rect 183575 113147 183609 113175
rect 183637 113147 183671 113175
rect 183699 113147 183747 113175
rect 183437 113113 183747 113147
rect 183437 113085 183485 113113
rect 183513 113085 183547 113113
rect 183575 113085 183609 113113
rect 183637 113085 183671 113113
rect 183699 113085 183747 113113
rect 183437 113051 183747 113085
rect 183437 113023 183485 113051
rect 183513 113023 183547 113051
rect 183575 113023 183609 113051
rect 183637 113023 183671 113051
rect 183699 113023 183747 113051
rect 183437 112989 183747 113023
rect 183437 112961 183485 112989
rect 183513 112961 183547 112989
rect 183575 112961 183609 112989
rect 183637 112961 183671 112989
rect 183699 112961 183747 112989
rect 183437 104175 183747 112961
rect 183437 104147 183485 104175
rect 183513 104147 183547 104175
rect 183575 104147 183609 104175
rect 183637 104147 183671 104175
rect 183699 104147 183747 104175
rect 183437 104113 183747 104147
rect 183437 104085 183485 104113
rect 183513 104085 183547 104113
rect 183575 104085 183609 104113
rect 183637 104085 183671 104113
rect 183699 104085 183747 104113
rect 183437 104051 183747 104085
rect 183437 104023 183485 104051
rect 183513 104023 183547 104051
rect 183575 104023 183609 104051
rect 183637 104023 183671 104051
rect 183699 104023 183747 104051
rect 183437 103989 183747 104023
rect 183437 103961 183485 103989
rect 183513 103961 183547 103989
rect 183575 103961 183609 103989
rect 183637 103961 183671 103989
rect 183699 103961 183747 103989
rect 183437 95175 183747 103961
rect 183437 95147 183485 95175
rect 183513 95147 183547 95175
rect 183575 95147 183609 95175
rect 183637 95147 183671 95175
rect 183699 95147 183747 95175
rect 183437 95113 183747 95147
rect 183437 95085 183485 95113
rect 183513 95085 183547 95113
rect 183575 95085 183609 95113
rect 183637 95085 183671 95113
rect 183699 95085 183747 95113
rect 183437 95051 183747 95085
rect 183437 95023 183485 95051
rect 183513 95023 183547 95051
rect 183575 95023 183609 95051
rect 183637 95023 183671 95051
rect 183699 95023 183747 95051
rect 183437 94989 183747 95023
rect 183437 94961 183485 94989
rect 183513 94961 183547 94989
rect 183575 94961 183609 94989
rect 183637 94961 183671 94989
rect 183699 94961 183747 94989
rect 183437 86175 183747 94961
rect 183437 86147 183485 86175
rect 183513 86147 183547 86175
rect 183575 86147 183609 86175
rect 183637 86147 183671 86175
rect 183699 86147 183747 86175
rect 183437 86113 183747 86147
rect 183437 86085 183485 86113
rect 183513 86085 183547 86113
rect 183575 86085 183609 86113
rect 183637 86085 183671 86113
rect 183699 86085 183747 86113
rect 183437 86051 183747 86085
rect 183437 86023 183485 86051
rect 183513 86023 183547 86051
rect 183575 86023 183609 86051
rect 183637 86023 183671 86051
rect 183699 86023 183747 86051
rect 183437 85989 183747 86023
rect 183437 85961 183485 85989
rect 183513 85961 183547 85989
rect 183575 85961 183609 85989
rect 183637 85961 183671 85989
rect 183699 85961 183747 85989
rect 183437 77175 183747 85961
rect 183437 77147 183485 77175
rect 183513 77147 183547 77175
rect 183575 77147 183609 77175
rect 183637 77147 183671 77175
rect 183699 77147 183747 77175
rect 183437 77113 183747 77147
rect 183437 77085 183485 77113
rect 183513 77085 183547 77113
rect 183575 77085 183609 77113
rect 183637 77085 183671 77113
rect 183699 77085 183747 77113
rect 183437 77051 183747 77085
rect 183437 77023 183485 77051
rect 183513 77023 183547 77051
rect 183575 77023 183609 77051
rect 183637 77023 183671 77051
rect 183699 77023 183747 77051
rect 183437 76989 183747 77023
rect 183437 76961 183485 76989
rect 183513 76961 183547 76989
rect 183575 76961 183609 76989
rect 183637 76961 183671 76989
rect 183699 76961 183747 76989
rect 183437 68175 183747 76961
rect 183437 68147 183485 68175
rect 183513 68147 183547 68175
rect 183575 68147 183609 68175
rect 183637 68147 183671 68175
rect 183699 68147 183747 68175
rect 183437 68113 183747 68147
rect 183437 68085 183485 68113
rect 183513 68085 183547 68113
rect 183575 68085 183609 68113
rect 183637 68085 183671 68113
rect 183699 68085 183747 68113
rect 183437 68051 183747 68085
rect 183437 68023 183485 68051
rect 183513 68023 183547 68051
rect 183575 68023 183609 68051
rect 183637 68023 183671 68051
rect 183699 68023 183747 68051
rect 183437 67989 183747 68023
rect 183437 67961 183485 67989
rect 183513 67961 183547 67989
rect 183575 67961 183609 67989
rect 183637 67961 183671 67989
rect 183699 67961 183747 67989
rect 183437 59175 183747 67961
rect 183437 59147 183485 59175
rect 183513 59147 183547 59175
rect 183575 59147 183609 59175
rect 183637 59147 183671 59175
rect 183699 59147 183747 59175
rect 183437 59113 183747 59147
rect 183437 59085 183485 59113
rect 183513 59085 183547 59113
rect 183575 59085 183609 59113
rect 183637 59085 183671 59113
rect 183699 59085 183747 59113
rect 183437 59051 183747 59085
rect 183437 59023 183485 59051
rect 183513 59023 183547 59051
rect 183575 59023 183609 59051
rect 183637 59023 183671 59051
rect 183699 59023 183747 59051
rect 183437 58989 183747 59023
rect 183437 58961 183485 58989
rect 183513 58961 183547 58989
rect 183575 58961 183609 58989
rect 183637 58961 183671 58989
rect 183699 58961 183747 58989
rect 183437 50175 183747 58961
rect 183437 50147 183485 50175
rect 183513 50147 183547 50175
rect 183575 50147 183609 50175
rect 183637 50147 183671 50175
rect 183699 50147 183747 50175
rect 183437 50113 183747 50147
rect 183437 50085 183485 50113
rect 183513 50085 183547 50113
rect 183575 50085 183609 50113
rect 183637 50085 183671 50113
rect 183699 50085 183747 50113
rect 183437 50051 183747 50085
rect 183437 50023 183485 50051
rect 183513 50023 183547 50051
rect 183575 50023 183609 50051
rect 183637 50023 183671 50051
rect 183699 50023 183747 50051
rect 183437 49989 183747 50023
rect 183437 49961 183485 49989
rect 183513 49961 183547 49989
rect 183575 49961 183609 49989
rect 183637 49961 183671 49989
rect 183699 49961 183747 49989
rect 183437 41175 183747 49961
rect 183437 41147 183485 41175
rect 183513 41147 183547 41175
rect 183575 41147 183609 41175
rect 183637 41147 183671 41175
rect 183699 41147 183747 41175
rect 183437 41113 183747 41147
rect 183437 41085 183485 41113
rect 183513 41085 183547 41113
rect 183575 41085 183609 41113
rect 183637 41085 183671 41113
rect 183699 41085 183747 41113
rect 183437 41051 183747 41085
rect 183437 41023 183485 41051
rect 183513 41023 183547 41051
rect 183575 41023 183609 41051
rect 183637 41023 183671 41051
rect 183699 41023 183747 41051
rect 183437 40989 183747 41023
rect 183437 40961 183485 40989
rect 183513 40961 183547 40989
rect 183575 40961 183609 40989
rect 183637 40961 183671 40989
rect 183699 40961 183747 40989
rect 183437 32175 183747 40961
rect 183437 32147 183485 32175
rect 183513 32147 183547 32175
rect 183575 32147 183609 32175
rect 183637 32147 183671 32175
rect 183699 32147 183747 32175
rect 183437 32113 183747 32147
rect 183437 32085 183485 32113
rect 183513 32085 183547 32113
rect 183575 32085 183609 32113
rect 183637 32085 183671 32113
rect 183699 32085 183747 32113
rect 183437 32051 183747 32085
rect 183437 32023 183485 32051
rect 183513 32023 183547 32051
rect 183575 32023 183609 32051
rect 183637 32023 183671 32051
rect 183699 32023 183747 32051
rect 183437 31989 183747 32023
rect 183437 31961 183485 31989
rect 183513 31961 183547 31989
rect 183575 31961 183609 31989
rect 183637 31961 183671 31989
rect 183699 31961 183747 31989
rect 183437 23175 183747 31961
rect 183437 23147 183485 23175
rect 183513 23147 183547 23175
rect 183575 23147 183609 23175
rect 183637 23147 183671 23175
rect 183699 23147 183747 23175
rect 183437 23113 183747 23147
rect 183437 23085 183485 23113
rect 183513 23085 183547 23113
rect 183575 23085 183609 23113
rect 183637 23085 183671 23113
rect 183699 23085 183747 23113
rect 183437 23051 183747 23085
rect 183437 23023 183485 23051
rect 183513 23023 183547 23051
rect 183575 23023 183609 23051
rect 183637 23023 183671 23051
rect 183699 23023 183747 23051
rect 183437 22989 183747 23023
rect 183437 22961 183485 22989
rect 183513 22961 183547 22989
rect 183575 22961 183609 22989
rect 183637 22961 183671 22989
rect 183699 22961 183747 22989
rect 183437 14175 183747 22961
rect 183437 14147 183485 14175
rect 183513 14147 183547 14175
rect 183575 14147 183609 14175
rect 183637 14147 183671 14175
rect 183699 14147 183747 14175
rect 183437 14113 183747 14147
rect 183437 14085 183485 14113
rect 183513 14085 183547 14113
rect 183575 14085 183609 14113
rect 183637 14085 183671 14113
rect 183699 14085 183747 14113
rect 183437 14051 183747 14085
rect 183437 14023 183485 14051
rect 183513 14023 183547 14051
rect 183575 14023 183609 14051
rect 183637 14023 183671 14051
rect 183699 14023 183747 14051
rect 183437 13989 183747 14023
rect 183437 13961 183485 13989
rect 183513 13961 183547 13989
rect 183575 13961 183609 13989
rect 183637 13961 183671 13989
rect 183699 13961 183747 13989
rect 183437 5175 183747 13961
rect 183437 5147 183485 5175
rect 183513 5147 183547 5175
rect 183575 5147 183609 5175
rect 183637 5147 183671 5175
rect 183699 5147 183747 5175
rect 183437 5113 183747 5147
rect 183437 5085 183485 5113
rect 183513 5085 183547 5113
rect 183575 5085 183609 5113
rect 183637 5085 183671 5113
rect 183699 5085 183747 5113
rect 183437 5051 183747 5085
rect 183437 5023 183485 5051
rect 183513 5023 183547 5051
rect 183575 5023 183609 5051
rect 183637 5023 183671 5051
rect 183699 5023 183747 5051
rect 183437 4989 183747 5023
rect 183437 4961 183485 4989
rect 183513 4961 183547 4989
rect 183575 4961 183609 4989
rect 183637 4961 183671 4989
rect 183699 4961 183747 4989
rect 183437 -560 183747 4961
rect 183437 -588 183485 -560
rect 183513 -588 183547 -560
rect 183575 -588 183609 -560
rect 183637 -588 183671 -560
rect 183699 -588 183747 -560
rect 183437 -622 183747 -588
rect 183437 -650 183485 -622
rect 183513 -650 183547 -622
rect 183575 -650 183609 -622
rect 183637 -650 183671 -622
rect 183699 -650 183747 -622
rect 183437 -684 183747 -650
rect 183437 -712 183485 -684
rect 183513 -712 183547 -684
rect 183575 -712 183609 -684
rect 183637 -712 183671 -684
rect 183699 -712 183747 -684
rect 183437 -746 183747 -712
rect 183437 -774 183485 -746
rect 183513 -774 183547 -746
rect 183575 -774 183609 -746
rect 183637 -774 183671 -746
rect 183699 -774 183747 -746
rect 183437 -822 183747 -774
rect 190577 298606 190887 299134
rect 190577 298578 190625 298606
rect 190653 298578 190687 298606
rect 190715 298578 190749 298606
rect 190777 298578 190811 298606
rect 190839 298578 190887 298606
rect 190577 298544 190887 298578
rect 190577 298516 190625 298544
rect 190653 298516 190687 298544
rect 190715 298516 190749 298544
rect 190777 298516 190811 298544
rect 190839 298516 190887 298544
rect 190577 298482 190887 298516
rect 190577 298454 190625 298482
rect 190653 298454 190687 298482
rect 190715 298454 190749 298482
rect 190777 298454 190811 298482
rect 190839 298454 190887 298482
rect 190577 298420 190887 298454
rect 190577 298392 190625 298420
rect 190653 298392 190687 298420
rect 190715 298392 190749 298420
rect 190777 298392 190811 298420
rect 190839 298392 190887 298420
rect 190577 290175 190887 298392
rect 190577 290147 190625 290175
rect 190653 290147 190687 290175
rect 190715 290147 190749 290175
rect 190777 290147 190811 290175
rect 190839 290147 190887 290175
rect 190577 290113 190887 290147
rect 190577 290085 190625 290113
rect 190653 290085 190687 290113
rect 190715 290085 190749 290113
rect 190777 290085 190811 290113
rect 190839 290085 190887 290113
rect 190577 290051 190887 290085
rect 190577 290023 190625 290051
rect 190653 290023 190687 290051
rect 190715 290023 190749 290051
rect 190777 290023 190811 290051
rect 190839 290023 190887 290051
rect 190577 289989 190887 290023
rect 190577 289961 190625 289989
rect 190653 289961 190687 289989
rect 190715 289961 190749 289989
rect 190777 289961 190811 289989
rect 190839 289961 190887 289989
rect 190577 281175 190887 289961
rect 190577 281147 190625 281175
rect 190653 281147 190687 281175
rect 190715 281147 190749 281175
rect 190777 281147 190811 281175
rect 190839 281147 190887 281175
rect 190577 281113 190887 281147
rect 190577 281085 190625 281113
rect 190653 281085 190687 281113
rect 190715 281085 190749 281113
rect 190777 281085 190811 281113
rect 190839 281085 190887 281113
rect 190577 281051 190887 281085
rect 190577 281023 190625 281051
rect 190653 281023 190687 281051
rect 190715 281023 190749 281051
rect 190777 281023 190811 281051
rect 190839 281023 190887 281051
rect 190577 280989 190887 281023
rect 190577 280961 190625 280989
rect 190653 280961 190687 280989
rect 190715 280961 190749 280989
rect 190777 280961 190811 280989
rect 190839 280961 190887 280989
rect 190577 272175 190887 280961
rect 190577 272147 190625 272175
rect 190653 272147 190687 272175
rect 190715 272147 190749 272175
rect 190777 272147 190811 272175
rect 190839 272147 190887 272175
rect 190577 272113 190887 272147
rect 190577 272085 190625 272113
rect 190653 272085 190687 272113
rect 190715 272085 190749 272113
rect 190777 272085 190811 272113
rect 190839 272085 190887 272113
rect 190577 272051 190887 272085
rect 190577 272023 190625 272051
rect 190653 272023 190687 272051
rect 190715 272023 190749 272051
rect 190777 272023 190811 272051
rect 190839 272023 190887 272051
rect 190577 271989 190887 272023
rect 190577 271961 190625 271989
rect 190653 271961 190687 271989
rect 190715 271961 190749 271989
rect 190777 271961 190811 271989
rect 190839 271961 190887 271989
rect 190577 263175 190887 271961
rect 190577 263147 190625 263175
rect 190653 263147 190687 263175
rect 190715 263147 190749 263175
rect 190777 263147 190811 263175
rect 190839 263147 190887 263175
rect 190577 263113 190887 263147
rect 190577 263085 190625 263113
rect 190653 263085 190687 263113
rect 190715 263085 190749 263113
rect 190777 263085 190811 263113
rect 190839 263085 190887 263113
rect 190577 263051 190887 263085
rect 190577 263023 190625 263051
rect 190653 263023 190687 263051
rect 190715 263023 190749 263051
rect 190777 263023 190811 263051
rect 190839 263023 190887 263051
rect 190577 262989 190887 263023
rect 190577 262961 190625 262989
rect 190653 262961 190687 262989
rect 190715 262961 190749 262989
rect 190777 262961 190811 262989
rect 190839 262961 190887 262989
rect 190577 254175 190887 262961
rect 190577 254147 190625 254175
rect 190653 254147 190687 254175
rect 190715 254147 190749 254175
rect 190777 254147 190811 254175
rect 190839 254147 190887 254175
rect 190577 254113 190887 254147
rect 190577 254085 190625 254113
rect 190653 254085 190687 254113
rect 190715 254085 190749 254113
rect 190777 254085 190811 254113
rect 190839 254085 190887 254113
rect 190577 254051 190887 254085
rect 190577 254023 190625 254051
rect 190653 254023 190687 254051
rect 190715 254023 190749 254051
rect 190777 254023 190811 254051
rect 190839 254023 190887 254051
rect 190577 253989 190887 254023
rect 190577 253961 190625 253989
rect 190653 253961 190687 253989
rect 190715 253961 190749 253989
rect 190777 253961 190811 253989
rect 190839 253961 190887 253989
rect 190577 245175 190887 253961
rect 190577 245147 190625 245175
rect 190653 245147 190687 245175
rect 190715 245147 190749 245175
rect 190777 245147 190811 245175
rect 190839 245147 190887 245175
rect 190577 245113 190887 245147
rect 190577 245085 190625 245113
rect 190653 245085 190687 245113
rect 190715 245085 190749 245113
rect 190777 245085 190811 245113
rect 190839 245085 190887 245113
rect 190577 245051 190887 245085
rect 190577 245023 190625 245051
rect 190653 245023 190687 245051
rect 190715 245023 190749 245051
rect 190777 245023 190811 245051
rect 190839 245023 190887 245051
rect 190577 244989 190887 245023
rect 190577 244961 190625 244989
rect 190653 244961 190687 244989
rect 190715 244961 190749 244989
rect 190777 244961 190811 244989
rect 190839 244961 190887 244989
rect 190577 236175 190887 244961
rect 190577 236147 190625 236175
rect 190653 236147 190687 236175
rect 190715 236147 190749 236175
rect 190777 236147 190811 236175
rect 190839 236147 190887 236175
rect 190577 236113 190887 236147
rect 190577 236085 190625 236113
rect 190653 236085 190687 236113
rect 190715 236085 190749 236113
rect 190777 236085 190811 236113
rect 190839 236085 190887 236113
rect 190577 236051 190887 236085
rect 190577 236023 190625 236051
rect 190653 236023 190687 236051
rect 190715 236023 190749 236051
rect 190777 236023 190811 236051
rect 190839 236023 190887 236051
rect 190577 235989 190887 236023
rect 190577 235961 190625 235989
rect 190653 235961 190687 235989
rect 190715 235961 190749 235989
rect 190777 235961 190811 235989
rect 190839 235961 190887 235989
rect 190577 227175 190887 235961
rect 190577 227147 190625 227175
rect 190653 227147 190687 227175
rect 190715 227147 190749 227175
rect 190777 227147 190811 227175
rect 190839 227147 190887 227175
rect 190577 227113 190887 227147
rect 190577 227085 190625 227113
rect 190653 227085 190687 227113
rect 190715 227085 190749 227113
rect 190777 227085 190811 227113
rect 190839 227085 190887 227113
rect 190577 227051 190887 227085
rect 190577 227023 190625 227051
rect 190653 227023 190687 227051
rect 190715 227023 190749 227051
rect 190777 227023 190811 227051
rect 190839 227023 190887 227051
rect 190577 226989 190887 227023
rect 190577 226961 190625 226989
rect 190653 226961 190687 226989
rect 190715 226961 190749 226989
rect 190777 226961 190811 226989
rect 190839 226961 190887 226989
rect 190577 218175 190887 226961
rect 190577 218147 190625 218175
rect 190653 218147 190687 218175
rect 190715 218147 190749 218175
rect 190777 218147 190811 218175
rect 190839 218147 190887 218175
rect 190577 218113 190887 218147
rect 190577 218085 190625 218113
rect 190653 218085 190687 218113
rect 190715 218085 190749 218113
rect 190777 218085 190811 218113
rect 190839 218085 190887 218113
rect 190577 218051 190887 218085
rect 190577 218023 190625 218051
rect 190653 218023 190687 218051
rect 190715 218023 190749 218051
rect 190777 218023 190811 218051
rect 190839 218023 190887 218051
rect 190577 217989 190887 218023
rect 190577 217961 190625 217989
rect 190653 217961 190687 217989
rect 190715 217961 190749 217989
rect 190777 217961 190811 217989
rect 190839 217961 190887 217989
rect 190577 209175 190887 217961
rect 190577 209147 190625 209175
rect 190653 209147 190687 209175
rect 190715 209147 190749 209175
rect 190777 209147 190811 209175
rect 190839 209147 190887 209175
rect 190577 209113 190887 209147
rect 190577 209085 190625 209113
rect 190653 209085 190687 209113
rect 190715 209085 190749 209113
rect 190777 209085 190811 209113
rect 190839 209085 190887 209113
rect 190577 209051 190887 209085
rect 190577 209023 190625 209051
rect 190653 209023 190687 209051
rect 190715 209023 190749 209051
rect 190777 209023 190811 209051
rect 190839 209023 190887 209051
rect 190577 208989 190887 209023
rect 190577 208961 190625 208989
rect 190653 208961 190687 208989
rect 190715 208961 190749 208989
rect 190777 208961 190811 208989
rect 190839 208961 190887 208989
rect 190577 200175 190887 208961
rect 190577 200147 190625 200175
rect 190653 200147 190687 200175
rect 190715 200147 190749 200175
rect 190777 200147 190811 200175
rect 190839 200147 190887 200175
rect 190577 200113 190887 200147
rect 190577 200085 190625 200113
rect 190653 200085 190687 200113
rect 190715 200085 190749 200113
rect 190777 200085 190811 200113
rect 190839 200085 190887 200113
rect 190577 200051 190887 200085
rect 190577 200023 190625 200051
rect 190653 200023 190687 200051
rect 190715 200023 190749 200051
rect 190777 200023 190811 200051
rect 190839 200023 190887 200051
rect 190577 199989 190887 200023
rect 190577 199961 190625 199989
rect 190653 199961 190687 199989
rect 190715 199961 190749 199989
rect 190777 199961 190811 199989
rect 190839 199961 190887 199989
rect 190577 191175 190887 199961
rect 190577 191147 190625 191175
rect 190653 191147 190687 191175
rect 190715 191147 190749 191175
rect 190777 191147 190811 191175
rect 190839 191147 190887 191175
rect 190577 191113 190887 191147
rect 190577 191085 190625 191113
rect 190653 191085 190687 191113
rect 190715 191085 190749 191113
rect 190777 191085 190811 191113
rect 190839 191085 190887 191113
rect 190577 191051 190887 191085
rect 190577 191023 190625 191051
rect 190653 191023 190687 191051
rect 190715 191023 190749 191051
rect 190777 191023 190811 191051
rect 190839 191023 190887 191051
rect 190577 190989 190887 191023
rect 190577 190961 190625 190989
rect 190653 190961 190687 190989
rect 190715 190961 190749 190989
rect 190777 190961 190811 190989
rect 190839 190961 190887 190989
rect 190577 182175 190887 190961
rect 190577 182147 190625 182175
rect 190653 182147 190687 182175
rect 190715 182147 190749 182175
rect 190777 182147 190811 182175
rect 190839 182147 190887 182175
rect 190577 182113 190887 182147
rect 190577 182085 190625 182113
rect 190653 182085 190687 182113
rect 190715 182085 190749 182113
rect 190777 182085 190811 182113
rect 190839 182085 190887 182113
rect 190577 182051 190887 182085
rect 190577 182023 190625 182051
rect 190653 182023 190687 182051
rect 190715 182023 190749 182051
rect 190777 182023 190811 182051
rect 190839 182023 190887 182051
rect 190577 181989 190887 182023
rect 190577 181961 190625 181989
rect 190653 181961 190687 181989
rect 190715 181961 190749 181989
rect 190777 181961 190811 181989
rect 190839 181961 190887 181989
rect 190577 173175 190887 181961
rect 190577 173147 190625 173175
rect 190653 173147 190687 173175
rect 190715 173147 190749 173175
rect 190777 173147 190811 173175
rect 190839 173147 190887 173175
rect 190577 173113 190887 173147
rect 190577 173085 190625 173113
rect 190653 173085 190687 173113
rect 190715 173085 190749 173113
rect 190777 173085 190811 173113
rect 190839 173085 190887 173113
rect 190577 173051 190887 173085
rect 190577 173023 190625 173051
rect 190653 173023 190687 173051
rect 190715 173023 190749 173051
rect 190777 173023 190811 173051
rect 190839 173023 190887 173051
rect 190577 172989 190887 173023
rect 190577 172961 190625 172989
rect 190653 172961 190687 172989
rect 190715 172961 190749 172989
rect 190777 172961 190811 172989
rect 190839 172961 190887 172989
rect 190577 164175 190887 172961
rect 190577 164147 190625 164175
rect 190653 164147 190687 164175
rect 190715 164147 190749 164175
rect 190777 164147 190811 164175
rect 190839 164147 190887 164175
rect 190577 164113 190887 164147
rect 190577 164085 190625 164113
rect 190653 164085 190687 164113
rect 190715 164085 190749 164113
rect 190777 164085 190811 164113
rect 190839 164085 190887 164113
rect 190577 164051 190887 164085
rect 190577 164023 190625 164051
rect 190653 164023 190687 164051
rect 190715 164023 190749 164051
rect 190777 164023 190811 164051
rect 190839 164023 190887 164051
rect 190577 163989 190887 164023
rect 190577 163961 190625 163989
rect 190653 163961 190687 163989
rect 190715 163961 190749 163989
rect 190777 163961 190811 163989
rect 190839 163961 190887 163989
rect 190577 155175 190887 163961
rect 190577 155147 190625 155175
rect 190653 155147 190687 155175
rect 190715 155147 190749 155175
rect 190777 155147 190811 155175
rect 190839 155147 190887 155175
rect 190577 155113 190887 155147
rect 190577 155085 190625 155113
rect 190653 155085 190687 155113
rect 190715 155085 190749 155113
rect 190777 155085 190811 155113
rect 190839 155085 190887 155113
rect 190577 155051 190887 155085
rect 190577 155023 190625 155051
rect 190653 155023 190687 155051
rect 190715 155023 190749 155051
rect 190777 155023 190811 155051
rect 190839 155023 190887 155051
rect 190577 154989 190887 155023
rect 190577 154961 190625 154989
rect 190653 154961 190687 154989
rect 190715 154961 190749 154989
rect 190777 154961 190811 154989
rect 190839 154961 190887 154989
rect 190577 146175 190887 154961
rect 190577 146147 190625 146175
rect 190653 146147 190687 146175
rect 190715 146147 190749 146175
rect 190777 146147 190811 146175
rect 190839 146147 190887 146175
rect 190577 146113 190887 146147
rect 190577 146085 190625 146113
rect 190653 146085 190687 146113
rect 190715 146085 190749 146113
rect 190777 146085 190811 146113
rect 190839 146085 190887 146113
rect 190577 146051 190887 146085
rect 190577 146023 190625 146051
rect 190653 146023 190687 146051
rect 190715 146023 190749 146051
rect 190777 146023 190811 146051
rect 190839 146023 190887 146051
rect 190577 145989 190887 146023
rect 190577 145961 190625 145989
rect 190653 145961 190687 145989
rect 190715 145961 190749 145989
rect 190777 145961 190811 145989
rect 190839 145961 190887 145989
rect 190577 137175 190887 145961
rect 190577 137147 190625 137175
rect 190653 137147 190687 137175
rect 190715 137147 190749 137175
rect 190777 137147 190811 137175
rect 190839 137147 190887 137175
rect 190577 137113 190887 137147
rect 190577 137085 190625 137113
rect 190653 137085 190687 137113
rect 190715 137085 190749 137113
rect 190777 137085 190811 137113
rect 190839 137085 190887 137113
rect 190577 137051 190887 137085
rect 190577 137023 190625 137051
rect 190653 137023 190687 137051
rect 190715 137023 190749 137051
rect 190777 137023 190811 137051
rect 190839 137023 190887 137051
rect 190577 136989 190887 137023
rect 190577 136961 190625 136989
rect 190653 136961 190687 136989
rect 190715 136961 190749 136989
rect 190777 136961 190811 136989
rect 190839 136961 190887 136989
rect 190577 128175 190887 136961
rect 190577 128147 190625 128175
rect 190653 128147 190687 128175
rect 190715 128147 190749 128175
rect 190777 128147 190811 128175
rect 190839 128147 190887 128175
rect 190577 128113 190887 128147
rect 190577 128085 190625 128113
rect 190653 128085 190687 128113
rect 190715 128085 190749 128113
rect 190777 128085 190811 128113
rect 190839 128085 190887 128113
rect 190577 128051 190887 128085
rect 190577 128023 190625 128051
rect 190653 128023 190687 128051
rect 190715 128023 190749 128051
rect 190777 128023 190811 128051
rect 190839 128023 190887 128051
rect 190577 127989 190887 128023
rect 190577 127961 190625 127989
rect 190653 127961 190687 127989
rect 190715 127961 190749 127989
rect 190777 127961 190811 127989
rect 190839 127961 190887 127989
rect 190577 119175 190887 127961
rect 190577 119147 190625 119175
rect 190653 119147 190687 119175
rect 190715 119147 190749 119175
rect 190777 119147 190811 119175
rect 190839 119147 190887 119175
rect 190577 119113 190887 119147
rect 190577 119085 190625 119113
rect 190653 119085 190687 119113
rect 190715 119085 190749 119113
rect 190777 119085 190811 119113
rect 190839 119085 190887 119113
rect 190577 119051 190887 119085
rect 190577 119023 190625 119051
rect 190653 119023 190687 119051
rect 190715 119023 190749 119051
rect 190777 119023 190811 119051
rect 190839 119023 190887 119051
rect 190577 118989 190887 119023
rect 190577 118961 190625 118989
rect 190653 118961 190687 118989
rect 190715 118961 190749 118989
rect 190777 118961 190811 118989
rect 190839 118961 190887 118989
rect 190577 110175 190887 118961
rect 190577 110147 190625 110175
rect 190653 110147 190687 110175
rect 190715 110147 190749 110175
rect 190777 110147 190811 110175
rect 190839 110147 190887 110175
rect 190577 110113 190887 110147
rect 190577 110085 190625 110113
rect 190653 110085 190687 110113
rect 190715 110085 190749 110113
rect 190777 110085 190811 110113
rect 190839 110085 190887 110113
rect 190577 110051 190887 110085
rect 190577 110023 190625 110051
rect 190653 110023 190687 110051
rect 190715 110023 190749 110051
rect 190777 110023 190811 110051
rect 190839 110023 190887 110051
rect 190577 109989 190887 110023
rect 190577 109961 190625 109989
rect 190653 109961 190687 109989
rect 190715 109961 190749 109989
rect 190777 109961 190811 109989
rect 190839 109961 190887 109989
rect 190577 101175 190887 109961
rect 190577 101147 190625 101175
rect 190653 101147 190687 101175
rect 190715 101147 190749 101175
rect 190777 101147 190811 101175
rect 190839 101147 190887 101175
rect 190577 101113 190887 101147
rect 190577 101085 190625 101113
rect 190653 101085 190687 101113
rect 190715 101085 190749 101113
rect 190777 101085 190811 101113
rect 190839 101085 190887 101113
rect 190577 101051 190887 101085
rect 190577 101023 190625 101051
rect 190653 101023 190687 101051
rect 190715 101023 190749 101051
rect 190777 101023 190811 101051
rect 190839 101023 190887 101051
rect 190577 100989 190887 101023
rect 190577 100961 190625 100989
rect 190653 100961 190687 100989
rect 190715 100961 190749 100989
rect 190777 100961 190811 100989
rect 190839 100961 190887 100989
rect 190577 92175 190887 100961
rect 190577 92147 190625 92175
rect 190653 92147 190687 92175
rect 190715 92147 190749 92175
rect 190777 92147 190811 92175
rect 190839 92147 190887 92175
rect 190577 92113 190887 92147
rect 190577 92085 190625 92113
rect 190653 92085 190687 92113
rect 190715 92085 190749 92113
rect 190777 92085 190811 92113
rect 190839 92085 190887 92113
rect 190577 92051 190887 92085
rect 190577 92023 190625 92051
rect 190653 92023 190687 92051
rect 190715 92023 190749 92051
rect 190777 92023 190811 92051
rect 190839 92023 190887 92051
rect 190577 91989 190887 92023
rect 190577 91961 190625 91989
rect 190653 91961 190687 91989
rect 190715 91961 190749 91989
rect 190777 91961 190811 91989
rect 190839 91961 190887 91989
rect 190577 83175 190887 91961
rect 190577 83147 190625 83175
rect 190653 83147 190687 83175
rect 190715 83147 190749 83175
rect 190777 83147 190811 83175
rect 190839 83147 190887 83175
rect 190577 83113 190887 83147
rect 190577 83085 190625 83113
rect 190653 83085 190687 83113
rect 190715 83085 190749 83113
rect 190777 83085 190811 83113
rect 190839 83085 190887 83113
rect 190577 83051 190887 83085
rect 190577 83023 190625 83051
rect 190653 83023 190687 83051
rect 190715 83023 190749 83051
rect 190777 83023 190811 83051
rect 190839 83023 190887 83051
rect 190577 82989 190887 83023
rect 190577 82961 190625 82989
rect 190653 82961 190687 82989
rect 190715 82961 190749 82989
rect 190777 82961 190811 82989
rect 190839 82961 190887 82989
rect 190577 74175 190887 82961
rect 190577 74147 190625 74175
rect 190653 74147 190687 74175
rect 190715 74147 190749 74175
rect 190777 74147 190811 74175
rect 190839 74147 190887 74175
rect 190577 74113 190887 74147
rect 190577 74085 190625 74113
rect 190653 74085 190687 74113
rect 190715 74085 190749 74113
rect 190777 74085 190811 74113
rect 190839 74085 190887 74113
rect 190577 74051 190887 74085
rect 190577 74023 190625 74051
rect 190653 74023 190687 74051
rect 190715 74023 190749 74051
rect 190777 74023 190811 74051
rect 190839 74023 190887 74051
rect 190577 73989 190887 74023
rect 190577 73961 190625 73989
rect 190653 73961 190687 73989
rect 190715 73961 190749 73989
rect 190777 73961 190811 73989
rect 190839 73961 190887 73989
rect 190577 65175 190887 73961
rect 190577 65147 190625 65175
rect 190653 65147 190687 65175
rect 190715 65147 190749 65175
rect 190777 65147 190811 65175
rect 190839 65147 190887 65175
rect 190577 65113 190887 65147
rect 190577 65085 190625 65113
rect 190653 65085 190687 65113
rect 190715 65085 190749 65113
rect 190777 65085 190811 65113
rect 190839 65085 190887 65113
rect 190577 65051 190887 65085
rect 190577 65023 190625 65051
rect 190653 65023 190687 65051
rect 190715 65023 190749 65051
rect 190777 65023 190811 65051
rect 190839 65023 190887 65051
rect 190577 64989 190887 65023
rect 190577 64961 190625 64989
rect 190653 64961 190687 64989
rect 190715 64961 190749 64989
rect 190777 64961 190811 64989
rect 190839 64961 190887 64989
rect 190577 56175 190887 64961
rect 190577 56147 190625 56175
rect 190653 56147 190687 56175
rect 190715 56147 190749 56175
rect 190777 56147 190811 56175
rect 190839 56147 190887 56175
rect 190577 56113 190887 56147
rect 190577 56085 190625 56113
rect 190653 56085 190687 56113
rect 190715 56085 190749 56113
rect 190777 56085 190811 56113
rect 190839 56085 190887 56113
rect 190577 56051 190887 56085
rect 190577 56023 190625 56051
rect 190653 56023 190687 56051
rect 190715 56023 190749 56051
rect 190777 56023 190811 56051
rect 190839 56023 190887 56051
rect 190577 55989 190887 56023
rect 190577 55961 190625 55989
rect 190653 55961 190687 55989
rect 190715 55961 190749 55989
rect 190777 55961 190811 55989
rect 190839 55961 190887 55989
rect 190577 47175 190887 55961
rect 190577 47147 190625 47175
rect 190653 47147 190687 47175
rect 190715 47147 190749 47175
rect 190777 47147 190811 47175
rect 190839 47147 190887 47175
rect 190577 47113 190887 47147
rect 190577 47085 190625 47113
rect 190653 47085 190687 47113
rect 190715 47085 190749 47113
rect 190777 47085 190811 47113
rect 190839 47085 190887 47113
rect 190577 47051 190887 47085
rect 190577 47023 190625 47051
rect 190653 47023 190687 47051
rect 190715 47023 190749 47051
rect 190777 47023 190811 47051
rect 190839 47023 190887 47051
rect 190577 46989 190887 47023
rect 190577 46961 190625 46989
rect 190653 46961 190687 46989
rect 190715 46961 190749 46989
rect 190777 46961 190811 46989
rect 190839 46961 190887 46989
rect 190577 38175 190887 46961
rect 190577 38147 190625 38175
rect 190653 38147 190687 38175
rect 190715 38147 190749 38175
rect 190777 38147 190811 38175
rect 190839 38147 190887 38175
rect 190577 38113 190887 38147
rect 190577 38085 190625 38113
rect 190653 38085 190687 38113
rect 190715 38085 190749 38113
rect 190777 38085 190811 38113
rect 190839 38085 190887 38113
rect 190577 38051 190887 38085
rect 190577 38023 190625 38051
rect 190653 38023 190687 38051
rect 190715 38023 190749 38051
rect 190777 38023 190811 38051
rect 190839 38023 190887 38051
rect 190577 37989 190887 38023
rect 190577 37961 190625 37989
rect 190653 37961 190687 37989
rect 190715 37961 190749 37989
rect 190777 37961 190811 37989
rect 190839 37961 190887 37989
rect 190577 29175 190887 37961
rect 190577 29147 190625 29175
rect 190653 29147 190687 29175
rect 190715 29147 190749 29175
rect 190777 29147 190811 29175
rect 190839 29147 190887 29175
rect 190577 29113 190887 29147
rect 190577 29085 190625 29113
rect 190653 29085 190687 29113
rect 190715 29085 190749 29113
rect 190777 29085 190811 29113
rect 190839 29085 190887 29113
rect 190577 29051 190887 29085
rect 190577 29023 190625 29051
rect 190653 29023 190687 29051
rect 190715 29023 190749 29051
rect 190777 29023 190811 29051
rect 190839 29023 190887 29051
rect 190577 28989 190887 29023
rect 190577 28961 190625 28989
rect 190653 28961 190687 28989
rect 190715 28961 190749 28989
rect 190777 28961 190811 28989
rect 190839 28961 190887 28989
rect 190577 20175 190887 28961
rect 190577 20147 190625 20175
rect 190653 20147 190687 20175
rect 190715 20147 190749 20175
rect 190777 20147 190811 20175
rect 190839 20147 190887 20175
rect 190577 20113 190887 20147
rect 190577 20085 190625 20113
rect 190653 20085 190687 20113
rect 190715 20085 190749 20113
rect 190777 20085 190811 20113
rect 190839 20085 190887 20113
rect 190577 20051 190887 20085
rect 190577 20023 190625 20051
rect 190653 20023 190687 20051
rect 190715 20023 190749 20051
rect 190777 20023 190811 20051
rect 190839 20023 190887 20051
rect 190577 19989 190887 20023
rect 190577 19961 190625 19989
rect 190653 19961 190687 19989
rect 190715 19961 190749 19989
rect 190777 19961 190811 19989
rect 190839 19961 190887 19989
rect 190577 11175 190887 19961
rect 190577 11147 190625 11175
rect 190653 11147 190687 11175
rect 190715 11147 190749 11175
rect 190777 11147 190811 11175
rect 190839 11147 190887 11175
rect 190577 11113 190887 11147
rect 190577 11085 190625 11113
rect 190653 11085 190687 11113
rect 190715 11085 190749 11113
rect 190777 11085 190811 11113
rect 190839 11085 190887 11113
rect 190577 11051 190887 11085
rect 190577 11023 190625 11051
rect 190653 11023 190687 11051
rect 190715 11023 190749 11051
rect 190777 11023 190811 11051
rect 190839 11023 190887 11051
rect 190577 10989 190887 11023
rect 190577 10961 190625 10989
rect 190653 10961 190687 10989
rect 190715 10961 190749 10989
rect 190777 10961 190811 10989
rect 190839 10961 190887 10989
rect 190577 2175 190887 10961
rect 190577 2147 190625 2175
rect 190653 2147 190687 2175
rect 190715 2147 190749 2175
rect 190777 2147 190811 2175
rect 190839 2147 190887 2175
rect 190577 2113 190887 2147
rect 190577 2085 190625 2113
rect 190653 2085 190687 2113
rect 190715 2085 190749 2113
rect 190777 2085 190811 2113
rect 190839 2085 190887 2113
rect 190577 2051 190887 2085
rect 190577 2023 190625 2051
rect 190653 2023 190687 2051
rect 190715 2023 190749 2051
rect 190777 2023 190811 2051
rect 190839 2023 190887 2051
rect 190577 1989 190887 2023
rect 190577 1961 190625 1989
rect 190653 1961 190687 1989
rect 190715 1961 190749 1989
rect 190777 1961 190811 1989
rect 190839 1961 190887 1989
rect 190577 -80 190887 1961
rect 190577 -108 190625 -80
rect 190653 -108 190687 -80
rect 190715 -108 190749 -80
rect 190777 -108 190811 -80
rect 190839 -108 190887 -80
rect 190577 -142 190887 -108
rect 190577 -170 190625 -142
rect 190653 -170 190687 -142
rect 190715 -170 190749 -142
rect 190777 -170 190811 -142
rect 190839 -170 190887 -142
rect 190577 -204 190887 -170
rect 190577 -232 190625 -204
rect 190653 -232 190687 -204
rect 190715 -232 190749 -204
rect 190777 -232 190811 -204
rect 190839 -232 190887 -204
rect 190577 -266 190887 -232
rect 190577 -294 190625 -266
rect 190653 -294 190687 -266
rect 190715 -294 190749 -266
rect 190777 -294 190811 -266
rect 190839 -294 190887 -266
rect 190577 -822 190887 -294
rect 192437 299086 192747 299134
rect 192437 299058 192485 299086
rect 192513 299058 192547 299086
rect 192575 299058 192609 299086
rect 192637 299058 192671 299086
rect 192699 299058 192747 299086
rect 192437 299024 192747 299058
rect 192437 298996 192485 299024
rect 192513 298996 192547 299024
rect 192575 298996 192609 299024
rect 192637 298996 192671 299024
rect 192699 298996 192747 299024
rect 192437 298962 192747 298996
rect 192437 298934 192485 298962
rect 192513 298934 192547 298962
rect 192575 298934 192609 298962
rect 192637 298934 192671 298962
rect 192699 298934 192747 298962
rect 192437 298900 192747 298934
rect 192437 298872 192485 298900
rect 192513 298872 192547 298900
rect 192575 298872 192609 298900
rect 192637 298872 192671 298900
rect 192699 298872 192747 298900
rect 192437 293175 192747 298872
rect 192437 293147 192485 293175
rect 192513 293147 192547 293175
rect 192575 293147 192609 293175
rect 192637 293147 192671 293175
rect 192699 293147 192747 293175
rect 192437 293113 192747 293147
rect 192437 293085 192485 293113
rect 192513 293085 192547 293113
rect 192575 293085 192609 293113
rect 192637 293085 192671 293113
rect 192699 293085 192747 293113
rect 192437 293051 192747 293085
rect 192437 293023 192485 293051
rect 192513 293023 192547 293051
rect 192575 293023 192609 293051
rect 192637 293023 192671 293051
rect 192699 293023 192747 293051
rect 192437 292989 192747 293023
rect 192437 292961 192485 292989
rect 192513 292961 192547 292989
rect 192575 292961 192609 292989
rect 192637 292961 192671 292989
rect 192699 292961 192747 292989
rect 192437 284175 192747 292961
rect 192437 284147 192485 284175
rect 192513 284147 192547 284175
rect 192575 284147 192609 284175
rect 192637 284147 192671 284175
rect 192699 284147 192747 284175
rect 192437 284113 192747 284147
rect 192437 284085 192485 284113
rect 192513 284085 192547 284113
rect 192575 284085 192609 284113
rect 192637 284085 192671 284113
rect 192699 284085 192747 284113
rect 192437 284051 192747 284085
rect 192437 284023 192485 284051
rect 192513 284023 192547 284051
rect 192575 284023 192609 284051
rect 192637 284023 192671 284051
rect 192699 284023 192747 284051
rect 192437 283989 192747 284023
rect 192437 283961 192485 283989
rect 192513 283961 192547 283989
rect 192575 283961 192609 283989
rect 192637 283961 192671 283989
rect 192699 283961 192747 283989
rect 192437 275175 192747 283961
rect 192437 275147 192485 275175
rect 192513 275147 192547 275175
rect 192575 275147 192609 275175
rect 192637 275147 192671 275175
rect 192699 275147 192747 275175
rect 192437 275113 192747 275147
rect 192437 275085 192485 275113
rect 192513 275085 192547 275113
rect 192575 275085 192609 275113
rect 192637 275085 192671 275113
rect 192699 275085 192747 275113
rect 192437 275051 192747 275085
rect 192437 275023 192485 275051
rect 192513 275023 192547 275051
rect 192575 275023 192609 275051
rect 192637 275023 192671 275051
rect 192699 275023 192747 275051
rect 192437 274989 192747 275023
rect 192437 274961 192485 274989
rect 192513 274961 192547 274989
rect 192575 274961 192609 274989
rect 192637 274961 192671 274989
rect 192699 274961 192747 274989
rect 192437 266175 192747 274961
rect 192437 266147 192485 266175
rect 192513 266147 192547 266175
rect 192575 266147 192609 266175
rect 192637 266147 192671 266175
rect 192699 266147 192747 266175
rect 192437 266113 192747 266147
rect 192437 266085 192485 266113
rect 192513 266085 192547 266113
rect 192575 266085 192609 266113
rect 192637 266085 192671 266113
rect 192699 266085 192747 266113
rect 192437 266051 192747 266085
rect 192437 266023 192485 266051
rect 192513 266023 192547 266051
rect 192575 266023 192609 266051
rect 192637 266023 192671 266051
rect 192699 266023 192747 266051
rect 192437 265989 192747 266023
rect 192437 265961 192485 265989
rect 192513 265961 192547 265989
rect 192575 265961 192609 265989
rect 192637 265961 192671 265989
rect 192699 265961 192747 265989
rect 192437 257175 192747 265961
rect 192437 257147 192485 257175
rect 192513 257147 192547 257175
rect 192575 257147 192609 257175
rect 192637 257147 192671 257175
rect 192699 257147 192747 257175
rect 192437 257113 192747 257147
rect 192437 257085 192485 257113
rect 192513 257085 192547 257113
rect 192575 257085 192609 257113
rect 192637 257085 192671 257113
rect 192699 257085 192747 257113
rect 192437 257051 192747 257085
rect 192437 257023 192485 257051
rect 192513 257023 192547 257051
rect 192575 257023 192609 257051
rect 192637 257023 192671 257051
rect 192699 257023 192747 257051
rect 192437 256989 192747 257023
rect 192437 256961 192485 256989
rect 192513 256961 192547 256989
rect 192575 256961 192609 256989
rect 192637 256961 192671 256989
rect 192699 256961 192747 256989
rect 192437 248175 192747 256961
rect 192437 248147 192485 248175
rect 192513 248147 192547 248175
rect 192575 248147 192609 248175
rect 192637 248147 192671 248175
rect 192699 248147 192747 248175
rect 192437 248113 192747 248147
rect 192437 248085 192485 248113
rect 192513 248085 192547 248113
rect 192575 248085 192609 248113
rect 192637 248085 192671 248113
rect 192699 248085 192747 248113
rect 192437 248051 192747 248085
rect 192437 248023 192485 248051
rect 192513 248023 192547 248051
rect 192575 248023 192609 248051
rect 192637 248023 192671 248051
rect 192699 248023 192747 248051
rect 192437 247989 192747 248023
rect 192437 247961 192485 247989
rect 192513 247961 192547 247989
rect 192575 247961 192609 247989
rect 192637 247961 192671 247989
rect 192699 247961 192747 247989
rect 192437 239175 192747 247961
rect 192437 239147 192485 239175
rect 192513 239147 192547 239175
rect 192575 239147 192609 239175
rect 192637 239147 192671 239175
rect 192699 239147 192747 239175
rect 192437 239113 192747 239147
rect 192437 239085 192485 239113
rect 192513 239085 192547 239113
rect 192575 239085 192609 239113
rect 192637 239085 192671 239113
rect 192699 239085 192747 239113
rect 192437 239051 192747 239085
rect 192437 239023 192485 239051
rect 192513 239023 192547 239051
rect 192575 239023 192609 239051
rect 192637 239023 192671 239051
rect 192699 239023 192747 239051
rect 192437 238989 192747 239023
rect 192437 238961 192485 238989
rect 192513 238961 192547 238989
rect 192575 238961 192609 238989
rect 192637 238961 192671 238989
rect 192699 238961 192747 238989
rect 192437 230175 192747 238961
rect 192437 230147 192485 230175
rect 192513 230147 192547 230175
rect 192575 230147 192609 230175
rect 192637 230147 192671 230175
rect 192699 230147 192747 230175
rect 192437 230113 192747 230147
rect 192437 230085 192485 230113
rect 192513 230085 192547 230113
rect 192575 230085 192609 230113
rect 192637 230085 192671 230113
rect 192699 230085 192747 230113
rect 192437 230051 192747 230085
rect 192437 230023 192485 230051
rect 192513 230023 192547 230051
rect 192575 230023 192609 230051
rect 192637 230023 192671 230051
rect 192699 230023 192747 230051
rect 192437 229989 192747 230023
rect 192437 229961 192485 229989
rect 192513 229961 192547 229989
rect 192575 229961 192609 229989
rect 192637 229961 192671 229989
rect 192699 229961 192747 229989
rect 192437 221175 192747 229961
rect 192437 221147 192485 221175
rect 192513 221147 192547 221175
rect 192575 221147 192609 221175
rect 192637 221147 192671 221175
rect 192699 221147 192747 221175
rect 192437 221113 192747 221147
rect 192437 221085 192485 221113
rect 192513 221085 192547 221113
rect 192575 221085 192609 221113
rect 192637 221085 192671 221113
rect 192699 221085 192747 221113
rect 192437 221051 192747 221085
rect 192437 221023 192485 221051
rect 192513 221023 192547 221051
rect 192575 221023 192609 221051
rect 192637 221023 192671 221051
rect 192699 221023 192747 221051
rect 192437 220989 192747 221023
rect 192437 220961 192485 220989
rect 192513 220961 192547 220989
rect 192575 220961 192609 220989
rect 192637 220961 192671 220989
rect 192699 220961 192747 220989
rect 192437 212175 192747 220961
rect 192437 212147 192485 212175
rect 192513 212147 192547 212175
rect 192575 212147 192609 212175
rect 192637 212147 192671 212175
rect 192699 212147 192747 212175
rect 192437 212113 192747 212147
rect 192437 212085 192485 212113
rect 192513 212085 192547 212113
rect 192575 212085 192609 212113
rect 192637 212085 192671 212113
rect 192699 212085 192747 212113
rect 192437 212051 192747 212085
rect 192437 212023 192485 212051
rect 192513 212023 192547 212051
rect 192575 212023 192609 212051
rect 192637 212023 192671 212051
rect 192699 212023 192747 212051
rect 192437 211989 192747 212023
rect 192437 211961 192485 211989
rect 192513 211961 192547 211989
rect 192575 211961 192609 211989
rect 192637 211961 192671 211989
rect 192699 211961 192747 211989
rect 192437 203175 192747 211961
rect 192437 203147 192485 203175
rect 192513 203147 192547 203175
rect 192575 203147 192609 203175
rect 192637 203147 192671 203175
rect 192699 203147 192747 203175
rect 192437 203113 192747 203147
rect 192437 203085 192485 203113
rect 192513 203085 192547 203113
rect 192575 203085 192609 203113
rect 192637 203085 192671 203113
rect 192699 203085 192747 203113
rect 192437 203051 192747 203085
rect 192437 203023 192485 203051
rect 192513 203023 192547 203051
rect 192575 203023 192609 203051
rect 192637 203023 192671 203051
rect 192699 203023 192747 203051
rect 192437 202989 192747 203023
rect 192437 202961 192485 202989
rect 192513 202961 192547 202989
rect 192575 202961 192609 202989
rect 192637 202961 192671 202989
rect 192699 202961 192747 202989
rect 192437 194175 192747 202961
rect 192437 194147 192485 194175
rect 192513 194147 192547 194175
rect 192575 194147 192609 194175
rect 192637 194147 192671 194175
rect 192699 194147 192747 194175
rect 192437 194113 192747 194147
rect 192437 194085 192485 194113
rect 192513 194085 192547 194113
rect 192575 194085 192609 194113
rect 192637 194085 192671 194113
rect 192699 194085 192747 194113
rect 192437 194051 192747 194085
rect 192437 194023 192485 194051
rect 192513 194023 192547 194051
rect 192575 194023 192609 194051
rect 192637 194023 192671 194051
rect 192699 194023 192747 194051
rect 192437 193989 192747 194023
rect 192437 193961 192485 193989
rect 192513 193961 192547 193989
rect 192575 193961 192609 193989
rect 192637 193961 192671 193989
rect 192699 193961 192747 193989
rect 192437 185175 192747 193961
rect 192437 185147 192485 185175
rect 192513 185147 192547 185175
rect 192575 185147 192609 185175
rect 192637 185147 192671 185175
rect 192699 185147 192747 185175
rect 192437 185113 192747 185147
rect 192437 185085 192485 185113
rect 192513 185085 192547 185113
rect 192575 185085 192609 185113
rect 192637 185085 192671 185113
rect 192699 185085 192747 185113
rect 192437 185051 192747 185085
rect 192437 185023 192485 185051
rect 192513 185023 192547 185051
rect 192575 185023 192609 185051
rect 192637 185023 192671 185051
rect 192699 185023 192747 185051
rect 192437 184989 192747 185023
rect 192437 184961 192485 184989
rect 192513 184961 192547 184989
rect 192575 184961 192609 184989
rect 192637 184961 192671 184989
rect 192699 184961 192747 184989
rect 192437 176175 192747 184961
rect 192437 176147 192485 176175
rect 192513 176147 192547 176175
rect 192575 176147 192609 176175
rect 192637 176147 192671 176175
rect 192699 176147 192747 176175
rect 192437 176113 192747 176147
rect 192437 176085 192485 176113
rect 192513 176085 192547 176113
rect 192575 176085 192609 176113
rect 192637 176085 192671 176113
rect 192699 176085 192747 176113
rect 192437 176051 192747 176085
rect 192437 176023 192485 176051
rect 192513 176023 192547 176051
rect 192575 176023 192609 176051
rect 192637 176023 192671 176051
rect 192699 176023 192747 176051
rect 192437 175989 192747 176023
rect 192437 175961 192485 175989
rect 192513 175961 192547 175989
rect 192575 175961 192609 175989
rect 192637 175961 192671 175989
rect 192699 175961 192747 175989
rect 192437 167175 192747 175961
rect 192437 167147 192485 167175
rect 192513 167147 192547 167175
rect 192575 167147 192609 167175
rect 192637 167147 192671 167175
rect 192699 167147 192747 167175
rect 192437 167113 192747 167147
rect 192437 167085 192485 167113
rect 192513 167085 192547 167113
rect 192575 167085 192609 167113
rect 192637 167085 192671 167113
rect 192699 167085 192747 167113
rect 192437 167051 192747 167085
rect 192437 167023 192485 167051
rect 192513 167023 192547 167051
rect 192575 167023 192609 167051
rect 192637 167023 192671 167051
rect 192699 167023 192747 167051
rect 192437 166989 192747 167023
rect 192437 166961 192485 166989
rect 192513 166961 192547 166989
rect 192575 166961 192609 166989
rect 192637 166961 192671 166989
rect 192699 166961 192747 166989
rect 192437 158175 192747 166961
rect 192437 158147 192485 158175
rect 192513 158147 192547 158175
rect 192575 158147 192609 158175
rect 192637 158147 192671 158175
rect 192699 158147 192747 158175
rect 192437 158113 192747 158147
rect 192437 158085 192485 158113
rect 192513 158085 192547 158113
rect 192575 158085 192609 158113
rect 192637 158085 192671 158113
rect 192699 158085 192747 158113
rect 192437 158051 192747 158085
rect 192437 158023 192485 158051
rect 192513 158023 192547 158051
rect 192575 158023 192609 158051
rect 192637 158023 192671 158051
rect 192699 158023 192747 158051
rect 192437 157989 192747 158023
rect 192437 157961 192485 157989
rect 192513 157961 192547 157989
rect 192575 157961 192609 157989
rect 192637 157961 192671 157989
rect 192699 157961 192747 157989
rect 192437 149175 192747 157961
rect 192437 149147 192485 149175
rect 192513 149147 192547 149175
rect 192575 149147 192609 149175
rect 192637 149147 192671 149175
rect 192699 149147 192747 149175
rect 192437 149113 192747 149147
rect 192437 149085 192485 149113
rect 192513 149085 192547 149113
rect 192575 149085 192609 149113
rect 192637 149085 192671 149113
rect 192699 149085 192747 149113
rect 192437 149051 192747 149085
rect 192437 149023 192485 149051
rect 192513 149023 192547 149051
rect 192575 149023 192609 149051
rect 192637 149023 192671 149051
rect 192699 149023 192747 149051
rect 192437 148989 192747 149023
rect 192437 148961 192485 148989
rect 192513 148961 192547 148989
rect 192575 148961 192609 148989
rect 192637 148961 192671 148989
rect 192699 148961 192747 148989
rect 192437 140175 192747 148961
rect 192437 140147 192485 140175
rect 192513 140147 192547 140175
rect 192575 140147 192609 140175
rect 192637 140147 192671 140175
rect 192699 140147 192747 140175
rect 192437 140113 192747 140147
rect 192437 140085 192485 140113
rect 192513 140085 192547 140113
rect 192575 140085 192609 140113
rect 192637 140085 192671 140113
rect 192699 140085 192747 140113
rect 192437 140051 192747 140085
rect 192437 140023 192485 140051
rect 192513 140023 192547 140051
rect 192575 140023 192609 140051
rect 192637 140023 192671 140051
rect 192699 140023 192747 140051
rect 192437 139989 192747 140023
rect 192437 139961 192485 139989
rect 192513 139961 192547 139989
rect 192575 139961 192609 139989
rect 192637 139961 192671 139989
rect 192699 139961 192747 139989
rect 192437 131175 192747 139961
rect 192437 131147 192485 131175
rect 192513 131147 192547 131175
rect 192575 131147 192609 131175
rect 192637 131147 192671 131175
rect 192699 131147 192747 131175
rect 192437 131113 192747 131147
rect 192437 131085 192485 131113
rect 192513 131085 192547 131113
rect 192575 131085 192609 131113
rect 192637 131085 192671 131113
rect 192699 131085 192747 131113
rect 192437 131051 192747 131085
rect 192437 131023 192485 131051
rect 192513 131023 192547 131051
rect 192575 131023 192609 131051
rect 192637 131023 192671 131051
rect 192699 131023 192747 131051
rect 192437 130989 192747 131023
rect 192437 130961 192485 130989
rect 192513 130961 192547 130989
rect 192575 130961 192609 130989
rect 192637 130961 192671 130989
rect 192699 130961 192747 130989
rect 192437 122175 192747 130961
rect 192437 122147 192485 122175
rect 192513 122147 192547 122175
rect 192575 122147 192609 122175
rect 192637 122147 192671 122175
rect 192699 122147 192747 122175
rect 192437 122113 192747 122147
rect 192437 122085 192485 122113
rect 192513 122085 192547 122113
rect 192575 122085 192609 122113
rect 192637 122085 192671 122113
rect 192699 122085 192747 122113
rect 192437 122051 192747 122085
rect 192437 122023 192485 122051
rect 192513 122023 192547 122051
rect 192575 122023 192609 122051
rect 192637 122023 192671 122051
rect 192699 122023 192747 122051
rect 192437 121989 192747 122023
rect 192437 121961 192485 121989
rect 192513 121961 192547 121989
rect 192575 121961 192609 121989
rect 192637 121961 192671 121989
rect 192699 121961 192747 121989
rect 192437 113175 192747 121961
rect 192437 113147 192485 113175
rect 192513 113147 192547 113175
rect 192575 113147 192609 113175
rect 192637 113147 192671 113175
rect 192699 113147 192747 113175
rect 192437 113113 192747 113147
rect 192437 113085 192485 113113
rect 192513 113085 192547 113113
rect 192575 113085 192609 113113
rect 192637 113085 192671 113113
rect 192699 113085 192747 113113
rect 192437 113051 192747 113085
rect 192437 113023 192485 113051
rect 192513 113023 192547 113051
rect 192575 113023 192609 113051
rect 192637 113023 192671 113051
rect 192699 113023 192747 113051
rect 192437 112989 192747 113023
rect 192437 112961 192485 112989
rect 192513 112961 192547 112989
rect 192575 112961 192609 112989
rect 192637 112961 192671 112989
rect 192699 112961 192747 112989
rect 192437 104175 192747 112961
rect 192437 104147 192485 104175
rect 192513 104147 192547 104175
rect 192575 104147 192609 104175
rect 192637 104147 192671 104175
rect 192699 104147 192747 104175
rect 192437 104113 192747 104147
rect 192437 104085 192485 104113
rect 192513 104085 192547 104113
rect 192575 104085 192609 104113
rect 192637 104085 192671 104113
rect 192699 104085 192747 104113
rect 192437 104051 192747 104085
rect 192437 104023 192485 104051
rect 192513 104023 192547 104051
rect 192575 104023 192609 104051
rect 192637 104023 192671 104051
rect 192699 104023 192747 104051
rect 192437 103989 192747 104023
rect 192437 103961 192485 103989
rect 192513 103961 192547 103989
rect 192575 103961 192609 103989
rect 192637 103961 192671 103989
rect 192699 103961 192747 103989
rect 192437 95175 192747 103961
rect 192437 95147 192485 95175
rect 192513 95147 192547 95175
rect 192575 95147 192609 95175
rect 192637 95147 192671 95175
rect 192699 95147 192747 95175
rect 192437 95113 192747 95147
rect 192437 95085 192485 95113
rect 192513 95085 192547 95113
rect 192575 95085 192609 95113
rect 192637 95085 192671 95113
rect 192699 95085 192747 95113
rect 192437 95051 192747 95085
rect 192437 95023 192485 95051
rect 192513 95023 192547 95051
rect 192575 95023 192609 95051
rect 192637 95023 192671 95051
rect 192699 95023 192747 95051
rect 192437 94989 192747 95023
rect 192437 94961 192485 94989
rect 192513 94961 192547 94989
rect 192575 94961 192609 94989
rect 192637 94961 192671 94989
rect 192699 94961 192747 94989
rect 192437 86175 192747 94961
rect 192437 86147 192485 86175
rect 192513 86147 192547 86175
rect 192575 86147 192609 86175
rect 192637 86147 192671 86175
rect 192699 86147 192747 86175
rect 192437 86113 192747 86147
rect 192437 86085 192485 86113
rect 192513 86085 192547 86113
rect 192575 86085 192609 86113
rect 192637 86085 192671 86113
rect 192699 86085 192747 86113
rect 192437 86051 192747 86085
rect 192437 86023 192485 86051
rect 192513 86023 192547 86051
rect 192575 86023 192609 86051
rect 192637 86023 192671 86051
rect 192699 86023 192747 86051
rect 192437 85989 192747 86023
rect 192437 85961 192485 85989
rect 192513 85961 192547 85989
rect 192575 85961 192609 85989
rect 192637 85961 192671 85989
rect 192699 85961 192747 85989
rect 192437 77175 192747 85961
rect 192437 77147 192485 77175
rect 192513 77147 192547 77175
rect 192575 77147 192609 77175
rect 192637 77147 192671 77175
rect 192699 77147 192747 77175
rect 192437 77113 192747 77147
rect 192437 77085 192485 77113
rect 192513 77085 192547 77113
rect 192575 77085 192609 77113
rect 192637 77085 192671 77113
rect 192699 77085 192747 77113
rect 192437 77051 192747 77085
rect 192437 77023 192485 77051
rect 192513 77023 192547 77051
rect 192575 77023 192609 77051
rect 192637 77023 192671 77051
rect 192699 77023 192747 77051
rect 192437 76989 192747 77023
rect 192437 76961 192485 76989
rect 192513 76961 192547 76989
rect 192575 76961 192609 76989
rect 192637 76961 192671 76989
rect 192699 76961 192747 76989
rect 192437 68175 192747 76961
rect 192437 68147 192485 68175
rect 192513 68147 192547 68175
rect 192575 68147 192609 68175
rect 192637 68147 192671 68175
rect 192699 68147 192747 68175
rect 192437 68113 192747 68147
rect 192437 68085 192485 68113
rect 192513 68085 192547 68113
rect 192575 68085 192609 68113
rect 192637 68085 192671 68113
rect 192699 68085 192747 68113
rect 192437 68051 192747 68085
rect 192437 68023 192485 68051
rect 192513 68023 192547 68051
rect 192575 68023 192609 68051
rect 192637 68023 192671 68051
rect 192699 68023 192747 68051
rect 192437 67989 192747 68023
rect 192437 67961 192485 67989
rect 192513 67961 192547 67989
rect 192575 67961 192609 67989
rect 192637 67961 192671 67989
rect 192699 67961 192747 67989
rect 192437 59175 192747 67961
rect 192437 59147 192485 59175
rect 192513 59147 192547 59175
rect 192575 59147 192609 59175
rect 192637 59147 192671 59175
rect 192699 59147 192747 59175
rect 192437 59113 192747 59147
rect 192437 59085 192485 59113
rect 192513 59085 192547 59113
rect 192575 59085 192609 59113
rect 192637 59085 192671 59113
rect 192699 59085 192747 59113
rect 192437 59051 192747 59085
rect 192437 59023 192485 59051
rect 192513 59023 192547 59051
rect 192575 59023 192609 59051
rect 192637 59023 192671 59051
rect 192699 59023 192747 59051
rect 192437 58989 192747 59023
rect 192437 58961 192485 58989
rect 192513 58961 192547 58989
rect 192575 58961 192609 58989
rect 192637 58961 192671 58989
rect 192699 58961 192747 58989
rect 192437 50175 192747 58961
rect 192437 50147 192485 50175
rect 192513 50147 192547 50175
rect 192575 50147 192609 50175
rect 192637 50147 192671 50175
rect 192699 50147 192747 50175
rect 192437 50113 192747 50147
rect 192437 50085 192485 50113
rect 192513 50085 192547 50113
rect 192575 50085 192609 50113
rect 192637 50085 192671 50113
rect 192699 50085 192747 50113
rect 192437 50051 192747 50085
rect 192437 50023 192485 50051
rect 192513 50023 192547 50051
rect 192575 50023 192609 50051
rect 192637 50023 192671 50051
rect 192699 50023 192747 50051
rect 192437 49989 192747 50023
rect 192437 49961 192485 49989
rect 192513 49961 192547 49989
rect 192575 49961 192609 49989
rect 192637 49961 192671 49989
rect 192699 49961 192747 49989
rect 192437 41175 192747 49961
rect 192437 41147 192485 41175
rect 192513 41147 192547 41175
rect 192575 41147 192609 41175
rect 192637 41147 192671 41175
rect 192699 41147 192747 41175
rect 192437 41113 192747 41147
rect 192437 41085 192485 41113
rect 192513 41085 192547 41113
rect 192575 41085 192609 41113
rect 192637 41085 192671 41113
rect 192699 41085 192747 41113
rect 192437 41051 192747 41085
rect 192437 41023 192485 41051
rect 192513 41023 192547 41051
rect 192575 41023 192609 41051
rect 192637 41023 192671 41051
rect 192699 41023 192747 41051
rect 192437 40989 192747 41023
rect 192437 40961 192485 40989
rect 192513 40961 192547 40989
rect 192575 40961 192609 40989
rect 192637 40961 192671 40989
rect 192699 40961 192747 40989
rect 192437 32175 192747 40961
rect 192437 32147 192485 32175
rect 192513 32147 192547 32175
rect 192575 32147 192609 32175
rect 192637 32147 192671 32175
rect 192699 32147 192747 32175
rect 192437 32113 192747 32147
rect 192437 32085 192485 32113
rect 192513 32085 192547 32113
rect 192575 32085 192609 32113
rect 192637 32085 192671 32113
rect 192699 32085 192747 32113
rect 192437 32051 192747 32085
rect 192437 32023 192485 32051
rect 192513 32023 192547 32051
rect 192575 32023 192609 32051
rect 192637 32023 192671 32051
rect 192699 32023 192747 32051
rect 192437 31989 192747 32023
rect 192437 31961 192485 31989
rect 192513 31961 192547 31989
rect 192575 31961 192609 31989
rect 192637 31961 192671 31989
rect 192699 31961 192747 31989
rect 192437 23175 192747 31961
rect 192437 23147 192485 23175
rect 192513 23147 192547 23175
rect 192575 23147 192609 23175
rect 192637 23147 192671 23175
rect 192699 23147 192747 23175
rect 192437 23113 192747 23147
rect 192437 23085 192485 23113
rect 192513 23085 192547 23113
rect 192575 23085 192609 23113
rect 192637 23085 192671 23113
rect 192699 23085 192747 23113
rect 192437 23051 192747 23085
rect 192437 23023 192485 23051
rect 192513 23023 192547 23051
rect 192575 23023 192609 23051
rect 192637 23023 192671 23051
rect 192699 23023 192747 23051
rect 192437 22989 192747 23023
rect 192437 22961 192485 22989
rect 192513 22961 192547 22989
rect 192575 22961 192609 22989
rect 192637 22961 192671 22989
rect 192699 22961 192747 22989
rect 192437 14175 192747 22961
rect 192437 14147 192485 14175
rect 192513 14147 192547 14175
rect 192575 14147 192609 14175
rect 192637 14147 192671 14175
rect 192699 14147 192747 14175
rect 192437 14113 192747 14147
rect 192437 14085 192485 14113
rect 192513 14085 192547 14113
rect 192575 14085 192609 14113
rect 192637 14085 192671 14113
rect 192699 14085 192747 14113
rect 192437 14051 192747 14085
rect 192437 14023 192485 14051
rect 192513 14023 192547 14051
rect 192575 14023 192609 14051
rect 192637 14023 192671 14051
rect 192699 14023 192747 14051
rect 192437 13989 192747 14023
rect 192437 13961 192485 13989
rect 192513 13961 192547 13989
rect 192575 13961 192609 13989
rect 192637 13961 192671 13989
rect 192699 13961 192747 13989
rect 192437 5175 192747 13961
rect 192437 5147 192485 5175
rect 192513 5147 192547 5175
rect 192575 5147 192609 5175
rect 192637 5147 192671 5175
rect 192699 5147 192747 5175
rect 192437 5113 192747 5147
rect 192437 5085 192485 5113
rect 192513 5085 192547 5113
rect 192575 5085 192609 5113
rect 192637 5085 192671 5113
rect 192699 5085 192747 5113
rect 192437 5051 192747 5085
rect 192437 5023 192485 5051
rect 192513 5023 192547 5051
rect 192575 5023 192609 5051
rect 192637 5023 192671 5051
rect 192699 5023 192747 5051
rect 192437 4989 192747 5023
rect 192437 4961 192485 4989
rect 192513 4961 192547 4989
rect 192575 4961 192609 4989
rect 192637 4961 192671 4989
rect 192699 4961 192747 4989
rect 192437 -560 192747 4961
rect 192437 -588 192485 -560
rect 192513 -588 192547 -560
rect 192575 -588 192609 -560
rect 192637 -588 192671 -560
rect 192699 -588 192747 -560
rect 192437 -622 192747 -588
rect 192437 -650 192485 -622
rect 192513 -650 192547 -622
rect 192575 -650 192609 -622
rect 192637 -650 192671 -622
rect 192699 -650 192747 -622
rect 192437 -684 192747 -650
rect 192437 -712 192485 -684
rect 192513 -712 192547 -684
rect 192575 -712 192609 -684
rect 192637 -712 192671 -684
rect 192699 -712 192747 -684
rect 192437 -746 192747 -712
rect 192437 -774 192485 -746
rect 192513 -774 192547 -746
rect 192575 -774 192609 -746
rect 192637 -774 192671 -746
rect 192699 -774 192747 -746
rect 192437 -822 192747 -774
rect 199577 298606 199887 299134
rect 199577 298578 199625 298606
rect 199653 298578 199687 298606
rect 199715 298578 199749 298606
rect 199777 298578 199811 298606
rect 199839 298578 199887 298606
rect 199577 298544 199887 298578
rect 199577 298516 199625 298544
rect 199653 298516 199687 298544
rect 199715 298516 199749 298544
rect 199777 298516 199811 298544
rect 199839 298516 199887 298544
rect 199577 298482 199887 298516
rect 199577 298454 199625 298482
rect 199653 298454 199687 298482
rect 199715 298454 199749 298482
rect 199777 298454 199811 298482
rect 199839 298454 199887 298482
rect 199577 298420 199887 298454
rect 199577 298392 199625 298420
rect 199653 298392 199687 298420
rect 199715 298392 199749 298420
rect 199777 298392 199811 298420
rect 199839 298392 199887 298420
rect 199577 290175 199887 298392
rect 199577 290147 199625 290175
rect 199653 290147 199687 290175
rect 199715 290147 199749 290175
rect 199777 290147 199811 290175
rect 199839 290147 199887 290175
rect 199577 290113 199887 290147
rect 199577 290085 199625 290113
rect 199653 290085 199687 290113
rect 199715 290085 199749 290113
rect 199777 290085 199811 290113
rect 199839 290085 199887 290113
rect 199577 290051 199887 290085
rect 199577 290023 199625 290051
rect 199653 290023 199687 290051
rect 199715 290023 199749 290051
rect 199777 290023 199811 290051
rect 199839 290023 199887 290051
rect 199577 289989 199887 290023
rect 199577 289961 199625 289989
rect 199653 289961 199687 289989
rect 199715 289961 199749 289989
rect 199777 289961 199811 289989
rect 199839 289961 199887 289989
rect 199577 281175 199887 289961
rect 199577 281147 199625 281175
rect 199653 281147 199687 281175
rect 199715 281147 199749 281175
rect 199777 281147 199811 281175
rect 199839 281147 199887 281175
rect 199577 281113 199887 281147
rect 199577 281085 199625 281113
rect 199653 281085 199687 281113
rect 199715 281085 199749 281113
rect 199777 281085 199811 281113
rect 199839 281085 199887 281113
rect 199577 281051 199887 281085
rect 199577 281023 199625 281051
rect 199653 281023 199687 281051
rect 199715 281023 199749 281051
rect 199777 281023 199811 281051
rect 199839 281023 199887 281051
rect 199577 280989 199887 281023
rect 199577 280961 199625 280989
rect 199653 280961 199687 280989
rect 199715 280961 199749 280989
rect 199777 280961 199811 280989
rect 199839 280961 199887 280989
rect 199577 272175 199887 280961
rect 199577 272147 199625 272175
rect 199653 272147 199687 272175
rect 199715 272147 199749 272175
rect 199777 272147 199811 272175
rect 199839 272147 199887 272175
rect 199577 272113 199887 272147
rect 199577 272085 199625 272113
rect 199653 272085 199687 272113
rect 199715 272085 199749 272113
rect 199777 272085 199811 272113
rect 199839 272085 199887 272113
rect 199577 272051 199887 272085
rect 199577 272023 199625 272051
rect 199653 272023 199687 272051
rect 199715 272023 199749 272051
rect 199777 272023 199811 272051
rect 199839 272023 199887 272051
rect 199577 271989 199887 272023
rect 199577 271961 199625 271989
rect 199653 271961 199687 271989
rect 199715 271961 199749 271989
rect 199777 271961 199811 271989
rect 199839 271961 199887 271989
rect 199577 263175 199887 271961
rect 199577 263147 199625 263175
rect 199653 263147 199687 263175
rect 199715 263147 199749 263175
rect 199777 263147 199811 263175
rect 199839 263147 199887 263175
rect 199577 263113 199887 263147
rect 199577 263085 199625 263113
rect 199653 263085 199687 263113
rect 199715 263085 199749 263113
rect 199777 263085 199811 263113
rect 199839 263085 199887 263113
rect 199577 263051 199887 263085
rect 199577 263023 199625 263051
rect 199653 263023 199687 263051
rect 199715 263023 199749 263051
rect 199777 263023 199811 263051
rect 199839 263023 199887 263051
rect 199577 262989 199887 263023
rect 199577 262961 199625 262989
rect 199653 262961 199687 262989
rect 199715 262961 199749 262989
rect 199777 262961 199811 262989
rect 199839 262961 199887 262989
rect 199577 254175 199887 262961
rect 199577 254147 199625 254175
rect 199653 254147 199687 254175
rect 199715 254147 199749 254175
rect 199777 254147 199811 254175
rect 199839 254147 199887 254175
rect 199577 254113 199887 254147
rect 199577 254085 199625 254113
rect 199653 254085 199687 254113
rect 199715 254085 199749 254113
rect 199777 254085 199811 254113
rect 199839 254085 199887 254113
rect 199577 254051 199887 254085
rect 199577 254023 199625 254051
rect 199653 254023 199687 254051
rect 199715 254023 199749 254051
rect 199777 254023 199811 254051
rect 199839 254023 199887 254051
rect 199577 253989 199887 254023
rect 199577 253961 199625 253989
rect 199653 253961 199687 253989
rect 199715 253961 199749 253989
rect 199777 253961 199811 253989
rect 199839 253961 199887 253989
rect 199577 245175 199887 253961
rect 199577 245147 199625 245175
rect 199653 245147 199687 245175
rect 199715 245147 199749 245175
rect 199777 245147 199811 245175
rect 199839 245147 199887 245175
rect 199577 245113 199887 245147
rect 199577 245085 199625 245113
rect 199653 245085 199687 245113
rect 199715 245085 199749 245113
rect 199777 245085 199811 245113
rect 199839 245085 199887 245113
rect 199577 245051 199887 245085
rect 199577 245023 199625 245051
rect 199653 245023 199687 245051
rect 199715 245023 199749 245051
rect 199777 245023 199811 245051
rect 199839 245023 199887 245051
rect 199577 244989 199887 245023
rect 199577 244961 199625 244989
rect 199653 244961 199687 244989
rect 199715 244961 199749 244989
rect 199777 244961 199811 244989
rect 199839 244961 199887 244989
rect 199577 236175 199887 244961
rect 199577 236147 199625 236175
rect 199653 236147 199687 236175
rect 199715 236147 199749 236175
rect 199777 236147 199811 236175
rect 199839 236147 199887 236175
rect 199577 236113 199887 236147
rect 199577 236085 199625 236113
rect 199653 236085 199687 236113
rect 199715 236085 199749 236113
rect 199777 236085 199811 236113
rect 199839 236085 199887 236113
rect 199577 236051 199887 236085
rect 199577 236023 199625 236051
rect 199653 236023 199687 236051
rect 199715 236023 199749 236051
rect 199777 236023 199811 236051
rect 199839 236023 199887 236051
rect 199577 235989 199887 236023
rect 199577 235961 199625 235989
rect 199653 235961 199687 235989
rect 199715 235961 199749 235989
rect 199777 235961 199811 235989
rect 199839 235961 199887 235989
rect 199577 227175 199887 235961
rect 199577 227147 199625 227175
rect 199653 227147 199687 227175
rect 199715 227147 199749 227175
rect 199777 227147 199811 227175
rect 199839 227147 199887 227175
rect 199577 227113 199887 227147
rect 199577 227085 199625 227113
rect 199653 227085 199687 227113
rect 199715 227085 199749 227113
rect 199777 227085 199811 227113
rect 199839 227085 199887 227113
rect 199577 227051 199887 227085
rect 199577 227023 199625 227051
rect 199653 227023 199687 227051
rect 199715 227023 199749 227051
rect 199777 227023 199811 227051
rect 199839 227023 199887 227051
rect 199577 226989 199887 227023
rect 199577 226961 199625 226989
rect 199653 226961 199687 226989
rect 199715 226961 199749 226989
rect 199777 226961 199811 226989
rect 199839 226961 199887 226989
rect 199577 218175 199887 226961
rect 199577 218147 199625 218175
rect 199653 218147 199687 218175
rect 199715 218147 199749 218175
rect 199777 218147 199811 218175
rect 199839 218147 199887 218175
rect 199577 218113 199887 218147
rect 199577 218085 199625 218113
rect 199653 218085 199687 218113
rect 199715 218085 199749 218113
rect 199777 218085 199811 218113
rect 199839 218085 199887 218113
rect 199577 218051 199887 218085
rect 199577 218023 199625 218051
rect 199653 218023 199687 218051
rect 199715 218023 199749 218051
rect 199777 218023 199811 218051
rect 199839 218023 199887 218051
rect 199577 217989 199887 218023
rect 199577 217961 199625 217989
rect 199653 217961 199687 217989
rect 199715 217961 199749 217989
rect 199777 217961 199811 217989
rect 199839 217961 199887 217989
rect 199577 209175 199887 217961
rect 199577 209147 199625 209175
rect 199653 209147 199687 209175
rect 199715 209147 199749 209175
rect 199777 209147 199811 209175
rect 199839 209147 199887 209175
rect 199577 209113 199887 209147
rect 199577 209085 199625 209113
rect 199653 209085 199687 209113
rect 199715 209085 199749 209113
rect 199777 209085 199811 209113
rect 199839 209085 199887 209113
rect 199577 209051 199887 209085
rect 199577 209023 199625 209051
rect 199653 209023 199687 209051
rect 199715 209023 199749 209051
rect 199777 209023 199811 209051
rect 199839 209023 199887 209051
rect 199577 208989 199887 209023
rect 199577 208961 199625 208989
rect 199653 208961 199687 208989
rect 199715 208961 199749 208989
rect 199777 208961 199811 208989
rect 199839 208961 199887 208989
rect 199577 200175 199887 208961
rect 199577 200147 199625 200175
rect 199653 200147 199687 200175
rect 199715 200147 199749 200175
rect 199777 200147 199811 200175
rect 199839 200147 199887 200175
rect 199577 200113 199887 200147
rect 199577 200085 199625 200113
rect 199653 200085 199687 200113
rect 199715 200085 199749 200113
rect 199777 200085 199811 200113
rect 199839 200085 199887 200113
rect 199577 200051 199887 200085
rect 199577 200023 199625 200051
rect 199653 200023 199687 200051
rect 199715 200023 199749 200051
rect 199777 200023 199811 200051
rect 199839 200023 199887 200051
rect 199577 199989 199887 200023
rect 199577 199961 199625 199989
rect 199653 199961 199687 199989
rect 199715 199961 199749 199989
rect 199777 199961 199811 199989
rect 199839 199961 199887 199989
rect 199577 191175 199887 199961
rect 199577 191147 199625 191175
rect 199653 191147 199687 191175
rect 199715 191147 199749 191175
rect 199777 191147 199811 191175
rect 199839 191147 199887 191175
rect 199577 191113 199887 191147
rect 199577 191085 199625 191113
rect 199653 191085 199687 191113
rect 199715 191085 199749 191113
rect 199777 191085 199811 191113
rect 199839 191085 199887 191113
rect 199577 191051 199887 191085
rect 199577 191023 199625 191051
rect 199653 191023 199687 191051
rect 199715 191023 199749 191051
rect 199777 191023 199811 191051
rect 199839 191023 199887 191051
rect 199577 190989 199887 191023
rect 199577 190961 199625 190989
rect 199653 190961 199687 190989
rect 199715 190961 199749 190989
rect 199777 190961 199811 190989
rect 199839 190961 199887 190989
rect 199577 182175 199887 190961
rect 199577 182147 199625 182175
rect 199653 182147 199687 182175
rect 199715 182147 199749 182175
rect 199777 182147 199811 182175
rect 199839 182147 199887 182175
rect 199577 182113 199887 182147
rect 199577 182085 199625 182113
rect 199653 182085 199687 182113
rect 199715 182085 199749 182113
rect 199777 182085 199811 182113
rect 199839 182085 199887 182113
rect 199577 182051 199887 182085
rect 199577 182023 199625 182051
rect 199653 182023 199687 182051
rect 199715 182023 199749 182051
rect 199777 182023 199811 182051
rect 199839 182023 199887 182051
rect 199577 181989 199887 182023
rect 199577 181961 199625 181989
rect 199653 181961 199687 181989
rect 199715 181961 199749 181989
rect 199777 181961 199811 181989
rect 199839 181961 199887 181989
rect 199577 173175 199887 181961
rect 199577 173147 199625 173175
rect 199653 173147 199687 173175
rect 199715 173147 199749 173175
rect 199777 173147 199811 173175
rect 199839 173147 199887 173175
rect 199577 173113 199887 173147
rect 199577 173085 199625 173113
rect 199653 173085 199687 173113
rect 199715 173085 199749 173113
rect 199777 173085 199811 173113
rect 199839 173085 199887 173113
rect 199577 173051 199887 173085
rect 199577 173023 199625 173051
rect 199653 173023 199687 173051
rect 199715 173023 199749 173051
rect 199777 173023 199811 173051
rect 199839 173023 199887 173051
rect 199577 172989 199887 173023
rect 199577 172961 199625 172989
rect 199653 172961 199687 172989
rect 199715 172961 199749 172989
rect 199777 172961 199811 172989
rect 199839 172961 199887 172989
rect 199577 164175 199887 172961
rect 199577 164147 199625 164175
rect 199653 164147 199687 164175
rect 199715 164147 199749 164175
rect 199777 164147 199811 164175
rect 199839 164147 199887 164175
rect 199577 164113 199887 164147
rect 199577 164085 199625 164113
rect 199653 164085 199687 164113
rect 199715 164085 199749 164113
rect 199777 164085 199811 164113
rect 199839 164085 199887 164113
rect 199577 164051 199887 164085
rect 199577 164023 199625 164051
rect 199653 164023 199687 164051
rect 199715 164023 199749 164051
rect 199777 164023 199811 164051
rect 199839 164023 199887 164051
rect 199577 163989 199887 164023
rect 199577 163961 199625 163989
rect 199653 163961 199687 163989
rect 199715 163961 199749 163989
rect 199777 163961 199811 163989
rect 199839 163961 199887 163989
rect 199577 155175 199887 163961
rect 199577 155147 199625 155175
rect 199653 155147 199687 155175
rect 199715 155147 199749 155175
rect 199777 155147 199811 155175
rect 199839 155147 199887 155175
rect 199577 155113 199887 155147
rect 199577 155085 199625 155113
rect 199653 155085 199687 155113
rect 199715 155085 199749 155113
rect 199777 155085 199811 155113
rect 199839 155085 199887 155113
rect 199577 155051 199887 155085
rect 199577 155023 199625 155051
rect 199653 155023 199687 155051
rect 199715 155023 199749 155051
rect 199777 155023 199811 155051
rect 199839 155023 199887 155051
rect 199577 154989 199887 155023
rect 199577 154961 199625 154989
rect 199653 154961 199687 154989
rect 199715 154961 199749 154989
rect 199777 154961 199811 154989
rect 199839 154961 199887 154989
rect 199577 146175 199887 154961
rect 199577 146147 199625 146175
rect 199653 146147 199687 146175
rect 199715 146147 199749 146175
rect 199777 146147 199811 146175
rect 199839 146147 199887 146175
rect 199577 146113 199887 146147
rect 199577 146085 199625 146113
rect 199653 146085 199687 146113
rect 199715 146085 199749 146113
rect 199777 146085 199811 146113
rect 199839 146085 199887 146113
rect 199577 146051 199887 146085
rect 199577 146023 199625 146051
rect 199653 146023 199687 146051
rect 199715 146023 199749 146051
rect 199777 146023 199811 146051
rect 199839 146023 199887 146051
rect 199577 145989 199887 146023
rect 199577 145961 199625 145989
rect 199653 145961 199687 145989
rect 199715 145961 199749 145989
rect 199777 145961 199811 145989
rect 199839 145961 199887 145989
rect 199577 137175 199887 145961
rect 199577 137147 199625 137175
rect 199653 137147 199687 137175
rect 199715 137147 199749 137175
rect 199777 137147 199811 137175
rect 199839 137147 199887 137175
rect 199577 137113 199887 137147
rect 199577 137085 199625 137113
rect 199653 137085 199687 137113
rect 199715 137085 199749 137113
rect 199777 137085 199811 137113
rect 199839 137085 199887 137113
rect 199577 137051 199887 137085
rect 199577 137023 199625 137051
rect 199653 137023 199687 137051
rect 199715 137023 199749 137051
rect 199777 137023 199811 137051
rect 199839 137023 199887 137051
rect 199577 136989 199887 137023
rect 199577 136961 199625 136989
rect 199653 136961 199687 136989
rect 199715 136961 199749 136989
rect 199777 136961 199811 136989
rect 199839 136961 199887 136989
rect 199577 128175 199887 136961
rect 199577 128147 199625 128175
rect 199653 128147 199687 128175
rect 199715 128147 199749 128175
rect 199777 128147 199811 128175
rect 199839 128147 199887 128175
rect 199577 128113 199887 128147
rect 199577 128085 199625 128113
rect 199653 128085 199687 128113
rect 199715 128085 199749 128113
rect 199777 128085 199811 128113
rect 199839 128085 199887 128113
rect 199577 128051 199887 128085
rect 199577 128023 199625 128051
rect 199653 128023 199687 128051
rect 199715 128023 199749 128051
rect 199777 128023 199811 128051
rect 199839 128023 199887 128051
rect 199577 127989 199887 128023
rect 199577 127961 199625 127989
rect 199653 127961 199687 127989
rect 199715 127961 199749 127989
rect 199777 127961 199811 127989
rect 199839 127961 199887 127989
rect 199577 119175 199887 127961
rect 199577 119147 199625 119175
rect 199653 119147 199687 119175
rect 199715 119147 199749 119175
rect 199777 119147 199811 119175
rect 199839 119147 199887 119175
rect 199577 119113 199887 119147
rect 199577 119085 199625 119113
rect 199653 119085 199687 119113
rect 199715 119085 199749 119113
rect 199777 119085 199811 119113
rect 199839 119085 199887 119113
rect 199577 119051 199887 119085
rect 199577 119023 199625 119051
rect 199653 119023 199687 119051
rect 199715 119023 199749 119051
rect 199777 119023 199811 119051
rect 199839 119023 199887 119051
rect 199577 118989 199887 119023
rect 199577 118961 199625 118989
rect 199653 118961 199687 118989
rect 199715 118961 199749 118989
rect 199777 118961 199811 118989
rect 199839 118961 199887 118989
rect 199577 110175 199887 118961
rect 199577 110147 199625 110175
rect 199653 110147 199687 110175
rect 199715 110147 199749 110175
rect 199777 110147 199811 110175
rect 199839 110147 199887 110175
rect 199577 110113 199887 110147
rect 199577 110085 199625 110113
rect 199653 110085 199687 110113
rect 199715 110085 199749 110113
rect 199777 110085 199811 110113
rect 199839 110085 199887 110113
rect 199577 110051 199887 110085
rect 199577 110023 199625 110051
rect 199653 110023 199687 110051
rect 199715 110023 199749 110051
rect 199777 110023 199811 110051
rect 199839 110023 199887 110051
rect 199577 109989 199887 110023
rect 199577 109961 199625 109989
rect 199653 109961 199687 109989
rect 199715 109961 199749 109989
rect 199777 109961 199811 109989
rect 199839 109961 199887 109989
rect 199577 101175 199887 109961
rect 199577 101147 199625 101175
rect 199653 101147 199687 101175
rect 199715 101147 199749 101175
rect 199777 101147 199811 101175
rect 199839 101147 199887 101175
rect 199577 101113 199887 101147
rect 199577 101085 199625 101113
rect 199653 101085 199687 101113
rect 199715 101085 199749 101113
rect 199777 101085 199811 101113
rect 199839 101085 199887 101113
rect 199577 101051 199887 101085
rect 199577 101023 199625 101051
rect 199653 101023 199687 101051
rect 199715 101023 199749 101051
rect 199777 101023 199811 101051
rect 199839 101023 199887 101051
rect 199577 100989 199887 101023
rect 199577 100961 199625 100989
rect 199653 100961 199687 100989
rect 199715 100961 199749 100989
rect 199777 100961 199811 100989
rect 199839 100961 199887 100989
rect 199577 92175 199887 100961
rect 199577 92147 199625 92175
rect 199653 92147 199687 92175
rect 199715 92147 199749 92175
rect 199777 92147 199811 92175
rect 199839 92147 199887 92175
rect 199577 92113 199887 92147
rect 199577 92085 199625 92113
rect 199653 92085 199687 92113
rect 199715 92085 199749 92113
rect 199777 92085 199811 92113
rect 199839 92085 199887 92113
rect 199577 92051 199887 92085
rect 199577 92023 199625 92051
rect 199653 92023 199687 92051
rect 199715 92023 199749 92051
rect 199777 92023 199811 92051
rect 199839 92023 199887 92051
rect 199577 91989 199887 92023
rect 199577 91961 199625 91989
rect 199653 91961 199687 91989
rect 199715 91961 199749 91989
rect 199777 91961 199811 91989
rect 199839 91961 199887 91989
rect 199577 83175 199887 91961
rect 199577 83147 199625 83175
rect 199653 83147 199687 83175
rect 199715 83147 199749 83175
rect 199777 83147 199811 83175
rect 199839 83147 199887 83175
rect 199577 83113 199887 83147
rect 199577 83085 199625 83113
rect 199653 83085 199687 83113
rect 199715 83085 199749 83113
rect 199777 83085 199811 83113
rect 199839 83085 199887 83113
rect 199577 83051 199887 83085
rect 199577 83023 199625 83051
rect 199653 83023 199687 83051
rect 199715 83023 199749 83051
rect 199777 83023 199811 83051
rect 199839 83023 199887 83051
rect 199577 82989 199887 83023
rect 199577 82961 199625 82989
rect 199653 82961 199687 82989
rect 199715 82961 199749 82989
rect 199777 82961 199811 82989
rect 199839 82961 199887 82989
rect 199577 74175 199887 82961
rect 199577 74147 199625 74175
rect 199653 74147 199687 74175
rect 199715 74147 199749 74175
rect 199777 74147 199811 74175
rect 199839 74147 199887 74175
rect 199577 74113 199887 74147
rect 199577 74085 199625 74113
rect 199653 74085 199687 74113
rect 199715 74085 199749 74113
rect 199777 74085 199811 74113
rect 199839 74085 199887 74113
rect 199577 74051 199887 74085
rect 199577 74023 199625 74051
rect 199653 74023 199687 74051
rect 199715 74023 199749 74051
rect 199777 74023 199811 74051
rect 199839 74023 199887 74051
rect 199577 73989 199887 74023
rect 199577 73961 199625 73989
rect 199653 73961 199687 73989
rect 199715 73961 199749 73989
rect 199777 73961 199811 73989
rect 199839 73961 199887 73989
rect 199577 65175 199887 73961
rect 199577 65147 199625 65175
rect 199653 65147 199687 65175
rect 199715 65147 199749 65175
rect 199777 65147 199811 65175
rect 199839 65147 199887 65175
rect 199577 65113 199887 65147
rect 199577 65085 199625 65113
rect 199653 65085 199687 65113
rect 199715 65085 199749 65113
rect 199777 65085 199811 65113
rect 199839 65085 199887 65113
rect 199577 65051 199887 65085
rect 199577 65023 199625 65051
rect 199653 65023 199687 65051
rect 199715 65023 199749 65051
rect 199777 65023 199811 65051
rect 199839 65023 199887 65051
rect 199577 64989 199887 65023
rect 199577 64961 199625 64989
rect 199653 64961 199687 64989
rect 199715 64961 199749 64989
rect 199777 64961 199811 64989
rect 199839 64961 199887 64989
rect 199577 56175 199887 64961
rect 199577 56147 199625 56175
rect 199653 56147 199687 56175
rect 199715 56147 199749 56175
rect 199777 56147 199811 56175
rect 199839 56147 199887 56175
rect 199577 56113 199887 56147
rect 199577 56085 199625 56113
rect 199653 56085 199687 56113
rect 199715 56085 199749 56113
rect 199777 56085 199811 56113
rect 199839 56085 199887 56113
rect 199577 56051 199887 56085
rect 199577 56023 199625 56051
rect 199653 56023 199687 56051
rect 199715 56023 199749 56051
rect 199777 56023 199811 56051
rect 199839 56023 199887 56051
rect 199577 55989 199887 56023
rect 199577 55961 199625 55989
rect 199653 55961 199687 55989
rect 199715 55961 199749 55989
rect 199777 55961 199811 55989
rect 199839 55961 199887 55989
rect 199577 47175 199887 55961
rect 199577 47147 199625 47175
rect 199653 47147 199687 47175
rect 199715 47147 199749 47175
rect 199777 47147 199811 47175
rect 199839 47147 199887 47175
rect 199577 47113 199887 47147
rect 199577 47085 199625 47113
rect 199653 47085 199687 47113
rect 199715 47085 199749 47113
rect 199777 47085 199811 47113
rect 199839 47085 199887 47113
rect 199577 47051 199887 47085
rect 199577 47023 199625 47051
rect 199653 47023 199687 47051
rect 199715 47023 199749 47051
rect 199777 47023 199811 47051
rect 199839 47023 199887 47051
rect 199577 46989 199887 47023
rect 199577 46961 199625 46989
rect 199653 46961 199687 46989
rect 199715 46961 199749 46989
rect 199777 46961 199811 46989
rect 199839 46961 199887 46989
rect 199577 38175 199887 46961
rect 199577 38147 199625 38175
rect 199653 38147 199687 38175
rect 199715 38147 199749 38175
rect 199777 38147 199811 38175
rect 199839 38147 199887 38175
rect 199577 38113 199887 38147
rect 199577 38085 199625 38113
rect 199653 38085 199687 38113
rect 199715 38085 199749 38113
rect 199777 38085 199811 38113
rect 199839 38085 199887 38113
rect 199577 38051 199887 38085
rect 199577 38023 199625 38051
rect 199653 38023 199687 38051
rect 199715 38023 199749 38051
rect 199777 38023 199811 38051
rect 199839 38023 199887 38051
rect 199577 37989 199887 38023
rect 199577 37961 199625 37989
rect 199653 37961 199687 37989
rect 199715 37961 199749 37989
rect 199777 37961 199811 37989
rect 199839 37961 199887 37989
rect 199577 29175 199887 37961
rect 199577 29147 199625 29175
rect 199653 29147 199687 29175
rect 199715 29147 199749 29175
rect 199777 29147 199811 29175
rect 199839 29147 199887 29175
rect 199577 29113 199887 29147
rect 199577 29085 199625 29113
rect 199653 29085 199687 29113
rect 199715 29085 199749 29113
rect 199777 29085 199811 29113
rect 199839 29085 199887 29113
rect 199577 29051 199887 29085
rect 199577 29023 199625 29051
rect 199653 29023 199687 29051
rect 199715 29023 199749 29051
rect 199777 29023 199811 29051
rect 199839 29023 199887 29051
rect 199577 28989 199887 29023
rect 199577 28961 199625 28989
rect 199653 28961 199687 28989
rect 199715 28961 199749 28989
rect 199777 28961 199811 28989
rect 199839 28961 199887 28989
rect 199577 20175 199887 28961
rect 199577 20147 199625 20175
rect 199653 20147 199687 20175
rect 199715 20147 199749 20175
rect 199777 20147 199811 20175
rect 199839 20147 199887 20175
rect 199577 20113 199887 20147
rect 199577 20085 199625 20113
rect 199653 20085 199687 20113
rect 199715 20085 199749 20113
rect 199777 20085 199811 20113
rect 199839 20085 199887 20113
rect 199577 20051 199887 20085
rect 199577 20023 199625 20051
rect 199653 20023 199687 20051
rect 199715 20023 199749 20051
rect 199777 20023 199811 20051
rect 199839 20023 199887 20051
rect 199577 19989 199887 20023
rect 199577 19961 199625 19989
rect 199653 19961 199687 19989
rect 199715 19961 199749 19989
rect 199777 19961 199811 19989
rect 199839 19961 199887 19989
rect 199577 11175 199887 19961
rect 199577 11147 199625 11175
rect 199653 11147 199687 11175
rect 199715 11147 199749 11175
rect 199777 11147 199811 11175
rect 199839 11147 199887 11175
rect 199577 11113 199887 11147
rect 199577 11085 199625 11113
rect 199653 11085 199687 11113
rect 199715 11085 199749 11113
rect 199777 11085 199811 11113
rect 199839 11085 199887 11113
rect 199577 11051 199887 11085
rect 199577 11023 199625 11051
rect 199653 11023 199687 11051
rect 199715 11023 199749 11051
rect 199777 11023 199811 11051
rect 199839 11023 199887 11051
rect 199577 10989 199887 11023
rect 199577 10961 199625 10989
rect 199653 10961 199687 10989
rect 199715 10961 199749 10989
rect 199777 10961 199811 10989
rect 199839 10961 199887 10989
rect 199577 2175 199887 10961
rect 199577 2147 199625 2175
rect 199653 2147 199687 2175
rect 199715 2147 199749 2175
rect 199777 2147 199811 2175
rect 199839 2147 199887 2175
rect 199577 2113 199887 2147
rect 199577 2085 199625 2113
rect 199653 2085 199687 2113
rect 199715 2085 199749 2113
rect 199777 2085 199811 2113
rect 199839 2085 199887 2113
rect 199577 2051 199887 2085
rect 199577 2023 199625 2051
rect 199653 2023 199687 2051
rect 199715 2023 199749 2051
rect 199777 2023 199811 2051
rect 199839 2023 199887 2051
rect 199577 1989 199887 2023
rect 199577 1961 199625 1989
rect 199653 1961 199687 1989
rect 199715 1961 199749 1989
rect 199777 1961 199811 1989
rect 199839 1961 199887 1989
rect 199577 -80 199887 1961
rect 199577 -108 199625 -80
rect 199653 -108 199687 -80
rect 199715 -108 199749 -80
rect 199777 -108 199811 -80
rect 199839 -108 199887 -80
rect 199577 -142 199887 -108
rect 199577 -170 199625 -142
rect 199653 -170 199687 -142
rect 199715 -170 199749 -142
rect 199777 -170 199811 -142
rect 199839 -170 199887 -142
rect 199577 -204 199887 -170
rect 199577 -232 199625 -204
rect 199653 -232 199687 -204
rect 199715 -232 199749 -204
rect 199777 -232 199811 -204
rect 199839 -232 199887 -204
rect 199577 -266 199887 -232
rect 199577 -294 199625 -266
rect 199653 -294 199687 -266
rect 199715 -294 199749 -266
rect 199777 -294 199811 -266
rect 199839 -294 199887 -266
rect 199577 -822 199887 -294
rect 201437 299086 201747 299134
rect 201437 299058 201485 299086
rect 201513 299058 201547 299086
rect 201575 299058 201609 299086
rect 201637 299058 201671 299086
rect 201699 299058 201747 299086
rect 201437 299024 201747 299058
rect 201437 298996 201485 299024
rect 201513 298996 201547 299024
rect 201575 298996 201609 299024
rect 201637 298996 201671 299024
rect 201699 298996 201747 299024
rect 201437 298962 201747 298996
rect 201437 298934 201485 298962
rect 201513 298934 201547 298962
rect 201575 298934 201609 298962
rect 201637 298934 201671 298962
rect 201699 298934 201747 298962
rect 201437 298900 201747 298934
rect 201437 298872 201485 298900
rect 201513 298872 201547 298900
rect 201575 298872 201609 298900
rect 201637 298872 201671 298900
rect 201699 298872 201747 298900
rect 201437 293175 201747 298872
rect 201437 293147 201485 293175
rect 201513 293147 201547 293175
rect 201575 293147 201609 293175
rect 201637 293147 201671 293175
rect 201699 293147 201747 293175
rect 201437 293113 201747 293147
rect 201437 293085 201485 293113
rect 201513 293085 201547 293113
rect 201575 293085 201609 293113
rect 201637 293085 201671 293113
rect 201699 293085 201747 293113
rect 201437 293051 201747 293085
rect 201437 293023 201485 293051
rect 201513 293023 201547 293051
rect 201575 293023 201609 293051
rect 201637 293023 201671 293051
rect 201699 293023 201747 293051
rect 201437 292989 201747 293023
rect 201437 292961 201485 292989
rect 201513 292961 201547 292989
rect 201575 292961 201609 292989
rect 201637 292961 201671 292989
rect 201699 292961 201747 292989
rect 201437 284175 201747 292961
rect 201437 284147 201485 284175
rect 201513 284147 201547 284175
rect 201575 284147 201609 284175
rect 201637 284147 201671 284175
rect 201699 284147 201747 284175
rect 201437 284113 201747 284147
rect 201437 284085 201485 284113
rect 201513 284085 201547 284113
rect 201575 284085 201609 284113
rect 201637 284085 201671 284113
rect 201699 284085 201747 284113
rect 201437 284051 201747 284085
rect 201437 284023 201485 284051
rect 201513 284023 201547 284051
rect 201575 284023 201609 284051
rect 201637 284023 201671 284051
rect 201699 284023 201747 284051
rect 201437 283989 201747 284023
rect 201437 283961 201485 283989
rect 201513 283961 201547 283989
rect 201575 283961 201609 283989
rect 201637 283961 201671 283989
rect 201699 283961 201747 283989
rect 201437 275175 201747 283961
rect 201437 275147 201485 275175
rect 201513 275147 201547 275175
rect 201575 275147 201609 275175
rect 201637 275147 201671 275175
rect 201699 275147 201747 275175
rect 201437 275113 201747 275147
rect 201437 275085 201485 275113
rect 201513 275085 201547 275113
rect 201575 275085 201609 275113
rect 201637 275085 201671 275113
rect 201699 275085 201747 275113
rect 201437 275051 201747 275085
rect 201437 275023 201485 275051
rect 201513 275023 201547 275051
rect 201575 275023 201609 275051
rect 201637 275023 201671 275051
rect 201699 275023 201747 275051
rect 201437 274989 201747 275023
rect 201437 274961 201485 274989
rect 201513 274961 201547 274989
rect 201575 274961 201609 274989
rect 201637 274961 201671 274989
rect 201699 274961 201747 274989
rect 201437 266175 201747 274961
rect 201437 266147 201485 266175
rect 201513 266147 201547 266175
rect 201575 266147 201609 266175
rect 201637 266147 201671 266175
rect 201699 266147 201747 266175
rect 201437 266113 201747 266147
rect 201437 266085 201485 266113
rect 201513 266085 201547 266113
rect 201575 266085 201609 266113
rect 201637 266085 201671 266113
rect 201699 266085 201747 266113
rect 201437 266051 201747 266085
rect 201437 266023 201485 266051
rect 201513 266023 201547 266051
rect 201575 266023 201609 266051
rect 201637 266023 201671 266051
rect 201699 266023 201747 266051
rect 201437 265989 201747 266023
rect 201437 265961 201485 265989
rect 201513 265961 201547 265989
rect 201575 265961 201609 265989
rect 201637 265961 201671 265989
rect 201699 265961 201747 265989
rect 201437 257175 201747 265961
rect 201437 257147 201485 257175
rect 201513 257147 201547 257175
rect 201575 257147 201609 257175
rect 201637 257147 201671 257175
rect 201699 257147 201747 257175
rect 201437 257113 201747 257147
rect 201437 257085 201485 257113
rect 201513 257085 201547 257113
rect 201575 257085 201609 257113
rect 201637 257085 201671 257113
rect 201699 257085 201747 257113
rect 201437 257051 201747 257085
rect 201437 257023 201485 257051
rect 201513 257023 201547 257051
rect 201575 257023 201609 257051
rect 201637 257023 201671 257051
rect 201699 257023 201747 257051
rect 201437 256989 201747 257023
rect 201437 256961 201485 256989
rect 201513 256961 201547 256989
rect 201575 256961 201609 256989
rect 201637 256961 201671 256989
rect 201699 256961 201747 256989
rect 201437 248175 201747 256961
rect 201437 248147 201485 248175
rect 201513 248147 201547 248175
rect 201575 248147 201609 248175
rect 201637 248147 201671 248175
rect 201699 248147 201747 248175
rect 201437 248113 201747 248147
rect 201437 248085 201485 248113
rect 201513 248085 201547 248113
rect 201575 248085 201609 248113
rect 201637 248085 201671 248113
rect 201699 248085 201747 248113
rect 201437 248051 201747 248085
rect 201437 248023 201485 248051
rect 201513 248023 201547 248051
rect 201575 248023 201609 248051
rect 201637 248023 201671 248051
rect 201699 248023 201747 248051
rect 201437 247989 201747 248023
rect 201437 247961 201485 247989
rect 201513 247961 201547 247989
rect 201575 247961 201609 247989
rect 201637 247961 201671 247989
rect 201699 247961 201747 247989
rect 201437 239175 201747 247961
rect 201437 239147 201485 239175
rect 201513 239147 201547 239175
rect 201575 239147 201609 239175
rect 201637 239147 201671 239175
rect 201699 239147 201747 239175
rect 201437 239113 201747 239147
rect 201437 239085 201485 239113
rect 201513 239085 201547 239113
rect 201575 239085 201609 239113
rect 201637 239085 201671 239113
rect 201699 239085 201747 239113
rect 201437 239051 201747 239085
rect 201437 239023 201485 239051
rect 201513 239023 201547 239051
rect 201575 239023 201609 239051
rect 201637 239023 201671 239051
rect 201699 239023 201747 239051
rect 201437 238989 201747 239023
rect 201437 238961 201485 238989
rect 201513 238961 201547 238989
rect 201575 238961 201609 238989
rect 201637 238961 201671 238989
rect 201699 238961 201747 238989
rect 201437 230175 201747 238961
rect 201437 230147 201485 230175
rect 201513 230147 201547 230175
rect 201575 230147 201609 230175
rect 201637 230147 201671 230175
rect 201699 230147 201747 230175
rect 201437 230113 201747 230147
rect 201437 230085 201485 230113
rect 201513 230085 201547 230113
rect 201575 230085 201609 230113
rect 201637 230085 201671 230113
rect 201699 230085 201747 230113
rect 201437 230051 201747 230085
rect 201437 230023 201485 230051
rect 201513 230023 201547 230051
rect 201575 230023 201609 230051
rect 201637 230023 201671 230051
rect 201699 230023 201747 230051
rect 201437 229989 201747 230023
rect 201437 229961 201485 229989
rect 201513 229961 201547 229989
rect 201575 229961 201609 229989
rect 201637 229961 201671 229989
rect 201699 229961 201747 229989
rect 201437 221175 201747 229961
rect 201437 221147 201485 221175
rect 201513 221147 201547 221175
rect 201575 221147 201609 221175
rect 201637 221147 201671 221175
rect 201699 221147 201747 221175
rect 201437 221113 201747 221147
rect 201437 221085 201485 221113
rect 201513 221085 201547 221113
rect 201575 221085 201609 221113
rect 201637 221085 201671 221113
rect 201699 221085 201747 221113
rect 201437 221051 201747 221085
rect 201437 221023 201485 221051
rect 201513 221023 201547 221051
rect 201575 221023 201609 221051
rect 201637 221023 201671 221051
rect 201699 221023 201747 221051
rect 201437 220989 201747 221023
rect 201437 220961 201485 220989
rect 201513 220961 201547 220989
rect 201575 220961 201609 220989
rect 201637 220961 201671 220989
rect 201699 220961 201747 220989
rect 201437 212175 201747 220961
rect 201437 212147 201485 212175
rect 201513 212147 201547 212175
rect 201575 212147 201609 212175
rect 201637 212147 201671 212175
rect 201699 212147 201747 212175
rect 201437 212113 201747 212147
rect 201437 212085 201485 212113
rect 201513 212085 201547 212113
rect 201575 212085 201609 212113
rect 201637 212085 201671 212113
rect 201699 212085 201747 212113
rect 201437 212051 201747 212085
rect 201437 212023 201485 212051
rect 201513 212023 201547 212051
rect 201575 212023 201609 212051
rect 201637 212023 201671 212051
rect 201699 212023 201747 212051
rect 201437 211989 201747 212023
rect 201437 211961 201485 211989
rect 201513 211961 201547 211989
rect 201575 211961 201609 211989
rect 201637 211961 201671 211989
rect 201699 211961 201747 211989
rect 201437 203175 201747 211961
rect 201437 203147 201485 203175
rect 201513 203147 201547 203175
rect 201575 203147 201609 203175
rect 201637 203147 201671 203175
rect 201699 203147 201747 203175
rect 201437 203113 201747 203147
rect 201437 203085 201485 203113
rect 201513 203085 201547 203113
rect 201575 203085 201609 203113
rect 201637 203085 201671 203113
rect 201699 203085 201747 203113
rect 201437 203051 201747 203085
rect 201437 203023 201485 203051
rect 201513 203023 201547 203051
rect 201575 203023 201609 203051
rect 201637 203023 201671 203051
rect 201699 203023 201747 203051
rect 201437 202989 201747 203023
rect 201437 202961 201485 202989
rect 201513 202961 201547 202989
rect 201575 202961 201609 202989
rect 201637 202961 201671 202989
rect 201699 202961 201747 202989
rect 201437 194175 201747 202961
rect 201437 194147 201485 194175
rect 201513 194147 201547 194175
rect 201575 194147 201609 194175
rect 201637 194147 201671 194175
rect 201699 194147 201747 194175
rect 201437 194113 201747 194147
rect 201437 194085 201485 194113
rect 201513 194085 201547 194113
rect 201575 194085 201609 194113
rect 201637 194085 201671 194113
rect 201699 194085 201747 194113
rect 201437 194051 201747 194085
rect 201437 194023 201485 194051
rect 201513 194023 201547 194051
rect 201575 194023 201609 194051
rect 201637 194023 201671 194051
rect 201699 194023 201747 194051
rect 201437 193989 201747 194023
rect 201437 193961 201485 193989
rect 201513 193961 201547 193989
rect 201575 193961 201609 193989
rect 201637 193961 201671 193989
rect 201699 193961 201747 193989
rect 201437 185175 201747 193961
rect 201437 185147 201485 185175
rect 201513 185147 201547 185175
rect 201575 185147 201609 185175
rect 201637 185147 201671 185175
rect 201699 185147 201747 185175
rect 201437 185113 201747 185147
rect 201437 185085 201485 185113
rect 201513 185085 201547 185113
rect 201575 185085 201609 185113
rect 201637 185085 201671 185113
rect 201699 185085 201747 185113
rect 201437 185051 201747 185085
rect 201437 185023 201485 185051
rect 201513 185023 201547 185051
rect 201575 185023 201609 185051
rect 201637 185023 201671 185051
rect 201699 185023 201747 185051
rect 201437 184989 201747 185023
rect 201437 184961 201485 184989
rect 201513 184961 201547 184989
rect 201575 184961 201609 184989
rect 201637 184961 201671 184989
rect 201699 184961 201747 184989
rect 201437 176175 201747 184961
rect 201437 176147 201485 176175
rect 201513 176147 201547 176175
rect 201575 176147 201609 176175
rect 201637 176147 201671 176175
rect 201699 176147 201747 176175
rect 201437 176113 201747 176147
rect 201437 176085 201485 176113
rect 201513 176085 201547 176113
rect 201575 176085 201609 176113
rect 201637 176085 201671 176113
rect 201699 176085 201747 176113
rect 201437 176051 201747 176085
rect 201437 176023 201485 176051
rect 201513 176023 201547 176051
rect 201575 176023 201609 176051
rect 201637 176023 201671 176051
rect 201699 176023 201747 176051
rect 201437 175989 201747 176023
rect 201437 175961 201485 175989
rect 201513 175961 201547 175989
rect 201575 175961 201609 175989
rect 201637 175961 201671 175989
rect 201699 175961 201747 175989
rect 201437 167175 201747 175961
rect 201437 167147 201485 167175
rect 201513 167147 201547 167175
rect 201575 167147 201609 167175
rect 201637 167147 201671 167175
rect 201699 167147 201747 167175
rect 201437 167113 201747 167147
rect 201437 167085 201485 167113
rect 201513 167085 201547 167113
rect 201575 167085 201609 167113
rect 201637 167085 201671 167113
rect 201699 167085 201747 167113
rect 201437 167051 201747 167085
rect 201437 167023 201485 167051
rect 201513 167023 201547 167051
rect 201575 167023 201609 167051
rect 201637 167023 201671 167051
rect 201699 167023 201747 167051
rect 201437 166989 201747 167023
rect 201437 166961 201485 166989
rect 201513 166961 201547 166989
rect 201575 166961 201609 166989
rect 201637 166961 201671 166989
rect 201699 166961 201747 166989
rect 201437 158175 201747 166961
rect 201437 158147 201485 158175
rect 201513 158147 201547 158175
rect 201575 158147 201609 158175
rect 201637 158147 201671 158175
rect 201699 158147 201747 158175
rect 201437 158113 201747 158147
rect 201437 158085 201485 158113
rect 201513 158085 201547 158113
rect 201575 158085 201609 158113
rect 201637 158085 201671 158113
rect 201699 158085 201747 158113
rect 201437 158051 201747 158085
rect 201437 158023 201485 158051
rect 201513 158023 201547 158051
rect 201575 158023 201609 158051
rect 201637 158023 201671 158051
rect 201699 158023 201747 158051
rect 201437 157989 201747 158023
rect 201437 157961 201485 157989
rect 201513 157961 201547 157989
rect 201575 157961 201609 157989
rect 201637 157961 201671 157989
rect 201699 157961 201747 157989
rect 201437 149175 201747 157961
rect 201437 149147 201485 149175
rect 201513 149147 201547 149175
rect 201575 149147 201609 149175
rect 201637 149147 201671 149175
rect 201699 149147 201747 149175
rect 201437 149113 201747 149147
rect 201437 149085 201485 149113
rect 201513 149085 201547 149113
rect 201575 149085 201609 149113
rect 201637 149085 201671 149113
rect 201699 149085 201747 149113
rect 201437 149051 201747 149085
rect 201437 149023 201485 149051
rect 201513 149023 201547 149051
rect 201575 149023 201609 149051
rect 201637 149023 201671 149051
rect 201699 149023 201747 149051
rect 201437 148989 201747 149023
rect 201437 148961 201485 148989
rect 201513 148961 201547 148989
rect 201575 148961 201609 148989
rect 201637 148961 201671 148989
rect 201699 148961 201747 148989
rect 201437 140175 201747 148961
rect 201437 140147 201485 140175
rect 201513 140147 201547 140175
rect 201575 140147 201609 140175
rect 201637 140147 201671 140175
rect 201699 140147 201747 140175
rect 201437 140113 201747 140147
rect 201437 140085 201485 140113
rect 201513 140085 201547 140113
rect 201575 140085 201609 140113
rect 201637 140085 201671 140113
rect 201699 140085 201747 140113
rect 201437 140051 201747 140085
rect 201437 140023 201485 140051
rect 201513 140023 201547 140051
rect 201575 140023 201609 140051
rect 201637 140023 201671 140051
rect 201699 140023 201747 140051
rect 201437 139989 201747 140023
rect 201437 139961 201485 139989
rect 201513 139961 201547 139989
rect 201575 139961 201609 139989
rect 201637 139961 201671 139989
rect 201699 139961 201747 139989
rect 201437 131175 201747 139961
rect 201437 131147 201485 131175
rect 201513 131147 201547 131175
rect 201575 131147 201609 131175
rect 201637 131147 201671 131175
rect 201699 131147 201747 131175
rect 201437 131113 201747 131147
rect 201437 131085 201485 131113
rect 201513 131085 201547 131113
rect 201575 131085 201609 131113
rect 201637 131085 201671 131113
rect 201699 131085 201747 131113
rect 201437 131051 201747 131085
rect 201437 131023 201485 131051
rect 201513 131023 201547 131051
rect 201575 131023 201609 131051
rect 201637 131023 201671 131051
rect 201699 131023 201747 131051
rect 201437 130989 201747 131023
rect 201437 130961 201485 130989
rect 201513 130961 201547 130989
rect 201575 130961 201609 130989
rect 201637 130961 201671 130989
rect 201699 130961 201747 130989
rect 201437 122175 201747 130961
rect 201437 122147 201485 122175
rect 201513 122147 201547 122175
rect 201575 122147 201609 122175
rect 201637 122147 201671 122175
rect 201699 122147 201747 122175
rect 201437 122113 201747 122147
rect 201437 122085 201485 122113
rect 201513 122085 201547 122113
rect 201575 122085 201609 122113
rect 201637 122085 201671 122113
rect 201699 122085 201747 122113
rect 201437 122051 201747 122085
rect 201437 122023 201485 122051
rect 201513 122023 201547 122051
rect 201575 122023 201609 122051
rect 201637 122023 201671 122051
rect 201699 122023 201747 122051
rect 201437 121989 201747 122023
rect 201437 121961 201485 121989
rect 201513 121961 201547 121989
rect 201575 121961 201609 121989
rect 201637 121961 201671 121989
rect 201699 121961 201747 121989
rect 201437 113175 201747 121961
rect 201437 113147 201485 113175
rect 201513 113147 201547 113175
rect 201575 113147 201609 113175
rect 201637 113147 201671 113175
rect 201699 113147 201747 113175
rect 201437 113113 201747 113147
rect 201437 113085 201485 113113
rect 201513 113085 201547 113113
rect 201575 113085 201609 113113
rect 201637 113085 201671 113113
rect 201699 113085 201747 113113
rect 201437 113051 201747 113085
rect 201437 113023 201485 113051
rect 201513 113023 201547 113051
rect 201575 113023 201609 113051
rect 201637 113023 201671 113051
rect 201699 113023 201747 113051
rect 201437 112989 201747 113023
rect 201437 112961 201485 112989
rect 201513 112961 201547 112989
rect 201575 112961 201609 112989
rect 201637 112961 201671 112989
rect 201699 112961 201747 112989
rect 201437 104175 201747 112961
rect 201437 104147 201485 104175
rect 201513 104147 201547 104175
rect 201575 104147 201609 104175
rect 201637 104147 201671 104175
rect 201699 104147 201747 104175
rect 201437 104113 201747 104147
rect 201437 104085 201485 104113
rect 201513 104085 201547 104113
rect 201575 104085 201609 104113
rect 201637 104085 201671 104113
rect 201699 104085 201747 104113
rect 201437 104051 201747 104085
rect 201437 104023 201485 104051
rect 201513 104023 201547 104051
rect 201575 104023 201609 104051
rect 201637 104023 201671 104051
rect 201699 104023 201747 104051
rect 201437 103989 201747 104023
rect 201437 103961 201485 103989
rect 201513 103961 201547 103989
rect 201575 103961 201609 103989
rect 201637 103961 201671 103989
rect 201699 103961 201747 103989
rect 201437 95175 201747 103961
rect 201437 95147 201485 95175
rect 201513 95147 201547 95175
rect 201575 95147 201609 95175
rect 201637 95147 201671 95175
rect 201699 95147 201747 95175
rect 201437 95113 201747 95147
rect 201437 95085 201485 95113
rect 201513 95085 201547 95113
rect 201575 95085 201609 95113
rect 201637 95085 201671 95113
rect 201699 95085 201747 95113
rect 201437 95051 201747 95085
rect 201437 95023 201485 95051
rect 201513 95023 201547 95051
rect 201575 95023 201609 95051
rect 201637 95023 201671 95051
rect 201699 95023 201747 95051
rect 201437 94989 201747 95023
rect 201437 94961 201485 94989
rect 201513 94961 201547 94989
rect 201575 94961 201609 94989
rect 201637 94961 201671 94989
rect 201699 94961 201747 94989
rect 201437 86175 201747 94961
rect 201437 86147 201485 86175
rect 201513 86147 201547 86175
rect 201575 86147 201609 86175
rect 201637 86147 201671 86175
rect 201699 86147 201747 86175
rect 201437 86113 201747 86147
rect 201437 86085 201485 86113
rect 201513 86085 201547 86113
rect 201575 86085 201609 86113
rect 201637 86085 201671 86113
rect 201699 86085 201747 86113
rect 201437 86051 201747 86085
rect 201437 86023 201485 86051
rect 201513 86023 201547 86051
rect 201575 86023 201609 86051
rect 201637 86023 201671 86051
rect 201699 86023 201747 86051
rect 201437 85989 201747 86023
rect 201437 85961 201485 85989
rect 201513 85961 201547 85989
rect 201575 85961 201609 85989
rect 201637 85961 201671 85989
rect 201699 85961 201747 85989
rect 201437 77175 201747 85961
rect 201437 77147 201485 77175
rect 201513 77147 201547 77175
rect 201575 77147 201609 77175
rect 201637 77147 201671 77175
rect 201699 77147 201747 77175
rect 201437 77113 201747 77147
rect 201437 77085 201485 77113
rect 201513 77085 201547 77113
rect 201575 77085 201609 77113
rect 201637 77085 201671 77113
rect 201699 77085 201747 77113
rect 201437 77051 201747 77085
rect 201437 77023 201485 77051
rect 201513 77023 201547 77051
rect 201575 77023 201609 77051
rect 201637 77023 201671 77051
rect 201699 77023 201747 77051
rect 201437 76989 201747 77023
rect 201437 76961 201485 76989
rect 201513 76961 201547 76989
rect 201575 76961 201609 76989
rect 201637 76961 201671 76989
rect 201699 76961 201747 76989
rect 201437 68175 201747 76961
rect 201437 68147 201485 68175
rect 201513 68147 201547 68175
rect 201575 68147 201609 68175
rect 201637 68147 201671 68175
rect 201699 68147 201747 68175
rect 201437 68113 201747 68147
rect 201437 68085 201485 68113
rect 201513 68085 201547 68113
rect 201575 68085 201609 68113
rect 201637 68085 201671 68113
rect 201699 68085 201747 68113
rect 201437 68051 201747 68085
rect 201437 68023 201485 68051
rect 201513 68023 201547 68051
rect 201575 68023 201609 68051
rect 201637 68023 201671 68051
rect 201699 68023 201747 68051
rect 201437 67989 201747 68023
rect 201437 67961 201485 67989
rect 201513 67961 201547 67989
rect 201575 67961 201609 67989
rect 201637 67961 201671 67989
rect 201699 67961 201747 67989
rect 201437 59175 201747 67961
rect 201437 59147 201485 59175
rect 201513 59147 201547 59175
rect 201575 59147 201609 59175
rect 201637 59147 201671 59175
rect 201699 59147 201747 59175
rect 201437 59113 201747 59147
rect 201437 59085 201485 59113
rect 201513 59085 201547 59113
rect 201575 59085 201609 59113
rect 201637 59085 201671 59113
rect 201699 59085 201747 59113
rect 201437 59051 201747 59085
rect 201437 59023 201485 59051
rect 201513 59023 201547 59051
rect 201575 59023 201609 59051
rect 201637 59023 201671 59051
rect 201699 59023 201747 59051
rect 201437 58989 201747 59023
rect 201437 58961 201485 58989
rect 201513 58961 201547 58989
rect 201575 58961 201609 58989
rect 201637 58961 201671 58989
rect 201699 58961 201747 58989
rect 201437 50175 201747 58961
rect 201437 50147 201485 50175
rect 201513 50147 201547 50175
rect 201575 50147 201609 50175
rect 201637 50147 201671 50175
rect 201699 50147 201747 50175
rect 201437 50113 201747 50147
rect 201437 50085 201485 50113
rect 201513 50085 201547 50113
rect 201575 50085 201609 50113
rect 201637 50085 201671 50113
rect 201699 50085 201747 50113
rect 201437 50051 201747 50085
rect 201437 50023 201485 50051
rect 201513 50023 201547 50051
rect 201575 50023 201609 50051
rect 201637 50023 201671 50051
rect 201699 50023 201747 50051
rect 201437 49989 201747 50023
rect 201437 49961 201485 49989
rect 201513 49961 201547 49989
rect 201575 49961 201609 49989
rect 201637 49961 201671 49989
rect 201699 49961 201747 49989
rect 201437 41175 201747 49961
rect 201437 41147 201485 41175
rect 201513 41147 201547 41175
rect 201575 41147 201609 41175
rect 201637 41147 201671 41175
rect 201699 41147 201747 41175
rect 201437 41113 201747 41147
rect 201437 41085 201485 41113
rect 201513 41085 201547 41113
rect 201575 41085 201609 41113
rect 201637 41085 201671 41113
rect 201699 41085 201747 41113
rect 201437 41051 201747 41085
rect 201437 41023 201485 41051
rect 201513 41023 201547 41051
rect 201575 41023 201609 41051
rect 201637 41023 201671 41051
rect 201699 41023 201747 41051
rect 201437 40989 201747 41023
rect 201437 40961 201485 40989
rect 201513 40961 201547 40989
rect 201575 40961 201609 40989
rect 201637 40961 201671 40989
rect 201699 40961 201747 40989
rect 201437 32175 201747 40961
rect 201437 32147 201485 32175
rect 201513 32147 201547 32175
rect 201575 32147 201609 32175
rect 201637 32147 201671 32175
rect 201699 32147 201747 32175
rect 201437 32113 201747 32147
rect 201437 32085 201485 32113
rect 201513 32085 201547 32113
rect 201575 32085 201609 32113
rect 201637 32085 201671 32113
rect 201699 32085 201747 32113
rect 201437 32051 201747 32085
rect 201437 32023 201485 32051
rect 201513 32023 201547 32051
rect 201575 32023 201609 32051
rect 201637 32023 201671 32051
rect 201699 32023 201747 32051
rect 201437 31989 201747 32023
rect 201437 31961 201485 31989
rect 201513 31961 201547 31989
rect 201575 31961 201609 31989
rect 201637 31961 201671 31989
rect 201699 31961 201747 31989
rect 201437 23175 201747 31961
rect 201437 23147 201485 23175
rect 201513 23147 201547 23175
rect 201575 23147 201609 23175
rect 201637 23147 201671 23175
rect 201699 23147 201747 23175
rect 201437 23113 201747 23147
rect 201437 23085 201485 23113
rect 201513 23085 201547 23113
rect 201575 23085 201609 23113
rect 201637 23085 201671 23113
rect 201699 23085 201747 23113
rect 201437 23051 201747 23085
rect 201437 23023 201485 23051
rect 201513 23023 201547 23051
rect 201575 23023 201609 23051
rect 201637 23023 201671 23051
rect 201699 23023 201747 23051
rect 201437 22989 201747 23023
rect 201437 22961 201485 22989
rect 201513 22961 201547 22989
rect 201575 22961 201609 22989
rect 201637 22961 201671 22989
rect 201699 22961 201747 22989
rect 201437 14175 201747 22961
rect 201437 14147 201485 14175
rect 201513 14147 201547 14175
rect 201575 14147 201609 14175
rect 201637 14147 201671 14175
rect 201699 14147 201747 14175
rect 201437 14113 201747 14147
rect 201437 14085 201485 14113
rect 201513 14085 201547 14113
rect 201575 14085 201609 14113
rect 201637 14085 201671 14113
rect 201699 14085 201747 14113
rect 201437 14051 201747 14085
rect 201437 14023 201485 14051
rect 201513 14023 201547 14051
rect 201575 14023 201609 14051
rect 201637 14023 201671 14051
rect 201699 14023 201747 14051
rect 201437 13989 201747 14023
rect 201437 13961 201485 13989
rect 201513 13961 201547 13989
rect 201575 13961 201609 13989
rect 201637 13961 201671 13989
rect 201699 13961 201747 13989
rect 201437 5175 201747 13961
rect 201437 5147 201485 5175
rect 201513 5147 201547 5175
rect 201575 5147 201609 5175
rect 201637 5147 201671 5175
rect 201699 5147 201747 5175
rect 201437 5113 201747 5147
rect 201437 5085 201485 5113
rect 201513 5085 201547 5113
rect 201575 5085 201609 5113
rect 201637 5085 201671 5113
rect 201699 5085 201747 5113
rect 201437 5051 201747 5085
rect 201437 5023 201485 5051
rect 201513 5023 201547 5051
rect 201575 5023 201609 5051
rect 201637 5023 201671 5051
rect 201699 5023 201747 5051
rect 201437 4989 201747 5023
rect 201437 4961 201485 4989
rect 201513 4961 201547 4989
rect 201575 4961 201609 4989
rect 201637 4961 201671 4989
rect 201699 4961 201747 4989
rect 201437 -560 201747 4961
rect 201437 -588 201485 -560
rect 201513 -588 201547 -560
rect 201575 -588 201609 -560
rect 201637 -588 201671 -560
rect 201699 -588 201747 -560
rect 201437 -622 201747 -588
rect 201437 -650 201485 -622
rect 201513 -650 201547 -622
rect 201575 -650 201609 -622
rect 201637 -650 201671 -622
rect 201699 -650 201747 -622
rect 201437 -684 201747 -650
rect 201437 -712 201485 -684
rect 201513 -712 201547 -684
rect 201575 -712 201609 -684
rect 201637 -712 201671 -684
rect 201699 -712 201747 -684
rect 201437 -746 201747 -712
rect 201437 -774 201485 -746
rect 201513 -774 201547 -746
rect 201575 -774 201609 -746
rect 201637 -774 201671 -746
rect 201699 -774 201747 -746
rect 201437 -822 201747 -774
rect 208577 298606 208887 299134
rect 208577 298578 208625 298606
rect 208653 298578 208687 298606
rect 208715 298578 208749 298606
rect 208777 298578 208811 298606
rect 208839 298578 208887 298606
rect 208577 298544 208887 298578
rect 208577 298516 208625 298544
rect 208653 298516 208687 298544
rect 208715 298516 208749 298544
rect 208777 298516 208811 298544
rect 208839 298516 208887 298544
rect 208577 298482 208887 298516
rect 208577 298454 208625 298482
rect 208653 298454 208687 298482
rect 208715 298454 208749 298482
rect 208777 298454 208811 298482
rect 208839 298454 208887 298482
rect 208577 298420 208887 298454
rect 208577 298392 208625 298420
rect 208653 298392 208687 298420
rect 208715 298392 208749 298420
rect 208777 298392 208811 298420
rect 208839 298392 208887 298420
rect 208577 290175 208887 298392
rect 208577 290147 208625 290175
rect 208653 290147 208687 290175
rect 208715 290147 208749 290175
rect 208777 290147 208811 290175
rect 208839 290147 208887 290175
rect 208577 290113 208887 290147
rect 208577 290085 208625 290113
rect 208653 290085 208687 290113
rect 208715 290085 208749 290113
rect 208777 290085 208811 290113
rect 208839 290085 208887 290113
rect 208577 290051 208887 290085
rect 208577 290023 208625 290051
rect 208653 290023 208687 290051
rect 208715 290023 208749 290051
rect 208777 290023 208811 290051
rect 208839 290023 208887 290051
rect 208577 289989 208887 290023
rect 208577 289961 208625 289989
rect 208653 289961 208687 289989
rect 208715 289961 208749 289989
rect 208777 289961 208811 289989
rect 208839 289961 208887 289989
rect 208577 281175 208887 289961
rect 208577 281147 208625 281175
rect 208653 281147 208687 281175
rect 208715 281147 208749 281175
rect 208777 281147 208811 281175
rect 208839 281147 208887 281175
rect 208577 281113 208887 281147
rect 208577 281085 208625 281113
rect 208653 281085 208687 281113
rect 208715 281085 208749 281113
rect 208777 281085 208811 281113
rect 208839 281085 208887 281113
rect 208577 281051 208887 281085
rect 208577 281023 208625 281051
rect 208653 281023 208687 281051
rect 208715 281023 208749 281051
rect 208777 281023 208811 281051
rect 208839 281023 208887 281051
rect 208577 280989 208887 281023
rect 208577 280961 208625 280989
rect 208653 280961 208687 280989
rect 208715 280961 208749 280989
rect 208777 280961 208811 280989
rect 208839 280961 208887 280989
rect 208577 272175 208887 280961
rect 208577 272147 208625 272175
rect 208653 272147 208687 272175
rect 208715 272147 208749 272175
rect 208777 272147 208811 272175
rect 208839 272147 208887 272175
rect 208577 272113 208887 272147
rect 208577 272085 208625 272113
rect 208653 272085 208687 272113
rect 208715 272085 208749 272113
rect 208777 272085 208811 272113
rect 208839 272085 208887 272113
rect 208577 272051 208887 272085
rect 208577 272023 208625 272051
rect 208653 272023 208687 272051
rect 208715 272023 208749 272051
rect 208777 272023 208811 272051
rect 208839 272023 208887 272051
rect 208577 271989 208887 272023
rect 208577 271961 208625 271989
rect 208653 271961 208687 271989
rect 208715 271961 208749 271989
rect 208777 271961 208811 271989
rect 208839 271961 208887 271989
rect 208577 263175 208887 271961
rect 208577 263147 208625 263175
rect 208653 263147 208687 263175
rect 208715 263147 208749 263175
rect 208777 263147 208811 263175
rect 208839 263147 208887 263175
rect 208577 263113 208887 263147
rect 208577 263085 208625 263113
rect 208653 263085 208687 263113
rect 208715 263085 208749 263113
rect 208777 263085 208811 263113
rect 208839 263085 208887 263113
rect 208577 263051 208887 263085
rect 208577 263023 208625 263051
rect 208653 263023 208687 263051
rect 208715 263023 208749 263051
rect 208777 263023 208811 263051
rect 208839 263023 208887 263051
rect 208577 262989 208887 263023
rect 208577 262961 208625 262989
rect 208653 262961 208687 262989
rect 208715 262961 208749 262989
rect 208777 262961 208811 262989
rect 208839 262961 208887 262989
rect 208577 254175 208887 262961
rect 208577 254147 208625 254175
rect 208653 254147 208687 254175
rect 208715 254147 208749 254175
rect 208777 254147 208811 254175
rect 208839 254147 208887 254175
rect 208577 254113 208887 254147
rect 208577 254085 208625 254113
rect 208653 254085 208687 254113
rect 208715 254085 208749 254113
rect 208777 254085 208811 254113
rect 208839 254085 208887 254113
rect 208577 254051 208887 254085
rect 208577 254023 208625 254051
rect 208653 254023 208687 254051
rect 208715 254023 208749 254051
rect 208777 254023 208811 254051
rect 208839 254023 208887 254051
rect 208577 253989 208887 254023
rect 208577 253961 208625 253989
rect 208653 253961 208687 253989
rect 208715 253961 208749 253989
rect 208777 253961 208811 253989
rect 208839 253961 208887 253989
rect 208577 245175 208887 253961
rect 208577 245147 208625 245175
rect 208653 245147 208687 245175
rect 208715 245147 208749 245175
rect 208777 245147 208811 245175
rect 208839 245147 208887 245175
rect 208577 245113 208887 245147
rect 208577 245085 208625 245113
rect 208653 245085 208687 245113
rect 208715 245085 208749 245113
rect 208777 245085 208811 245113
rect 208839 245085 208887 245113
rect 208577 245051 208887 245085
rect 208577 245023 208625 245051
rect 208653 245023 208687 245051
rect 208715 245023 208749 245051
rect 208777 245023 208811 245051
rect 208839 245023 208887 245051
rect 208577 244989 208887 245023
rect 208577 244961 208625 244989
rect 208653 244961 208687 244989
rect 208715 244961 208749 244989
rect 208777 244961 208811 244989
rect 208839 244961 208887 244989
rect 208577 236175 208887 244961
rect 208577 236147 208625 236175
rect 208653 236147 208687 236175
rect 208715 236147 208749 236175
rect 208777 236147 208811 236175
rect 208839 236147 208887 236175
rect 208577 236113 208887 236147
rect 208577 236085 208625 236113
rect 208653 236085 208687 236113
rect 208715 236085 208749 236113
rect 208777 236085 208811 236113
rect 208839 236085 208887 236113
rect 208577 236051 208887 236085
rect 208577 236023 208625 236051
rect 208653 236023 208687 236051
rect 208715 236023 208749 236051
rect 208777 236023 208811 236051
rect 208839 236023 208887 236051
rect 208577 235989 208887 236023
rect 208577 235961 208625 235989
rect 208653 235961 208687 235989
rect 208715 235961 208749 235989
rect 208777 235961 208811 235989
rect 208839 235961 208887 235989
rect 208577 227175 208887 235961
rect 208577 227147 208625 227175
rect 208653 227147 208687 227175
rect 208715 227147 208749 227175
rect 208777 227147 208811 227175
rect 208839 227147 208887 227175
rect 208577 227113 208887 227147
rect 208577 227085 208625 227113
rect 208653 227085 208687 227113
rect 208715 227085 208749 227113
rect 208777 227085 208811 227113
rect 208839 227085 208887 227113
rect 208577 227051 208887 227085
rect 208577 227023 208625 227051
rect 208653 227023 208687 227051
rect 208715 227023 208749 227051
rect 208777 227023 208811 227051
rect 208839 227023 208887 227051
rect 208577 226989 208887 227023
rect 208577 226961 208625 226989
rect 208653 226961 208687 226989
rect 208715 226961 208749 226989
rect 208777 226961 208811 226989
rect 208839 226961 208887 226989
rect 208577 218175 208887 226961
rect 208577 218147 208625 218175
rect 208653 218147 208687 218175
rect 208715 218147 208749 218175
rect 208777 218147 208811 218175
rect 208839 218147 208887 218175
rect 208577 218113 208887 218147
rect 208577 218085 208625 218113
rect 208653 218085 208687 218113
rect 208715 218085 208749 218113
rect 208777 218085 208811 218113
rect 208839 218085 208887 218113
rect 208577 218051 208887 218085
rect 208577 218023 208625 218051
rect 208653 218023 208687 218051
rect 208715 218023 208749 218051
rect 208777 218023 208811 218051
rect 208839 218023 208887 218051
rect 208577 217989 208887 218023
rect 208577 217961 208625 217989
rect 208653 217961 208687 217989
rect 208715 217961 208749 217989
rect 208777 217961 208811 217989
rect 208839 217961 208887 217989
rect 208577 209175 208887 217961
rect 208577 209147 208625 209175
rect 208653 209147 208687 209175
rect 208715 209147 208749 209175
rect 208777 209147 208811 209175
rect 208839 209147 208887 209175
rect 208577 209113 208887 209147
rect 208577 209085 208625 209113
rect 208653 209085 208687 209113
rect 208715 209085 208749 209113
rect 208777 209085 208811 209113
rect 208839 209085 208887 209113
rect 208577 209051 208887 209085
rect 208577 209023 208625 209051
rect 208653 209023 208687 209051
rect 208715 209023 208749 209051
rect 208777 209023 208811 209051
rect 208839 209023 208887 209051
rect 208577 208989 208887 209023
rect 208577 208961 208625 208989
rect 208653 208961 208687 208989
rect 208715 208961 208749 208989
rect 208777 208961 208811 208989
rect 208839 208961 208887 208989
rect 208577 200175 208887 208961
rect 208577 200147 208625 200175
rect 208653 200147 208687 200175
rect 208715 200147 208749 200175
rect 208777 200147 208811 200175
rect 208839 200147 208887 200175
rect 208577 200113 208887 200147
rect 208577 200085 208625 200113
rect 208653 200085 208687 200113
rect 208715 200085 208749 200113
rect 208777 200085 208811 200113
rect 208839 200085 208887 200113
rect 208577 200051 208887 200085
rect 208577 200023 208625 200051
rect 208653 200023 208687 200051
rect 208715 200023 208749 200051
rect 208777 200023 208811 200051
rect 208839 200023 208887 200051
rect 208577 199989 208887 200023
rect 208577 199961 208625 199989
rect 208653 199961 208687 199989
rect 208715 199961 208749 199989
rect 208777 199961 208811 199989
rect 208839 199961 208887 199989
rect 208577 191175 208887 199961
rect 208577 191147 208625 191175
rect 208653 191147 208687 191175
rect 208715 191147 208749 191175
rect 208777 191147 208811 191175
rect 208839 191147 208887 191175
rect 208577 191113 208887 191147
rect 208577 191085 208625 191113
rect 208653 191085 208687 191113
rect 208715 191085 208749 191113
rect 208777 191085 208811 191113
rect 208839 191085 208887 191113
rect 208577 191051 208887 191085
rect 208577 191023 208625 191051
rect 208653 191023 208687 191051
rect 208715 191023 208749 191051
rect 208777 191023 208811 191051
rect 208839 191023 208887 191051
rect 208577 190989 208887 191023
rect 208577 190961 208625 190989
rect 208653 190961 208687 190989
rect 208715 190961 208749 190989
rect 208777 190961 208811 190989
rect 208839 190961 208887 190989
rect 208577 182175 208887 190961
rect 208577 182147 208625 182175
rect 208653 182147 208687 182175
rect 208715 182147 208749 182175
rect 208777 182147 208811 182175
rect 208839 182147 208887 182175
rect 208577 182113 208887 182147
rect 208577 182085 208625 182113
rect 208653 182085 208687 182113
rect 208715 182085 208749 182113
rect 208777 182085 208811 182113
rect 208839 182085 208887 182113
rect 208577 182051 208887 182085
rect 208577 182023 208625 182051
rect 208653 182023 208687 182051
rect 208715 182023 208749 182051
rect 208777 182023 208811 182051
rect 208839 182023 208887 182051
rect 208577 181989 208887 182023
rect 208577 181961 208625 181989
rect 208653 181961 208687 181989
rect 208715 181961 208749 181989
rect 208777 181961 208811 181989
rect 208839 181961 208887 181989
rect 208577 173175 208887 181961
rect 208577 173147 208625 173175
rect 208653 173147 208687 173175
rect 208715 173147 208749 173175
rect 208777 173147 208811 173175
rect 208839 173147 208887 173175
rect 208577 173113 208887 173147
rect 208577 173085 208625 173113
rect 208653 173085 208687 173113
rect 208715 173085 208749 173113
rect 208777 173085 208811 173113
rect 208839 173085 208887 173113
rect 208577 173051 208887 173085
rect 208577 173023 208625 173051
rect 208653 173023 208687 173051
rect 208715 173023 208749 173051
rect 208777 173023 208811 173051
rect 208839 173023 208887 173051
rect 208577 172989 208887 173023
rect 208577 172961 208625 172989
rect 208653 172961 208687 172989
rect 208715 172961 208749 172989
rect 208777 172961 208811 172989
rect 208839 172961 208887 172989
rect 208577 164175 208887 172961
rect 208577 164147 208625 164175
rect 208653 164147 208687 164175
rect 208715 164147 208749 164175
rect 208777 164147 208811 164175
rect 208839 164147 208887 164175
rect 208577 164113 208887 164147
rect 208577 164085 208625 164113
rect 208653 164085 208687 164113
rect 208715 164085 208749 164113
rect 208777 164085 208811 164113
rect 208839 164085 208887 164113
rect 208577 164051 208887 164085
rect 208577 164023 208625 164051
rect 208653 164023 208687 164051
rect 208715 164023 208749 164051
rect 208777 164023 208811 164051
rect 208839 164023 208887 164051
rect 208577 163989 208887 164023
rect 208577 163961 208625 163989
rect 208653 163961 208687 163989
rect 208715 163961 208749 163989
rect 208777 163961 208811 163989
rect 208839 163961 208887 163989
rect 208577 155175 208887 163961
rect 208577 155147 208625 155175
rect 208653 155147 208687 155175
rect 208715 155147 208749 155175
rect 208777 155147 208811 155175
rect 208839 155147 208887 155175
rect 208577 155113 208887 155147
rect 208577 155085 208625 155113
rect 208653 155085 208687 155113
rect 208715 155085 208749 155113
rect 208777 155085 208811 155113
rect 208839 155085 208887 155113
rect 208577 155051 208887 155085
rect 208577 155023 208625 155051
rect 208653 155023 208687 155051
rect 208715 155023 208749 155051
rect 208777 155023 208811 155051
rect 208839 155023 208887 155051
rect 208577 154989 208887 155023
rect 208577 154961 208625 154989
rect 208653 154961 208687 154989
rect 208715 154961 208749 154989
rect 208777 154961 208811 154989
rect 208839 154961 208887 154989
rect 208577 146175 208887 154961
rect 208577 146147 208625 146175
rect 208653 146147 208687 146175
rect 208715 146147 208749 146175
rect 208777 146147 208811 146175
rect 208839 146147 208887 146175
rect 208577 146113 208887 146147
rect 208577 146085 208625 146113
rect 208653 146085 208687 146113
rect 208715 146085 208749 146113
rect 208777 146085 208811 146113
rect 208839 146085 208887 146113
rect 208577 146051 208887 146085
rect 208577 146023 208625 146051
rect 208653 146023 208687 146051
rect 208715 146023 208749 146051
rect 208777 146023 208811 146051
rect 208839 146023 208887 146051
rect 208577 145989 208887 146023
rect 208577 145961 208625 145989
rect 208653 145961 208687 145989
rect 208715 145961 208749 145989
rect 208777 145961 208811 145989
rect 208839 145961 208887 145989
rect 208577 137175 208887 145961
rect 208577 137147 208625 137175
rect 208653 137147 208687 137175
rect 208715 137147 208749 137175
rect 208777 137147 208811 137175
rect 208839 137147 208887 137175
rect 208577 137113 208887 137147
rect 208577 137085 208625 137113
rect 208653 137085 208687 137113
rect 208715 137085 208749 137113
rect 208777 137085 208811 137113
rect 208839 137085 208887 137113
rect 208577 137051 208887 137085
rect 208577 137023 208625 137051
rect 208653 137023 208687 137051
rect 208715 137023 208749 137051
rect 208777 137023 208811 137051
rect 208839 137023 208887 137051
rect 208577 136989 208887 137023
rect 208577 136961 208625 136989
rect 208653 136961 208687 136989
rect 208715 136961 208749 136989
rect 208777 136961 208811 136989
rect 208839 136961 208887 136989
rect 208577 128175 208887 136961
rect 208577 128147 208625 128175
rect 208653 128147 208687 128175
rect 208715 128147 208749 128175
rect 208777 128147 208811 128175
rect 208839 128147 208887 128175
rect 208577 128113 208887 128147
rect 208577 128085 208625 128113
rect 208653 128085 208687 128113
rect 208715 128085 208749 128113
rect 208777 128085 208811 128113
rect 208839 128085 208887 128113
rect 208577 128051 208887 128085
rect 208577 128023 208625 128051
rect 208653 128023 208687 128051
rect 208715 128023 208749 128051
rect 208777 128023 208811 128051
rect 208839 128023 208887 128051
rect 208577 127989 208887 128023
rect 208577 127961 208625 127989
rect 208653 127961 208687 127989
rect 208715 127961 208749 127989
rect 208777 127961 208811 127989
rect 208839 127961 208887 127989
rect 208577 119175 208887 127961
rect 208577 119147 208625 119175
rect 208653 119147 208687 119175
rect 208715 119147 208749 119175
rect 208777 119147 208811 119175
rect 208839 119147 208887 119175
rect 208577 119113 208887 119147
rect 208577 119085 208625 119113
rect 208653 119085 208687 119113
rect 208715 119085 208749 119113
rect 208777 119085 208811 119113
rect 208839 119085 208887 119113
rect 208577 119051 208887 119085
rect 208577 119023 208625 119051
rect 208653 119023 208687 119051
rect 208715 119023 208749 119051
rect 208777 119023 208811 119051
rect 208839 119023 208887 119051
rect 208577 118989 208887 119023
rect 208577 118961 208625 118989
rect 208653 118961 208687 118989
rect 208715 118961 208749 118989
rect 208777 118961 208811 118989
rect 208839 118961 208887 118989
rect 208577 110175 208887 118961
rect 208577 110147 208625 110175
rect 208653 110147 208687 110175
rect 208715 110147 208749 110175
rect 208777 110147 208811 110175
rect 208839 110147 208887 110175
rect 208577 110113 208887 110147
rect 208577 110085 208625 110113
rect 208653 110085 208687 110113
rect 208715 110085 208749 110113
rect 208777 110085 208811 110113
rect 208839 110085 208887 110113
rect 208577 110051 208887 110085
rect 208577 110023 208625 110051
rect 208653 110023 208687 110051
rect 208715 110023 208749 110051
rect 208777 110023 208811 110051
rect 208839 110023 208887 110051
rect 208577 109989 208887 110023
rect 208577 109961 208625 109989
rect 208653 109961 208687 109989
rect 208715 109961 208749 109989
rect 208777 109961 208811 109989
rect 208839 109961 208887 109989
rect 208577 101175 208887 109961
rect 208577 101147 208625 101175
rect 208653 101147 208687 101175
rect 208715 101147 208749 101175
rect 208777 101147 208811 101175
rect 208839 101147 208887 101175
rect 208577 101113 208887 101147
rect 208577 101085 208625 101113
rect 208653 101085 208687 101113
rect 208715 101085 208749 101113
rect 208777 101085 208811 101113
rect 208839 101085 208887 101113
rect 208577 101051 208887 101085
rect 208577 101023 208625 101051
rect 208653 101023 208687 101051
rect 208715 101023 208749 101051
rect 208777 101023 208811 101051
rect 208839 101023 208887 101051
rect 208577 100989 208887 101023
rect 208577 100961 208625 100989
rect 208653 100961 208687 100989
rect 208715 100961 208749 100989
rect 208777 100961 208811 100989
rect 208839 100961 208887 100989
rect 208577 92175 208887 100961
rect 208577 92147 208625 92175
rect 208653 92147 208687 92175
rect 208715 92147 208749 92175
rect 208777 92147 208811 92175
rect 208839 92147 208887 92175
rect 208577 92113 208887 92147
rect 208577 92085 208625 92113
rect 208653 92085 208687 92113
rect 208715 92085 208749 92113
rect 208777 92085 208811 92113
rect 208839 92085 208887 92113
rect 208577 92051 208887 92085
rect 208577 92023 208625 92051
rect 208653 92023 208687 92051
rect 208715 92023 208749 92051
rect 208777 92023 208811 92051
rect 208839 92023 208887 92051
rect 208577 91989 208887 92023
rect 208577 91961 208625 91989
rect 208653 91961 208687 91989
rect 208715 91961 208749 91989
rect 208777 91961 208811 91989
rect 208839 91961 208887 91989
rect 208577 83175 208887 91961
rect 208577 83147 208625 83175
rect 208653 83147 208687 83175
rect 208715 83147 208749 83175
rect 208777 83147 208811 83175
rect 208839 83147 208887 83175
rect 208577 83113 208887 83147
rect 208577 83085 208625 83113
rect 208653 83085 208687 83113
rect 208715 83085 208749 83113
rect 208777 83085 208811 83113
rect 208839 83085 208887 83113
rect 208577 83051 208887 83085
rect 208577 83023 208625 83051
rect 208653 83023 208687 83051
rect 208715 83023 208749 83051
rect 208777 83023 208811 83051
rect 208839 83023 208887 83051
rect 208577 82989 208887 83023
rect 208577 82961 208625 82989
rect 208653 82961 208687 82989
rect 208715 82961 208749 82989
rect 208777 82961 208811 82989
rect 208839 82961 208887 82989
rect 208577 74175 208887 82961
rect 208577 74147 208625 74175
rect 208653 74147 208687 74175
rect 208715 74147 208749 74175
rect 208777 74147 208811 74175
rect 208839 74147 208887 74175
rect 208577 74113 208887 74147
rect 208577 74085 208625 74113
rect 208653 74085 208687 74113
rect 208715 74085 208749 74113
rect 208777 74085 208811 74113
rect 208839 74085 208887 74113
rect 208577 74051 208887 74085
rect 208577 74023 208625 74051
rect 208653 74023 208687 74051
rect 208715 74023 208749 74051
rect 208777 74023 208811 74051
rect 208839 74023 208887 74051
rect 208577 73989 208887 74023
rect 208577 73961 208625 73989
rect 208653 73961 208687 73989
rect 208715 73961 208749 73989
rect 208777 73961 208811 73989
rect 208839 73961 208887 73989
rect 208577 65175 208887 73961
rect 208577 65147 208625 65175
rect 208653 65147 208687 65175
rect 208715 65147 208749 65175
rect 208777 65147 208811 65175
rect 208839 65147 208887 65175
rect 208577 65113 208887 65147
rect 208577 65085 208625 65113
rect 208653 65085 208687 65113
rect 208715 65085 208749 65113
rect 208777 65085 208811 65113
rect 208839 65085 208887 65113
rect 208577 65051 208887 65085
rect 208577 65023 208625 65051
rect 208653 65023 208687 65051
rect 208715 65023 208749 65051
rect 208777 65023 208811 65051
rect 208839 65023 208887 65051
rect 208577 64989 208887 65023
rect 208577 64961 208625 64989
rect 208653 64961 208687 64989
rect 208715 64961 208749 64989
rect 208777 64961 208811 64989
rect 208839 64961 208887 64989
rect 208577 56175 208887 64961
rect 208577 56147 208625 56175
rect 208653 56147 208687 56175
rect 208715 56147 208749 56175
rect 208777 56147 208811 56175
rect 208839 56147 208887 56175
rect 208577 56113 208887 56147
rect 208577 56085 208625 56113
rect 208653 56085 208687 56113
rect 208715 56085 208749 56113
rect 208777 56085 208811 56113
rect 208839 56085 208887 56113
rect 208577 56051 208887 56085
rect 208577 56023 208625 56051
rect 208653 56023 208687 56051
rect 208715 56023 208749 56051
rect 208777 56023 208811 56051
rect 208839 56023 208887 56051
rect 208577 55989 208887 56023
rect 208577 55961 208625 55989
rect 208653 55961 208687 55989
rect 208715 55961 208749 55989
rect 208777 55961 208811 55989
rect 208839 55961 208887 55989
rect 208577 47175 208887 55961
rect 208577 47147 208625 47175
rect 208653 47147 208687 47175
rect 208715 47147 208749 47175
rect 208777 47147 208811 47175
rect 208839 47147 208887 47175
rect 208577 47113 208887 47147
rect 208577 47085 208625 47113
rect 208653 47085 208687 47113
rect 208715 47085 208749 47113
rect 208777 47085 208811 47113
rect 208839 47085 208887 47113
rect 208577 47051 208887 47085
rect 208577 47023 208625 47051
rect 208653 47023 208687 47051
rect 208715 47023 208749 47051
rect 208777 47023 208811 47051
rect 208839 47023 208887 47051
rect 208577 46989 208887 47023
rect 208577 46961 208625 46989
rect 208653 46961 208687 46989
rect 208715 46961 208749 46989
rect 208777 46961 208811 46989
rect 208839 46961 208887 46989
rect 208577 38175 208887 46961
rect 208577 38147 208625 38175
rect 208653 38147 208687 38175
rect 208715 38147 208749 38175
rect 208777 38147 208811 38175
rect 208839 38147 208887 38175
rect 208577 38113 208887 38147
rect 208577 38085 208625 38113
rect 208653 38085 208687 38113
rect 208715 38085 208749 38113
rect 208777 38085 208811 38113
rect 208839 38085 208887 38113
rect 208577 38051 208887 38085
rect 208577 38023 208625 38051
rect 208653 38023 208687 38051
rect 208715 38023 208749 38051
rect 208777 38023 208811 38051
rect 208839 38023 208887 38051
rect 208577 37989 208887 38023
rect 208577 37961 208625 37989
rect 208653 37961 208687 37989
rect 208715 37961 208749 37989
rect 208777 37961 208811 37989
rect 208839 37961 208887 37989
rect 208577 29175 208887 37961
rect 208577 29147 208625 29175
rect 208653 29147 208687 29175
rect 208715 29147 208749 29175
rect 208777 29147 208811 29175
rect 208839 29147 208887 29175
rect 208577 29113 208887 29147
rect 208577 29085 208625 29113
rect 208653 29085 208687 29113
rect 208715 29085 208749 29113
rect 208777 29085 208811 29113
rect 208839 29085 208887 29113
rect 208577 29051 208887 29085
rect 208577 29023 208625 29051
rect 208653 29023 208687 29051
rect 208715 29023 208749 29051
rect 208777 29023 208811 29051
rect 208839 29023 208887 29051
rect 208577 28989 208887 29023
rect 208577 28961 208625 28989
rect 208653 28961 208687 28989
rect 208715 28961 208749 28989
rect 208777 28961 208811 28989
rect 208839 28961 208887 28989
rect 208577 20175 208887 28961
rect 208577 20147 208625 20175
rect 208653 20147 208687 20175
rect 208715 20147 208749 20175
rect 208777 20147 208811 20175
rect 208839 20147 208887 20175
rect 208577 20113 208887 20147
rect 208577 20085 208625 20113
rect 208653 20085 208687 20113
rect 208715 20085 208749 20113
rect 208777 20085 208811 20113
rect 208839 20085 208887 20113
rect 208577 20051 208887 20085
rect 208577 20023 208625 20051
rect 208653 20023 208687 20051
rect 208715 20023 208749 20051
rect 208777 20023 208811 20051
rect 208839 20023 208887 20051
rect 208577 19989 208887 20023
rect 208577 19961 208625 19989
rect 208653 19961 208687 19989
rect 208715 19961 208749 19989
rect 208777 19961 208811 19989
rect 208839 19961 208887 19989
rect 208577 11175 208887 19961
rect 208577 11147 208625 11175
rect 208653 11147 208687 11175
rect 208715 11147 208749 11175
rect 208777 11147 208811 11175
rect 208839 11147 208887 11175
rect 208577 11113 208887 11147
rect 208577 11085 208625 11113
rect 208653 11085 208687 11113
rect 208715 11085 208749 11113
rect 208777 11085 208811 11113
rect 208839 11085 208887 11113
rect 208577 11051 208887 11085
rect 208577 11023 208625 11051
rect 208653 11023 208687 11051
rect 208715 11023 208749 11051
rect 208777 11023 208811 11051
rect 208839 11023 208887 11051
rect 208577 10989 208887 11023
rect 208577 10961 208625 10989
rect 208653 10961 208687 10989
rect 208715 10961 208749 10989
rect 208777 10961 208811 10989
rect 208839 10961 208887 10989
rect 208577 2175 208887 10961
rect 208577 2147 208625 2175
rect 208653 2147 208687 2175
rect 208715 2147 208749 2175
rect 208777 2147 208811 2175
rect 208839 2147 208887 2175
rect 208577 2113 208887 2147
rect 208577 2085 208625 2113
rect 208653 2085 208687 2113
rect 208715 2085 208749 2113
rect 208777 2085 208811 2113
rect 208839 2085 208887 2113
rect 208577 2051 208887 2085
rect 208577 2023 208625 2051
rect 208653 2023 208687 2051
rect 208715 2023 208749 2051
rect 208777 2023 208811 2051
rect 208839 2023 208887 2051
rect 208577 1989 208887 2023
rect 208577 1961 208625 1989
rect 208653 1961 208687 1989
rect 208715 1961 208749 1989
rect 208777 1961 208811 1989
rect 208839 1961 208887 1989
rect 208577 -80 208887 1961
rect 208577 -108 208625 -80
rect 208653 -108 208687 -80
rect 208715 -108 208749 -80
rect 208777 -108 208811 -80
rect 208839 -108 208887 -80
rect 208577 -142 208887 -108
rect 208577 -170 208625 -142
rect 208653 -170 208687 -142
rect 208715 -170 208749 -142
rect 208777 -170 208811 -142
rect 208839 -170 208887 -142
rect 208577 -204 208887 -170
rect 208577 -232 208625 -204
rect 208653 -232 208687 -204
rect 208715 -232 208749 -204
rect 208777 -232 208811 -204
rect 208839 -232 208887 -204
rect 208577 -266 208887 -232
rect 208577 -294 208625 -266
rect 208653 -294 208687 -266
rect 208715 -294 208749 -266
rect 208777 -294 208811 -266
rect 208839 -294 208887 -266
rect 208577 -822 208887 -294
rect 210437 299086 210747 299134
rect 210437 299058 210485 299086
rect 210513 299058 210547 299086
rect 210575 299058 210609 299086
rect 210637 299058 210671 299086
rect 210699 299058 210747 299086
rect 210437 299024 210747 299058
rect 210437 298996 210485 299024
rect 210513 298996 210547 299024
rect 210575 298996 210609 299024
rect 210637 298996 210671 299024
rect 210699 298996 210747 299024
rect 210437 298962 210747 298996
rect 210437 298934 210485 298962
rect 210513 298934 210547 298962
rect 210575 298934 210609 298962
rect 210637 298934 210671 298962
rect 210699 298934 210747 298962
rect 210437 298900 210747 298934
rect 210437 298872 210485 298900
rect 210513 298872 210547 298900
rect 210575 298872 210609 298900
rect 210637 298872 210671 298900
rect 210699 298872 210747 298900
rect 210437 293175 210747 298872
rect 210437 293147 210485 293175
rect 210513 293147 210547 293175
rect 210575 293147 210609 293175
rect 210637 293147 210671 293175
rect 210699 293147 210747 293175
rect 210437 293113 210747 293147
rect 210437 293085 210485 293113
rect 210513 293085 210547 293113
rect 210575 293085 210609 293113
rect 210637 293085 210671 293113
rect 210699 293085 210747 293113
rect 210437 293051 210747 293085
rect 210437 293023 210485 293051
rect 210513 293023 210547 293051
rect 210575 293023 210609 293051
rect 210637 293023 210671 293051
rect 210699 293023 210747 293051
rect 210437 292989 210747 293023
rect 210437 292961 210485 292989
rect 210513 292961 210547 292989
rect 210575 292961 210609 292989
rect 210637 292961 210671 292989
rect 210699 292961 210747 292989
rect 210437 284175 210747 292961
rect 210437 284147 210485 284175
rect 210513 284147 210547 284175
rect 210575 284147 210609 284175
rect 210637 284147 210671 284175
rect 210699 284147 210747 284175
rect 210437 284113 210747 284147
rect 210437 284085 210485 284113
rect 210513 284085 210547 284113
rect 210575 284085 210609 284113
rect 210637 284085 210671 284113
rect 210699 284085 210747 284113
rect 210437 284051 210747 284085
rect 210437 284023 210485 284051
rect 210513 284023 210547 284051
rect 210575 284023 210609 284051
rect 210637 284023 210671 284051
rect 210699 284023 210747 284051
rect 210437 283989 210747 284023
rect 210437 283961 210485 283989
rect 210513 283961 210547 283989
rect 210575 283961 210609 283989
rect 210637 283961 210671 283989
rect 210699 283961 210747 283989
rect 210437 275175 210747 283961
rect 210437 275147 210485 275175
rect 210513 275147 210547 275175
rect 210575 275147 210609 275175
rect 210637 275147 210671 275175
rect 210699 275147 210747 275175
rect 210437 275113 210747 275147
rect 210437 275085 210485 275113
rect 210513 275085 210547 275113
rect 210575 275085 210609 275113
rect 210637 275085 210671 275113
rect 210699 275085 210747 275113
rect 210437 275051 210747 275085
rect 210437 275023 210485 275051
rect 210513 275023 210547 275051
rect 210575 275023 210609 275051
rect 210637 275023 210671 275051
rect 210699 275023 210747 275051
rect 210437 274989 210747 275023
rect 210437 274961 210485 274989
rect 210513 274961 210547 274989
rect 210575 274961 210609 274989
rect 210637 274961 210671 274989
rect 210699 274961 210747 274989
rect 210437 266175 210747 274961
rect 210437 266147 210485 266175
rect 210513 266147 210547 266175
rect 210575 266147 210609 266175
rect 210637 266147 210671 266175
rect 210699 266147 210747 266175
rect 210437 266113 210747 266147
rect 210437 266085 210485 266113
rect 210513 266085 210547 266113
rect 210575 266085 210609 266113
rect 210637 266085 210671 266113
rect 210699 266085 210747 266113
rect 210437 266051 210747 266085
rect 210437 266023 210485 266051
rect 210513 266023 210547 266051
rect 210575 266023 210609 266051
rect 210637 266023 210671 266051
rect 210699 266023 210747 266051
rect 210437 265989 210747 266023
rect 210437 265961 210485 265989
rect 210513 265961 210547 265989
rect 210575 265961 210609 265989
rect 210637 265961 210671 265989
rect 210699 265961 210747 265989
rect 210437 257175 210747 265961
rect 210437 257147 210485 257175
rect 210513 257147 210547 257175
rect 210575 257147 210609 257175
rect 210637 257147 210671 257175
rect 210699 257147 210747 257175
rect 210437 257113 210747 257147
rect 210437 257085 210485 257113
rect 210513 257085 210547 257113
rect 210575 257085 210609 257113
rect 210637 257085 210671 257113
rect 210699 257085 210747 257113
rect 210437 257051 210747 257085
rect 210437 257023 210485 257051
rect 210513 257023 210547 257051
rect 210575 257023 210609 257051
rect 210637 257023 210671 257051
rect 210699 257023 210747 257051
rect 210437 256989 210747 257023
rect 210437 256961 210485 256989
rect 210513 256961 210547 256989
rect 210575 256961 210609 256989
rect 210637 256961 210671 256989
rect 210699 256961 210747 256989
rect 210437 248175 210747 256961
rect 210437 248147 210485 248175
rect 210513 248147 210547 248175
rect 210575 248147 210609 248175
rect 210637 248147 210671 248175
rect 210699 248147 210747 248175
rect 210437 248113 210747 248147
rect 210437 248085 210485 248113
rect 210513 248085 210547 248113
rect 210575 248085 210609 248113
rect 210637 248085 210671 248113
rect 210699 248085 210747 248113
rect 210437 248051 210747 248085
rect 210437 248023 210485 248051
rect 210513 248023 210547 248051
rect 210575 248023 210609 248051
rect 210637 248023 210671 248051
rect 210699 248023 210747 248051
rect 210437 247989 210747 248023
rect 210437 247961 210485 247989
rect 210513 247961 210547 247989
rect 210575 247961 210609 247989
rect 210637 247961 210671 247989
rect 210699 247961 210747 247989
rect 210437 239175 210747 247961
rect 210437 239147 210485 239175
rect 210513 239147 210547 239175
rect 210575 239147 210609 239175
rect 210637 239147 210671 239175
rect 210699 239147 210747 239175
rect 210437 239113 210747 239147
rect 210437 239085 210485 239113
rect 210513 239085 210547 239113
rect 210575 239085 210609 239113
rect 210637 239085 210671 239113
rect 210699 239085 210747 239113
rect 210437 239051 210747 239085
rect 210437 239023 210485 239051
rect 210513 239023 210547 239051
rect 210575 239023 210609 239051
rect 210637 239023 210671 239051
rect 210699 239023 210747 239051
rect 210437 238989 210747 239023
rect 210437 238961 210485 238989
rect 210513 238961 210547 238989
rect 210575 238961 210609 238989
rect 210637 238961 210671 238989
rect 210699 238961 210747 238989
rect 210437 230175 210747 238961
rect 210437 230147 210485 230175
rect 210513 230147 210547 230175
rect 210575 230147 210609 230175
rect 210637 230147 210671 230175
rect 210699 230147 210747 230175
rect 210437 230113 210747 230147
rect 210437 230085 210485 230113
rect 210513 230085 210547 230113
rect 210575 230085 210609 230113
rect 210637 230085 210671 230113
rect 210699 230085 210747 230113
rect 210437 230051 210747 230085
rect 210437 230023 210485 230051
rect 210513 230023 210547 230051
rect 210575 230023 210609 230051
rect 210637 230023 210671 230051
rect 210699 230023 210747 230051
rect 210437 229989 210747 230023
rect 210437 229961 210485 229989
rect 210513 229961 210547 229989
rect 210575 229961 210609 229989
rect 210637 229961 210671 229989
rect 210699 229961 210747 229989
rect 210437 221175 210747 229961
rect 210437 221147 210485 221175
rect 210513 221147 210547 221175
rect 210575 221147 210609 221175
rect 210637 221147 210671 221175
rect 210699 221147 210747 221175
rect 210437 221113 210747 221147
rect 210437 221085 210485 221113
rect 210513 221085 210547 221113
rect 210575 221085 210609 221113
rect 210637 221085 210671 221113
rect 210699 221085 210747 221113
rect 210437 221051 210747 221085
rect 210437 221023 210485 221051
rect 210513 221023 210547 221051
rect 210575 221023 210609 221051
rect 210637 221023 210671 221051
rect 210699 221023 210747 221051
rect 210437 220989 210747 221023
rect 210437 220961 210485 220989
rect 210513 220961 210547 220989
rect 210575 220961 210609 220989
rect 210637 220961 210671 220989
rect 210699 220961 210747 220989
rect 210437 212175 210747 220961
rect 210437 212147 210485 212175
rect 210513 212147 210547 212175
rect 210575 212147 210609 212175
rect 210637 212147 210671 212175
rect 210699 212147 210747 212175
rect 210437 212113 210747 212147
rect 210437 212085 210485 212113
rect 210513 212085 210547 212113
rect 210575 212085 210609 212113
rect 210637 212085 210671 212113
rect 210699 212085 210747 212113
rect 210437 212051 210747 212085
rect 210437 212023 210485 212051
rect 210513 212023 210547 212051
rect 210575 212023 210609 212051
rect 210637 212023 210671 212051
rect 210699 212023 210747 212051
rect 210437 211989 210747 212023
rect 210437 211961 210485 211989
rect 210513 211961 210547 211989
rect 210575 211961 210609 211989
rect 210637 211961 210671 211989
rect 210699 211961 210747 211989
rect 210437 203175 210747 211961
rect 210437 203147 210485 203175
rect 210513 203147 210547 203175
rect 210575 203147 210609 203175
rect 210637 203147 210671 203175
rect 210699 203147 210747 203175
rect 210437 203113 210747 203147
rect 210437 203085 210485 203113
rect 210513 203085 210547 203113
rect 210575 203085 210609 203113
rect 210637 203085 210671 203113
rect 210699 203085 210747 203113
rect 210437 203051 210747 203085
rect 210437 203023 210485 203051
rect 210513 203023 210547 203051
rect 210575 203023 210609 203051
rect 210637 203023 210671 203051
rect 210699 203023 210747 203051
rect 210437 202989 210747 203023
rect 210437 202961 210485 202989
rect 210513 202961 210547 202989
rect 210575 202961 210609 202989
rect 210637 202961 210671 202989
rect 210699 202961 210747 202989
rect 210437 194175 210747 202961
rect 210437 194147 210485 194175
rect 210513 194147 210547 194175
rect 210575 194147 210609 194175
rect 210637 194147 210671 194175
rect 210699 194147 210747 194175
rect 210437 194113 210747 194147
rect 210437 194085 210485 194113
rect 210513 194085 210547 194113
rect 210575 194085 210609 194113
rect 210637 194085 210671 194113
rect 210699 194085 210747 194113
rect 210437 194051 210747 194085
rect 210437 194023 210485 194051
rect 210513 194023 210547 194051
rect 210575 194023 210609 194051
rect 210637 194023 210671 194051
rect 210699 194023 210747 194051
rect 210437 193989 210747 194023
rect 210437 193961 210485 193989
rect 210513 193961 210547 193989
rect 210575 193961 210609 193989
rect 210637 193961 210671 193989
rect 210699 193961 210747 193989
rect 210437 185175 210747 193961
rect 210437 185147 210485 185175
rect 210513 185147 210547 185175
rect 210575 185147 210609 185175
rect 210637 185147 210671 185175
rect 210699 185147 210747 185175
rect 210437 185113 210747 185147
rect 210437 185085 210485 185113
rect 210513 185085 210547 185113
rect 210575 185085 210609 185113
rect 210637 185085 210671 185113
rect 210699 185085 210747 185113
rect 210437 185051 210747 185085
rect 210437 185023 210485 185051
rect 210513 185023 210547 185051
rect 210575 185023 210609 185051
rect 210637 185023 210671 185051
rect 210699 185023 210747 185051
rect 210437 184989 210747 185023
rect 210437 184961 210485 184989
rect 210513 184961 210547 184989
rect 210575 184961 210609 184989
rect 210637 184961 210671 184989
rect 210699 184961 210747 184989
rect 210437 176175 210747 184961
rect 210437 176147 210485 176175
rect 210513 176147 210547 176175
rect 210575 176147 210609 176175
rect 210637 176147 210671 176175
rect 210699 176147 210747 176175
rect 210437 176113 210747 176147
rect 210437 176085 210485 176113
rect 210513 176085 210547 176113
rect 210575 176085 210609 176113
rect 210637 176085 210671 176113
rect 210699 176085 210747 176113
rect 210437 176051 210747 176085
rect 210437 176023 210485 176051
rect 210513 176023 210547 176051
rect 210575 176023 210609 176051
rect 210637 176023 210671 176051
rect 210699 176023 210747 176051
rect 210437 175989 210747 176023
rect 210437 175961 210485 175989
rect 210513 175961 210547 175989
rect 210575 175961 210609 175989
rect 210637 175961 210671 175989
rect 210699 175961 210747 175989
rect 210437 167175 210747 175961
rect 210437 167147 210485 167175
rect 210513 167147 210547 167175
rect 210575 167147 210609 167175
rect 210637 167147 210671 167175
rect 210699 167147 210747 167175
rect 210437 167113 210747 167147
rect 210437 167085 210485 167113
rect 210513 167085 210547 167113
rect 210575 167085 210609 167113
rect 210637 167085 210671 167113
rect 210699 167085 210747 167113
rect 210437 167051 210747 167085
rect 210437 167023 210485 167051
rect 210513 167023 210547 167051
rect 210575 167023 210609 167051
rect 210637 167023 210671 167051
rect 210699 167023 210747 167051
rect 210437 166989 210747 167023
rect 210437 166961 210485 166989
rect 210513 166961 210547 166989
rect 210575 166961 210609 166989
rect 210637 166961 210671 166989
rect 210699 166961 210747 166989
rect 210437 158175 210747 166961
rect 210437 158147 210485 158175
rect 210513 158147 210547 158175
rect 210575 158147 210609 158175
rect 210637 158147 210671 158175
rect 210699 158147 210747 158175
rect 210437 158113 210747 158147
rect 210437 158085 210485 158113
rect 210513 158085 210547 158113
rect 210575 158085 210609 158113
rect 210637 158085 210671 158113
rect 210699 158085 210747 158113
rect 210437 158051 210747 158085
rect 210437 158023 210485 158051
rect 210513 158023 210547 158051
rect 210575 158023 210609 158051
rect 210637 158023 210671 158051
rect 210699 158023 210747 158051
rect 210437 157989 210747 158023
rect 210437 157961 210485 157989
rect 210513 157961 210547 157989
rect 210575 157961 210609 157989
rect 210637 157961 210671 157989
rect 210699 157961 210747 157989
rect 210437 149175 210747 157961
rect 210437 149147 210485 149175
rect 210513 149147 210547 149175
rect 210575 149147 210609 149175
rect 210637 149147 210671 149175
rect 210699 149147 210747 149175
rect 210437 149113 210747 149147
rect 210437 149085 210485 149113
rect 210513 149085 210547 149113
rect 210575 149085 210609 149113
rect 210637 149085 210671 149113
rect 210699 149085 210747 149113
rect 210437 149051 210747 149085
rect 210437 149023 210485 149051
rect 210513 149023 210547 149051
rect 210575 149023 210609 149051
rect 210637 149023 210671 149051
rect 210699 149023 210747 149051
rect 210437 148989 210747 149023
rect 210437 148961 210485 148989
rect 210513 148961 210547 148989
rect 210575 148961 210609 148989
rect 210637 148961 210671 148989
rect 210699 148961 210747 148989
rect 210437 140175 210747 148961
rect 210437 140147 210485 140175
rect 210513 140147 210547 140175
rect 210575 140147 210609 140175
rect 210637 140147 210671 140175
rect 210699 140147 210747 140175
rect 210437 140113 210747 140147
rect 210437 140085 210485 140113
rect 210513 140085 210547 140113
rect 210575 140085 210609 140113
rect 210637 140085 210671 140113
rect 210699 140085 210747 140113
rect 210437 140051 210747 140085
rect 210437 140023 210485 140051
rect 210513 140023 210547 140051
rect 210575 140023 210609 140051
rect 210637 140023 210671 140051
rect 210699 140023 210747 140051
rect 210437 139989 210747 140023
rect 210437 139961 210485 139989
rect 210513 139961 210547 139989
rect 210575 139961 210609 139989
rect 210637 139961 210671 139989
rect 210699 139961 210747 139989
rect 210437 131175 210747 139961
rect 210437 131147 210485 131175
rect 210513 131147 210547 131175
rect 210575 131147 210609 131175
rect 210637 131147 210671 131175
rect 210699 131147 210747 131175
rect 210437 131113 210747 131147
rect 210437 131085 210485 131113
rect 210513 131085 210547 131113
rect 210575 131085 210609 131113
rect 210637 131085 210671 131113
rect 210699 131085 210747 131113
rect 210437 131051 210747 131085
rect 210437 131023 210485 131051
rect 210513 131023 210547 131051
rect 210575 131023 210609 131051
rect 210637 131023 210671 131051
rect 210699 131023 210747 131051
rect 210437 130989 210747 131023
rect 210437 130961 210485 130989
rect 210513 130961 210547 130989
rect 210575 130961 210609 130989
rect 210637 130961 210671 130989
rect 210699 130961 210747 130989
rect 210437 122175 210747 130961
rect 210437 122147 210485 122175
rect 210513 122147 210547 122175
rect 210575 122147 210609 122175
rect 210637 122147 210671 122175
rect 210699 122147 210747 122175
rect 210437 122113 210747 122147
rect 210437 122085 210485 122113
rect 210513 122085 210547 122113
rect 210575 122085 210609 122113
rect 210637 122085 210671 122113
rect 210699 122085 210747 122113
rect 210437 122051 210747 122085
rect 210437 122023 210485 122051
rect 210513 122023 210547 122051
rect 210575 122023 210609 122051
rect 210637 122023 210671 122051
rect 210699 122023 210747 122051
rect 210437 121989 210747 122023
rect 210437 121961 210485 121989
rect 210513 121961 210547 121989
rect 210575 121961 210609 121989
rect 210637 121961 210671 121989
rect 210699 121961 210747 121989
rect 210437 113175 210747 121961
rect 210437 113147 210485 113175
rect 210513 113147 210547 113175
rect 210575 113147 210609 113175
rect 210637 113147 210671 113175
rect 210699 113147 210747 113175
rect 210437 113113 210747 113147
rect 210437 113085 210485 113113
rect 210513 113085 210547 113113
rect 210575 113085 210609 113113
rect 210637 113085 210671 113113
rect 210699 113085 210747 113113
rect 210437 113051 210747 113085
rect 210437 113023 210485 113051
rect 210513 113023 210547 113051
rect 210575 113023 210609 113051
rect 210637 113023 210671 113051
rect 210699 113023 210747 113051
rect 210437 112989 210747 113023
rect 210437 112961 210485 112989
rect 210513 112961 210547 112989
rect 210575 112961 210609 112989
rect 210637 112961 210671 112989
rect 210699 112961 210747 112989
rect 210437 104175 210747 112961
rect 210437 104147 210485 104175
rect 210513 104147 210547 104175
rect 210575 104147 210609 104175
rect 210637 104147 210671 104175
rect 210699 104147 210747 104175
rect 210437 104113 210747 104147
rect 210437 104085 210485 104113
rect 210513 104085 210547 104113
rect 210575 104085 210609 104113
rect 210637 104085 210671 104113
rect 210699 104085 210747 104113
rect 210437 104051 210747 104085
rect 210437 104023 210485 104051
rect 210513 104023 210547 104051
rect 210575 104023 210609 104051
rect 210637 104023 210671 104051
rect 210699 104023 210747 104051
rect 210437 103989 210747 104023
rect 210437 103961 210485 103989
rect 210513 103961 210547 103989
rect 210575 103961 210609 103989
rect 210637 103961 210671 103989
rect 210699 103961 210747 103989
rect 210437 95175 210747 103961
rect 210437 95147 210485 95175
rect 210513 95147 210547 95175
rect 210575 95147 210609 95175
rect 210637 95147 210671 95175
rect 210699 95147 210747 95175
rect 210437 95113 210747 95147
rect 210437 95085 210485 95113
rect 210513 95085 210547 95113
rect 210575 95085 210609 95113
rect 210637 95085 210671 95113
rect 210699 95085 210747 95113
rect 210437 95051 210747 95085
rect 210437 95023 210485 95051
rect 210513 95023 210547 95051
rect 210575 95023 210609 95051
rect 210637 95023 210671 95051
rect 210699 95023 210747 95051
rect 210437 94989 210747 95023
rect 210437 94961 210485 94989
rect 210513 94961 210547 94989
rect 210575 94961 210609 94989
rect 210637 94961 210671 94989
rect 210699 94961 210747 94989
rect 210437 86175 210747 94961
rect 210437 86147 210485 86175
rect 210513 86147 210547 86175
rect 210575 86147 210609 86175
rect 210637 86147 210671 86175
rect 210699 86147 210747 86175
rect 210437 86113 210747 86147
rect 210437 86085 210485 86113
rect 210513 86085 210547 86113
rect 210575 86085 210609 86113
rect 210637 86085 210671 86113
rect 210699 86085 210747 86113
rect 210437 86051 210747 86085
rect 210437 86023 210485 86051
rect 210513 86023 210547 86051
rect 210575 86023 210609 86051
rect 210637 86023 210671 86051
rect 210699 86023 210747 86051
rect 210437 85989 210747 86023
rect 210437 85961 210485 85989
rect 210513 85961 210547 85989
rect 210575 85961 210609 85989
rect 210637 85961 210671 85989
rect 210699 85961 210747 85989
rect 210437 77175 210747 85961
rect 210437 77147 210485 77175
rect 210513 77147 210547 77175
rect 210575 77147 210609 77175
rect 210637 77147 210671 77175
rect 210699 77147 210747 77175
rect 210437 77113 210747 77147
rect 210437 77085 210485 77113
rect 210513 77085 210547 77113
rect 210575 77085 210609 77113
rect 210637 77085 210671 77113
rect 210699 77085 210747 77113
rect 210437 77051 210747 77085
rect 210437 77023 210485 77051
rect 210513 77023 210547 77051
rect 210575 77023 210609 77051
rect 210637 77023 210671 77051
rect 210699 77023 210747 77051
rect 210437 76989 210747 77023
rect 210437 76961 210485 76989
rect 210513 76961 210547 76989
rect 210575 76961 210609 76989
rect 210637 76961 210671 76989
rect 210699 76961 210747 76989
rect 210437 68175 210747 76961
rect 210437 68147 210485 68175
rect 210513 68147 210547 68175
rect 210575 68147 210609 68175
rect 210637 68147 210671 68175
rect 210699 68147 210747 68175
rect 210437 68113 210747 68147
rect 210437 68085 210485 68113
rect 210513 68085 210547 68113
rect 210575 68085 210609 68113
rect 210637 68085 210671 68113
rect 210699 68085 210747 68113
rect 210437 68051 210747 68085
rect 210437 68023 210485 68051
rect 210513 68023 210547 68051
rect 210575 68023 210609 68051
rect 210637 68023 210671 68051
rect 210699 68023 210747 68051
rect 210437 67989 210747 68023
rect 210437 67961 210485 67989
rect 210513 67961 210547 67989
rect 210575 67961 210609 67989
rect 210637 67961 210671 67989
rect 210699 67961 210747 67989
rect 210437 59175 210747 67961
rect 210437 59147 210485 59175
rect 210513 59147 210547 59175
rect 210575 59147 210609 59175
rect 210637 59147 210671 59175
rect 210699 59147 210747 59175
rect 210437 59113 210747 59147
rect 210437 59085 210485 59113
rect 210513 59085 210547 59113
rect 210575 59085 210609 59113
rect 210637 59085 210671 59113
rect 210699 59085 210747 59113
rect 210437 59051 210747 59085
rect 210437 59023 210485 59051
rect 210513 59023 210547 59051
rect 210575 59023 210609 59051
rect 210637 59023 210671 59051
rect 210699 59023 210747 59051
rect 210437 58989 210747 59023
rect 210437 58961 210485 58989
rect 210513 58961 210547 58989
rect 210575 58961 210609 58989
rect 210637 58961 210671 58989
rect 210699 58961 210747 58989
rect 210437 50175 210747 58961
rect 210437 50147 210485 50175
rect 210513 50147 210547 50175
rect 210575 50147 210609 50175
rect 210637 50147 210671 50175
rect 210699 50147 210747 50175
rect 210437 50113 210747 50147
rect 210437 50085 210485 50113
rect 210513 50085 210547 50113
rect 210575 50085 210609 50113
rect 210637 50085 210671 50113
rect 210699 50085 210747 50113
rect 210437 50051 210747 50085
rect 210437 50023 210485 50051
rect 210513 50023 210547 50051
rect 210575 50023 210609 50051
rect 210637 50023 210671 50051
rect 210699 50023 210747 50051
rect 210437 49989 210747 50023
rect 210437 49961 210485 49989
rect 210513 49961 210547 49989
rect 210575 49961 210609 49989
rect 210637 49961 210671 49989
rect 210699 49961 210747 49989
rect 210437 41175 210747 49961
rect 210437 41147 210485 41175
rect 210513 41147 210547 41175
rect 210575 41147 210609 41175
rect 210637 41147 210671 41175
rect 210699 41147 210747 41175
rect 210437 41113 210747 41147
rect 210437 41085 210485 41113
rect 210513 41085 210547 41113
rect 210575 41085 210609 41113
rect 210637 41085 210671 41113
rect 210699 41085 210747 41113
rect 210437 41051 210747 41085
rect 210437 41023 210485 41051
rect 210513 41023 210547 41051
rect 210575 41023 210609 41051
rect 210637 41023 210671 41051
rect 210699 41023 210747 41051
rect 210437 40989 210747 41023
rect 210437 40961 210485 40989
rect 210513 40961 210547 40989
rect 210575 40961 210609 40989
rect 210637 40961 210671 40989
rect 210699 40961 210747 40989
rect 210437 32175 210747 40961
rect 210437 32147 210485 32175
rect 210513 32147 210547 32175
rect 210575 32147 210609 32175
rect 210637 32147 210671 32175
rect 210699 32147 210747 32175
rect 210437 32113 210747 32147
rect 210437 32085 210485 32113
rect 210513 32085 210547 32113
rect 210575 32085 210609 32113
rect 210637 32085 210671 32113
rect 210699 32085 210747 32113
rect 210437 32051 210747 32085
rect 210437 32023 210485 32051
rect 210513 32023 210547 32051
rect 210575 32023 210609 32051
rect 210637 32023 210671 32051
rect 210699 32023 210747 32051
rect 210437 31989 210747 32023
rect 210437 31961 210485 31989
rect 210513 31961 210547 31989
rect 210575 31961 210609 31989
rect 210637 31961 210671 31989
rect 210699 31961 210747 31989
rect 210437 23175 210747 31961
rect 210437 23147 210485 23175
rect 210513 23147 210547 23175
rect 210575 23147 210609 23175
rect 210637 23147 210671 23175
rect 210699 23147 210747 23175
rect 210437 23113 210747 23147
rect 210437 23085 210485 23113
rect 210513 23085 210547 23113
rect 210575 23085 210609 23113
rect 210637 23085 210671 23113
rect 210699 23085 210747 23113
rect 210437 23051 210747 23085
rect 210437 23023 210485 23051
rect 210513 23023 210547 23051
rect 210575 23023 210609 23051
rect 210637 23023 210671 23051
rect 210699 23023 210747 23051
rect 210437 22989 210747 23023
rect 210437 22961 210485 22989
rect 210513 22961 210547 22989
rect 210575 22961 210609 22989
rect 210637 22961 210671 22989
rect 210699 22961 210747 22989
rect 210437 14175 210747 22961
rect 210437 14147 210485 14175
rect 210513 14147 210547 14175
rect 210575 14147 210609 14175
rect 210637 14147 210671 14175
rect 210699 14147 210747 14175
rect 210437 14113 210747 14147
rect 210437 14085 210485 14113
rect 210513 14085 210547 14113
rect 210575 14085 210609 14113
rect 210637 14085 210671 14113
rect 210699 14085 210747 14113
rect 210437 14051 210747 14085
rect 210437 14023 210485 14051
rect 210513 14023 210547 14051
rect 210575 14023 210609 14051
rect 210637 14023 210671 14051
rect 210699 14023 210747 14051
rect 210437 13989 210747 14023
rect 210437 13961 210485 13989
rect 210513 13961 210547 13989
rect 210575 13961 210609 13989
rect 210637 13961 210671 13989
rect 210699 13961 210747 13989
rect 210437 5175 210747 13961
rect 210437 5147 210485 5175
rect 210513 5147 210547 5175
rect 210575 5147 210609 5175
rect 210637 5147 210671 5175
rect 210699 5147 210747 5175
rect 210437 5113 210747 5147
rect 210437 5085 210485 5113
rect 210513 5085 210547 5113
rect 210575 5085 210609 5113
rect 210637 5085 210671 5113
rect 210699 5085 210747 5113
rect 210437 5051 210747 5085
rect 210437 5023 210485 5051
rect 210513 5023 210547 5051
rect 210575 5023 210609 5051
rect 210637 5023 210671 5051
rect 210699 5023 210747 5051
rect 210437 4989 210747 5023
rect 210437 4961 210485 4989
rect 210513 4961 210547 4989
rect 210575 4961 210609 4989
rect 210637 4961 210671 4989
rect 210699 4961 210747 4989
rect 210437 -560 210747 4961
rect 210437 -588 210485 -560
rect 210513 -588 210547 -560
rect 210575 -588 210609 -560
rect 210637 -588 210671 -560
rect 210699 -588 210747 -560
rect 210437 -622 210747 -588
rect 210437 -650 210485 -622
rect 210513 -650 210547 -622
rect 210575 -650 210609 -622
rect 210637 -650 210671 -622
rect 210699 -650 210747 -622
rect 210437 -684 210747 -650
rect 210437 -712 210485 -684
rect 210513 -712 210547 -684
rect 210575 -712 210609 -684
rect 210637 -712 210671 -684
rect 210699 -712 210747 -684
rect 210437 -746 210747 -712
rect 210437 -774 210485 -746
rect 210513 -774 210547 -746
rect 210575 -774 210609 -746
rect 210637 -774 210671 -746
rect 210699 -774 210747 -746
rect 210437 -822 210747 -774
rect 217577 298606 217887 299134
rect 217577 298578 217625 298606
rect 217653 298578 217687 298606
rect 217715 298578 217749 298606
rect 217777 298578 217811 298606
rect 217839 298578 217887 298606
rect 217577 298544 217887 298578
rect 217577 298516 217625 298544
rect 217653 298516 217687 298544
rect 217715 298516 217749 298544
rect 217777 298516 217811 298544
rect 217839 298516 217887 298544
rect 217577 298482 217887 298516
rect 217577 298454 217625 298482
rect 217653 298454 217687 298482
rect 217715 298454 217749 298482
rect 217777 298454 217811 298482
rect 217839 298454 217887 298482
rect 217577 298420 217887 298454
rect 217577 298392 217625 298420
rect 217653 298392 217687 298420
rect 217715 298392 217749 298420
rect 217777 298392 217811 298420
rect 217839 298392 217887 298420
rect 217577 290175 217887 298392
rect 217577 290147 217625 290175
rect 217653 290147 217687 290175
rect 217715 290147 217749 290175
rect 217777 290147 217811 290175
rect 217839 290147 217887 290175
rect 217577 290113 217887 290147
rect 217577 290085 217625 290113
rect 217653 290085 217687 290113
rect 217715 290085 217749 290113
rect 217777 290085 217811 290113
rect 217839 290085 217887 290113
rect 217577 290051 217887 290085
rect 217577 290023 217625 290051
rect 217653 290023 217687 290051
rect 217715 290023 217749 290051
rect 217777 290023 217811 290051
rect 217839 290023 217887 290051
rect 217577 289989 217887 290023
rect 217577 289961 217625 289989
rect 217653 289961 217687 289989
rect 217715 289961 217749 289989
rect 217777 289961 217811 289989
rect 217839 289961 217887 289989
rect 217577 281175 217887 289961
rect 217577 281147 217625 281175
rect 217653 281147 217687 281175
rect 217715 281147 217749 281175
rect 217777 281147 217811 281175
rect 217839 281147 217887 281175
rect 217577 281113 217887 281147
rect 217577 281085 217625 281113
rect 217653 281085 217687 281113
rect 217715 281085 217749 281113
rect 217777 281085 217811 281113
rect 217839 281085 217887 281113
rect 217577 281051 217887 281085
rect 217577 281023 217625 281051
rect 217653 281023 217687 281051
rect 217715 281023 217749 281051
rect 217777 281023 217811 281051
rect 217839 281023 217887 281051
rect 217577 280989 217887 281023
rect 217577 280961 217625 280989
rect 217653 280961 217687 280989
rect 217715 280961 217749 280989
rect 217777 280961 217811 280989
rect 217839 280961 217887 280989
rect 217577 272175 217887 280961
rect 217577 272147 217625 272175
rect 217653 272147 217687 272175
rect 217715 272147 217749 272175
rect 217777 272147 217811 272175
rect 217839 272147 217887 272175
rect 217577 272113 217887 272147
rect 217577 272085 217625 272113
rect 217653 272085 217687 272113
rect 217715 272085 217749 272113
rect 217777 272085 217811 272113
rect 217839 272085 217887 272113
rect 217577 272051 217887 272085
rect 217577 272023 217625 272051
rect 217653 272023 217687 272051
rect 217715 272023 217749 272051
rect 217777 272023 217811 272051
rect 217839 272023 217887 272051
rect 217577 271989 217887 272023
rect 217577 271961 217625 271989
rect 217653 271961 217687 271989
rect 217715 271961 217749 271989
rect 217777 271961 217811 271989
rect 217839 271961 217887 271989
rect 217577 263175 217887 271961
rect 217577 263147 217625 263175
rect 217653 263147 217687 263175
rect 217715 263147 217749 263175
rect 217777 263147 217811 263175
rect 217839 263147 217887 263175
rect 217577 263113 217887 263147
rect 217577 263085 217625 263113
rect 217653 263085 217687 263113
rect 217715 263085 217749 263113
rect 217777 263085 217811 263113
rect 217839 263085 217887 263113
rect 217577 263051 217887 263085
rect 217577 263023 217625 263051
rect 217653 263023 217687 263051
rect 217715 263023 217749 263051
rect 217777 263023 217811 263051
rect 217839 263023 217887 263051
rect 217577 262989 217887 263023
rect 217577 262961 217625 262989
rect 217653 262961 217687 262989
rect 217715 262961 217749 262989
rect 217777 262961 217811 262989
rect 217839 262961 217887 262989
rect 217577 254175 217887 262961
rect 217577 254147 217625 254175
rect 217653 254147 217687 254175
rect 217715 254147 217749 254175
rect 217777 254147 217811 254175
rect 217839 254147 217887 254175
rect 217577 254113 217887 254147
rect 217577 254085 217625 254113
rect 217653 254085 217687 254113
rect 217715 254085 217749 254113
rect 217777 254085 217811 254113
rect 217839 254085 217887 254113
rect 217577 254051 217887 254085
rect 217577 254023 217625 254051
rect 217653 254023 217687 254051
rect 217715 254023 217749 254051
rect 217777 254023 217811 254051
rect 217839 254023 217887 254051
rect 217577 253989 217887 254023
rect 217577 253961 217625 253989
rect 217653 253961 217687 253989
rect 217715 253961 217749 253989
rect 217777 253961 217811 253989
rect 217839 253961 217887 253989
rect 217577 245175 217887 253961
rect 217577 245147 217625 245175
rect 217653 245147 217687 245175
rect 217715 245147 217749 245175
rect 217777 245147 217811 245175
rect 217839 245147 217887 245175
rect 217577 245113 217887 245147
rect 217577 245085 217625 245113
rect 217653 245085 217687 245113
rect 217715 245085 217749 245113
rect 217777 245085 217811 245113
rect 217839 245085 217887 245113
rect 217577 245051 217887 245085
rect 217577 245023 217625 245051
rect 217653 245023 217687 245051
rect 217715 245023 217749 245051
rect 217777 245023 217811 245051
rect 217839 245023 217887 245051
rect 217577 244989 217887 245023
rect 217577 244961 217625 244989
rect 217653 244961 217687 244989
rect 217715 244961 217749 244989
rect 217777 244961 217811 244989
rect 217839 244961 217887 244989
rect 217577 236175 217887 244961
rect 217577 236147 217625 236175
rect 217653 236147 217687 236175
rect 217715 236147 217749 236175
rect 217777 236147 217811 236175
rect 217839 236147 217887 236175
rect 217577 236113 217887 236147
rect 217577 236085 217625 236113
rect 217653 236085 217687 236113
rect 217715 236085 217749 236113
rect 217777 236085 217811 236113
rect 217839 236085 217887 236113
rect 217577 236051 217887 236085
rect 217577 236023 217625 236051
rect 217653 236023 217687 236051
rect 217715 236023 217749 236051
rect 217777 236023 217811 236051
rect 217839 236023 217887 236051
rect 217577 235989 217887 236023
rect 217577 235961 217625 235989
rect 217653 235961 217687 235989
rect 217715 235961 217749 235989
rect 217777 235961 217811 235989
rect 217839 235961 217887 235989
rect 217577 227175 217887 235961
rect 217577 227147 217625 227175
rect 217653 227147 217687 227175
rect 217715 227147 217749 227175
rect 217777 227147 217811 227175
rect 217839 227147 217887 227175
rect 217577 227113 217887 227147
rect 217577 227085 217625 227113
rect 217653 227085 217687 227113
rect 217715 227085 217749 227113
rect 217777 227085 217811 227113
rect 217839 227085 217887 227113
rect 217577 227051 217887 227085
rect 217577 227023 217625 227051
rect 217653 227023 217687 227051
rect 217715 227023 217749 227051
rect 217777 227023 217811 227051
rect 217839 227023 217887 227051
rect 217577 226989 217887 227023
rect 217577 226961 217625 226989
rect 217653 226961 217687 226989
rect 217715 226961 217749 226989
rect 217777 226961 217811 226989
rect 217839 226961 217887 226989
rect 217577 218175 217887 226961
rect 217577 218147 217625 218175
rect 217653 218147 217687 218175
rect 217715 218147 217749 218175
rect 217777 218147 217811 218175
rect 217839 218147 217887 218175
rect 217577 218113 217887 218147
rect 217577 218085 217625 218113
rect 217653 218085 217687 218113
rect 217715 218085 217749 218113
rect 217777 218085 217811 218113
rect 217839 218085 217887 218113
rect 217577 218051 217887 218085
rect 217577 218023 217625 218051
rect 217653 218023 217687 218051
rect 217715 218023 217749 218051
rect 217777 218023 217811 218051
rect 217839 218023 217887 218051
rect 217577 217989 217887 218023
rect 217577 217961 217625 217989
rect 217653 217961 217687 217989
rect 217715 217961 217749 217989
rect 217777 217961 217811 217989
rect 217839 217961 217887 217989
rect 217577 209175 217887 217961
rect 217577 209147 217625 209175
rect 217653 209147 217687 209175
rect 217715 209147 217749 209175
rect 217777 209147 217811 209175
rect 217839 209147 217887 209175
rect 217577 209113 217887 209147
rect 217577 209085 217625 209113
rect 217653 209085 217687 209113
rect 217715 209085 217749 209113
rect 217777 209085 217811 209113
rect 217839 209085 217887 209113
rect 217577 209051 217887 209085
rect 217577 209023 217625 209051
rect 217653 209023 217687 209051
rect 217715 209023 217749 209051
rect 217777 209023 217811 209051
rect 217839 209023 217887 209051
rect 217577 208989 217887 209023
rect 217577 208961 217625 208989
rect 217653 208961 217687 208989
rect 217715 208961 217749 208989
rect 217777 208961 217811 208989
rect 217839 208961 217887 208989
rect 217577 200175 217887 208961
rect 217577 200147 217625 200175
rect 217653 200147 217687 200175
rect 217715 200147 217749 200175
rect 217777 200147 217811 200175
rect 217839 200147 217887 200175
rect 217577 200113 217887 200147
rect 217577 200085 217625 200113
rect 217653 200085 217687 200113
rect 217715 200085 217749 200113
rect 217777 200085 217811 200113
rect 217839 200085 217887 200113
rect 217577 200051 217887 200085
rect 217577 200023 217625 200051
rect 217653 200023 217687 200051
rect 217715 200023 217749 200051
rect 217777 200023 217811 200051
rect 217839 200023 217887 200051
rect 217577 199989 217887 200023
rect 217577 199961 217625 199989
rect 217653 199961 217687 199989
rect 217715 199961 217749 199989
rect 217777 199961 217811 199989
rect 217839 199961 217887 199989
rect 217577 191175 217887 199961
rect 217577 191147 217625 191175
rect 217653 191147 217687 191175
rect 217715 191147 217749 191175
rect 217777 191147 217811 191175
rect 217839 191147 217887 191175
rect 217577 191113 217887 191147
rect 217577 191085 217625 191113
rect 217653 191085 217687 191113
rect 217715 191085 217749 191113
rect 217777 191085 217811 191113
rect 217839 191085 217887 191113
rect 217577 191051 217887 191085
rect 217577 191023 217625 191051
rect 217653 191023 217687 191051
rect 217715 191023 217749 191051
rect 217777 191023 217811 191051
rect 217839 191023 217887 191051
rect 217577 190989 217887 191023
rect 217577 190961 217625 190989
rect 217653 190961 217687 190989
rect 217715 190961 217749 190989
rect 217777 190961 217811 190989
rect 217839 190961 217887 190989
rect 217577 182175 217887 190961
rect 217577 182147 217625 182175
rect 217653 182147 217687 182175
rect 217715 182147 217749 182175
rect 217777 182147 217811 182175
rect 217839 182147 217887 182175
rect 217577 182113 217887 182147
rect 217577 182085 217625 182113
rect 217653 182085 217687 182113
rect 217715 182085 217749 182113
rect 217777 182085 217811 182113
rect 217839 182085 217887 182113
rect 217577 182051 217887 182085
rect 217577 182023 217625 182051
rect 217653 182023 217687 182051
rect 217715 182023 217749 182051
rect 217777 182023 217811 182051
rect 217839 182023 217887 182051
rect 217577 181989 217887 182023
rect 217577 181961 217625 181989
rect 217653 181961 217687 181989
rect 217715 181961 217749 181989
rect 217777 181961 217811 181989
rect 217839 181961 217887 181989
rect 217577 173175 217887 181961
rect 217577 173147 217625 173175
rect 217653 173147 217687 173175
rect 217715 173147 217749 173175
rect 217777 173147 217811 173175
rect 217839 173147 217887 173175
rect 217577 173113 217887 173147
rect 217577 173085 217625 173113
rect 217653 173085 217687 173113
rect 217715 173085 217749 173113
rect 217777 173085 217811 173113
rect 217839 173085 217887 173113
rect 217577 173051 217887 173085
rect 217577 173023 217625 173051
rect 217653 173023 217687 173051
rect 217715 173023 217749 173051
rect 217777 173023 217811 173051
rect 217839 173023 217887 173051
rect 217577 172989 217887 173023
rect 217577 172961 217625 172989
rect 217653 172961 217687 172989
rect 217715 172961 217749 172989
rect 217777 172961 217811 172989
rect 217839 172961 217887 172989
rect 217577 164175 217887 172961
rect 217577 164147 217625 164175
rect 217653 164147 217687 164175
rect 217715 164147 217749 164175
rect 217777 164147 217811 164175
rect 217839 164147 217887 164175
rect 217577 164113 217887 164147
rect 217577 164085 217625 164113
rect 217653 164085 217687 164113
rect 217715 164085 217749 164113
rect 217777 164085 217811 164113
rect 217839 164085 217887 164113
rect 217577 164051 217887 164085
rect 217577 164023 217625 164051
rect 217653 164023 217687 164051
rect 217715 164023 217749 164051
rect 217777 164023 217811 164051
rect 217839 164023 217887 164051
rect 217577 163989 217887 164023
rect 217577 163961 217625 163989
rect 217653 163961 217687 163989
rect 217715 163961 217749 163989
rect 217777 163961 217811 163989
rect 217839 163961 217887 163989
rect 217577 155175 217887 163961
rect 217577 155147 217625 155175
rect 217653 155147 217687 155175
rect 217715 155147 217749 155175
rect 217777 155147 217811 155175
rect 217839 155147 217887 155175
rect 217577 155113 217887 155147
rect 217577 155085 217625 155113
rect 217653 155085 217687 155113
rect 217715 155085 217749 155113
rect 217777 155085 217811 155113
rect 217839 155085 217887 155113
rect 217577 155051 217887 155085
rect 217577 155023 217625 155051
rect 217653 155023 217687 155051
rect 217715 155023 217749 155051
rect 217777 155023 217811 155051
rect 217839 155023 217887 155051
rect 217577 154989 217887 155023
rect 217577 154961 217625 154989
rect 217653 154961 217687 154989
rect 217715 154961 217749 154989
rect 217777 154961 217811 154989
rect 217839 154961 217887 154989
rect 217577 146175 217887 154961
rect 217577 146147 217625 146175
rect 217653 146147 217687 146175
rect 217715 146147 217749 146175
rect 217777 146147 217811 146175
rect 217839 146147 217887 146175
rect 217577 146113 217887 146147
rect 217577 146085 217625 146113
rect 217653 146085 217687 146113
rect 217715 146085 217749 146113
rect 217777 146085 217811 146113
rect 217839 146085 217887 146113
rect 217577 146051 217887 146085
rect 217577 146023 217625 146051
rect 217653 146023 217687 146051
rect 217715 146023 217749 146051
rect 217777 146023 217811 146051
rect 217839 146023 217887 146051
rect 217577 145989 217887 146023
rect 217577 145961 217625 145989
rect 217653 145961 217687 145989
rect 217715 145961 217749 145989
rect 217777 145961 217811 145989
rect 217839 145961 217887 145989
rect 217577 137175 217887 145961
rect 217577 137147 217625 137175
rect 217653 137147 217687 137175
rect 217715 137147 217749 137175
rect 217777 137147 217811 137175
rect 217839 137147 217887 137175
rect 217577 137113 217887 137147
rect 217577 137085 217625 137113
rect 217653 137085 217687 137113
rect 217715 137085 217749 137113
rect 217777 137085 217811 137113
rect 217839 137085 217887 137113
rect 217577 137051 217887 137085
rect 217577 137023 217625 137051
rect 217653 137023 217687 137051
rect 217715 137023 217749 137051
rect 217777 137023 217811 137051
rect 217839 137023 217887 137051
rect 217577 136989 217887 137023
rect 217577 136961 217625 136989
rect 217653 136961 217687 136989
rect 217715 136961 217749 136989
rect 217777 136961 217811 136989
rect 217839 136961 217887 136989
rect 217577 128175 217887 136961
rect 217577 128147 217625 128175
rect 217653 128147 217687 128175
rect 217715 128147 217749 128175
rect 217777 128147 217811 128175
rect 217839 128147 217887 128175
rect 217577 128113 217887 128147
rect 217577 128085 217625 128113
rect 217653 128085 217687 128113
rect 217715 128085 217749 128113
rect 217777 128085 217811 128113
rect 217839 128085 217887 128113
rect 217577 128051 217887 128085
rect 217577 128023 217625 128051
rect 217653 128023 217687 128051
rect 217715 128023 217749 128051
rect 217777 128023 217811 128051
rect 217839 128023 217887 128051
rect 217577 127989 217887 128023
rect 217577 127961 217625 127989
rect 217653 127961 217687 127989
rect 217715 127961 217749 127989
rect 217777 127961 217811 127989
rect 217839 127961 217887 127989
rect 217577 119175 217887 127961
rect 217577 119147 217625 119175
rect 217653 119147 217687 119175
rect 217715 119147 217749 119175
rect 217777 119147 217811 119175
rect 217839 119147 217887 119175
rect 217577 119113 217887 119147
rect 217577 119085 217625 119113
rect 217653 119085 217687 119113
rect 217715 119085 217749 119113
rect 217777 119085 217811 119113
rect 217839 119085 217887 119113
rect 217577 119051 217887 119085
rect 217577 119023 217625 119051
rect 217653 119023 217687 119051
rect 217715 119023 217749 119051
rect 217777 119023 217811 119051
rect 217839 119023 217887 119051
rect 217577 118989 217887 119023
rect 217577 118961 217625 118989
rect 217653 118961 217687 118989
rect 217715 118961 217749 118989
rect 217777 118961 217811 118989
rect 217839 118961 217887 118989
rect 217577 110175 217887 118961
rect 217577 110147 217625 110175
rect 217653 110147 217687 110175
rect 217715 110147 217749 110175
rect 217777 110147 217811 110175
rect 217839 110147 217887 110175
rect 217577 110113 217887 110147
rect 217577 110085 217625 110113
rect 217653 110085 217687 110113
rect 217715 110085 217749 110113
rect 217777 110085 217811 110113
rect 217839 110085 217887 110113
rect 217577 110051 217887 110085
rect 217577 110023 217625 110051
rect 217653 110023 217687 110051
rect 217715 110023 217749 110051
rect 217777 110023 217811 110051
rect 217839 110023 217887 110051
rect 217577 109989 217887 110023
rect 217577 109961 217625 109989
rect 217653 109961 217687 109989
rect 217715 109961 217749 109989
rect 217777 109961 217811 109989
rect 217839 109961 217887 109989
rect 217577 101175 217887 109961
rect 217577 101147 217625 101175
rect 217653 101147 217687 101175
rect 217715 101147 217749 101175
rect 217777 101147 217811 101175
rect 217839 101147 217887 101175
rect 217577 101113 217887 101147
rect 217577 101085 217625 101113
rect 217653 101085 217687 101113
rect 217715 101085 217749 101113
rect 217777 101085 217811 101113
rect 217839 101085 217887 101113
rect 217577 101051 217887 101085
rect 217577 101023 217625 101051
rect 217653 101023 217687 101051
rect 217715 101023 217749 101051
rect 217777 101023 217811 101051
rect 217839 101023 217887 101051
rect 217577 100989 217887 101023
rect 217577 100961 217625 100989
rect 217653 100961 217687 100989
rect 217715 100961 217749 100989
rect 217777 100961 217811 100989
rect 217839 100961 217887 100989
rect 217577 92175 217887 100961
rect 217577 92147 217625 92175
rect 217653 92147 217687 92175
rect 217715 92147 217749 92175
rect 217777 92147 217811 92175
rect 217839 92147 217887 92175
rect 217577 92113 217887 92147
rect 217577 92085 217625 92113
rect 217653 92085 217687 92113
rect 217715 92085 217749 92113
rect 217777 92085 217811 92113
rect 217839 92085 217887 92113
rect 217577 92051 217887 92085
rect 217577 92023 217625 92051
rect 217653 92023 217687 92051
rect 217715 92023 217749 92051
rect 217777 92023 217811 92051
rect 217839 92023 217887 92051
rect 217577 91989 217887 92023
rect 217577 91961 217625 91989
rect 217653 91961 217687 91989
rect 217715 91961 217749 91989
rect 217777 91961 217811 91989
rect 217839 91961 217887 91989
rect 217577 83175 217887 91961
rect 217577 83147 217625 83175
rect 217653 83147 217687 83175
rect 217715 83147 217749 83175
rect 217777 83147 217811 83175
rect 217839 83147 217887 83175
rect 217577 83113 217887 83147
rect 217577 83085 217625 83113
rect 217653 83085 217687 83113
rect 217715 83085 217749 83113
rect 217777 83085 217811 83113
rect 217839 83085 217887 83113
rect 217577 83051 217887 83085
rect 217577 83023 217625 83051
rect 217653 83023 217687 83051
rect 217715 83023 217749 83051
rect 217777 83023 217811 83051
rect 217839 83023 217887 83051
rect 217577 82989 217887 83023
rect 217577 82961 217625 82989
rect 217653 82961 217687 82989
rect 217715 82961 217749 82989
rect 217777 82961 217811 82989
rect 217839 82961 217887 82989
rect 217577 74175 217887 82961
rect 217577 74147 217625 74175
rect 217653 74147 217687 74175
rect 217715 74147 217749 74175
rect 217777 74147 217811 74175
rect 217839 74147 217887 74175
rect 217577 74113 217887 74147
rect 217577 74085 217625 74113
rect 217653 74085 217687 74113
rect 217715 74085 217749 74113
rect 217777 74085 217811 74113
rect 217839 74085 217887 74113
rect 217577 74051 217887 74085
rect 217577 74023 217625 74051
rect 217653 74023 217687 74051
rect 217715 74023 217749 74051
rect 217777 74023 217811 74051
rect 217839 74023 217887 74051
rect 217577 73989 217887 74023
rect 217577 73961 217625 73989
rect 217653 73961 217687 73989
rect 217715 73961 217749 73989
rect 217777 73961 217811 73989
rect 217839 73961 217887 73989
rect 217577 65175 217887 73961
rect 217577 65147 217625 65175
rect 217653 65147 217687 65175
rect 217715 65147 217749 65175
rect 217777 65147 217811 65175
rect 217839 65147 217887 65175
rect 217577 65113 217887 65147
rect 217577 65085 217625 65113
rect 217653 65085 217687 65113
rect 217715 65085 217749 65113
rect 217777 65085 217811 65113
rect 217839 65085 217887 65113
rect 217577 65051 217887 65085
rect 217577 65023 217625 65051
rect 217653 65023 217687 65051
rect 217715 65023 217749 65051
rect 217777 65023 217811 65051
rect 217839 65023 217887 65051
rect 217577 64989 217887 65023
rect 217577 64961 217625 64989
rect 217653 64961 217687 64989
rect 217715 64961 217749 64989
rect 217777 64961 217811 64989
rect 217839 64961 217887 64989
rect 217577 56175 217887 64961
rect 217577 56147 217625 56175
rect 217653 56147 217687 56175
rect 217715 56147 217749 56175
rect 217777 56147 217811 56175
rect 217839 56147 217887 56175
rect 217577 56113 217887 56147
rect 217577 56085 217625 56113
rect 217653 56085 217687 56113
rect 217715 56085 217749 56113
rect 217777 56085 217811 56113
rect 217839 56085 217887 56113
rect 217577 56051 217887 56085
rect 217577 56023 217625 56051
rect 217653 56023 217687 56051
rect 217715 56023 217749 56051
rect 217777 56023 217811 56051
rect 217839 56023 217887 56051
rect 217577 55989 217887 56023
rect 217577 55961 217625 55989
rect 217653 55961 217687 55989
rect 217715 55961 217749 55989
rect 217777 55961 217811 55989
rect 217839 55961 217887 55989
rect 217577 47175 217887 55961
rect 217577 47147 217625 47175
rect 217653 47147 217687 47175
rect 217715 47147 217749 47175
rect 217777 47147 217811 47175
rect 217839 47147 217887 47175
rect 217577 47113 217887 47147
rect 217577 47085 217625 47113
rect 217653 47085 217687 47113
rect 217715 47085 217749 47113
rect 217777 47085 217811 47113
rect 217839 47085 217887 47113
rect 217577 47051 217887 47085
rect 217577 47023 217625 47051
rect 217653 47023 217687 47051
rect 217715 47023 217749 47051
rect 217777 47023 217811 47051
rect 217839 47023 217887 47051
rect 217577 46989 217887 47023
rect 217577 46961 217625 46989
rect 217653 46961 217687 46989
rect 217715 46961 217749 46989
rect 217777 46961 217811 46989
rect 217839 46961 217887 46989
rect 217577 38175 217887 46961
rect 217577 38147 217625 38175
rect 217653 38147 217687 38175
rect 217715 38147 217749 38175
rect 217777 38147 217811 38175
rect 217839 38147 217887 38175
rect 217577 38113 217887 38147
rect 217577 38085 217625 38113
rect 217653 38085 217687 38113
rect 217715 38085 217749 38113
rect 217777 38085 217811 38113
rect 217839 38085 217887 38113
rect 217577 38051 217887 38085
rect 217577 38023 217625 38051
rect 217653 38023 217687 38051
rect 217715 38023 217749 38051
rect 217777 38023 217811 38051
rect 217839 38023 217887 38051
rect 217577 37989 217887 38023
rect 217577 37961 217625 37989
rect 217653 37961 217687 37989
rect 217715 37961 217749 37989
rect 217777 37961 217811 37989
rect 217839 37961 217887 37989
rect 217577 29175 217887 37961
rect 217577 29147 217625 29175
rect 217653 29147 217687 29175
rect 217715 29147 217749 29175
rect 217777 29147 217811 29175
rect 217839 29147 217887 29175
rect 217577 29113 217887 29147
rect 217577 29085 217625 29113
rect 217653 29085 217687 29113
rect 217715 29085 217749 29113
rect 217777 29085 217811 29113
rect 217839 29085 217887 29113
rect 217577 29051 217887 29085
rect 217577 29023 217625 29051
rect 217653 29023 217687 29051
rect 217715 29023 217749 29051
rect 217777 29023 217811 29051
rect 217839 29023 217887 29051
rect 217577 28989 217887 29023
rect 217577 28961 217625 28989
rect 217653 28961 217687 28989
rect 217715 28961 217749 28989
rect 217777 28961 217811 28989
rect 217839 28961 217887 28989
rect 217577 20175 217887 28961
rect 217577 20147 217625 20175
rect 217653 20147 217687 20175
rect 217715 20147 217749 20175
rect 217777 20147 217811 20175
rect 217839 20147 217887 20175
rect 217577 20113 217887 20147
rect 217577 20085 217625 20113
rect 217653 20085 217687 20113
rect 217715 20085 217749 20113
rect 217777 20085 217811 20113
rect 217839 20085 217887 20113
rect 217577 20051 217887 20085
rect 217577 20023 217625 20051
rect 217653 20023 217687 20051
rect 217715 20023 217749 20051
rect 217777 20023 217811 20051
rect 217839 20023 217887 20051
rect 217577 19989 217887 20023
rect 217577 19961 217625 19989
rect 217653 19961 217687 19989
rect 217715 19961 217749 19989
rect 217777 19961 217811 19989
rect 217839 19961 217887 19989
rect 217577 11175 217887 19961
rect 217577 11147 217625 11175
rect 217653 11147 217687 11175
rect 217715 11147 217749 11175
rect 217777 11147 217811 11175
rect 217839 11147 217887 11175
rect 217577 11113 217887 11147
rect 217577 11085 217625 11113
rect 217653 11085 217687 11113
rect 217715 11085 217749 11113
rect 217777 11085 217811 11113
rect 217839 11085 217887 11113
rect 217577 11051 217887 11085
rect 217577 11023 217625 11051
rect 217653 11023 217687 11051
rect 217715 11023 217749 11051
rect 217777 11023 217811 11051
rect 217839 11023 217887 11051
rect 217577 10989 217887 11023
rect 217577 10961 217625 10989
rect 217653 10961 217687 10989
rect 217715 10961 217749 10989
rect 217777 10961 217811 10989
rect 217839 10961 217887 10989
rect 217577 2175 217887 10961
rect 217577 2147 217625 2175
rect 217653 2147 217687 2175
rect 217715 2147 217749 2175
rect 217777 2147 217811 2175
rect 217839 2147 217887 2175
rect 217577 2113 217887 2147
rect 217577 2085 217625 2113
rect 217653 2085 217687 2113
rect 217715 2085 217749 2113
rect 217777 2085 217811 2113
rect 217839 2085 217887 2113
rect 217577 2051 217887 2085
rect 217577 2023 217625 2051
rect 217653 2023 217687 2051
rect 217715 2023 217749 2051
rect 217777 2023 217811 2051
rect 217839 2023 217887 2051
rect 217577 1989 217887 2023
rect 217577 1961 217625 1989
rect 217653 1961 217687 1989
rect 217715 1961 217749 1989
rect 217777 1961 217811 1989
rect 217839 1961 217887 1989
rect 217577 -80 217887 1961
rect 217577 -108 217625 -80
rect 217653 -108 217687 -80
rect 217715 -108 217749 -80
rect 217777 -108 217811 -80
rect 217839 -108 217887 -80
rect 217577 -142 217887 -108
rect 217577 -170 217625 -142
rect 217653 -170 217687 -142
rect 217715 -170 217749 -142
rect 217777 -170 217811 -142
rect 217839 -170 217887 -142
rect 217577 -204 217887 -170
rect 217577 -232 217625 -204
rect 217653 -232 217687 -204
rect 217715 -232 217749 -204
rect 217777 -232 217811 -204
rect 217839 -232 217887 -204
rect 217577 -266 217887 -232
rect 217577 -294 217625 -266
rect 217653 -294 217687 -266
rect 217715 -294 217749 -266
rect 217777 -294 217811 -266
rect 217839 -294 217887 -266
rect 217577 -822 217887 -294
rect 219437 299086 219747 299134
rect 219437 299058 219485 299086
rect 219513 299058 219547 299086
rect 219575 299058 219609 299086
rect 219637 299058 219671 299086
rect 219699 299058 219747 299086
rect 219437 299024 219747 299058
rect 219437 298996 219485 299024
rect 219513 298996 219547 299024
rect 219575 298996 219609 299024
rect 219637 298996 219671 299024
rect 219699 298996 219747 299024
rect 219437 298962 219747 298996
rect 219437 298934 219485 298962
rect 219513 298934 219547 298962
rect 219575 298934 219609 298962
rect 219637 298934 219671 298962
rect 219699 298934 219747 298962
rect 219437 298900 219747 298934
rect 219437 298872 219485 298900
rect 219513 298872 219547 298900
rect 219575 298872 219609 298900
rect 219637 298872 219671 298900
rect 219699 298872 219747 298900
rect 219437 293175 219747 298872
rect 219437 293147 219485 293175
rect 219513 293147 219547 293175
rect 219575 293147 219609 293175
rect 219637 293147 219671 293175
rect 219699 293147 219747 293175
rect 219437 293113 219747 293147
rect 219437 293085 219485 293113
rect 219513 293085 219547 293113
rect 219575 293085 219609 293113
rect 219637 293085 219671 293113
rect 219699 293085 219747 293113
rect 219437 293051 219747 293085
rect 219437 293023 219485 293051
rect 219513 293023 219547 293051
rect 219575 293023 219609 293051
rect 219637 293023 219671 293051
rect 219699 293023 219747 293051
rect 219437 292989 219747 293023
rect 219437 292961 219485 292989
rect 219513 292961 219547 292989
rect 219575 292961 219609 292989
rect 219637 292961 219671 292989
rect 219699 292961 219747 292989
rect 219437 284175 219747 292961
rect 219437 284147 219485 284175
rect 219513 284147 219547 284175
rect 219575 284147 219609 284175
rect 219637 284147 219671 284175
rect 219699 284147 219747 284175
rect 219437 284113 219747 284147
rect 219437 284085 219485 284113
rect 219513 284085 219547 284113
rect 219575 284085 219609 284113
rect 219637 284085 219671 284113
rect 219699 284085 219747 284113
rect 219437 284051 219747 284085
rect 219437 284023 219485 284051
rect 219513 284023 219547 284051
rect 219575 284023 219609 284051
rect 219637 284023 219671 284051
rect 219699 284023 219747 284051
rect 219437 283989 219747 284023
rect 219437 283961 219485 283989
rect 219513 283961 219547 283989
rect 219575 283961 219609 283989
rect 219637 283961 219671 283989
rect 219699 283961 219747 283989
rect 219437 275175 219747 283961
rect 219437 275147 219485 275175
rect 219513 275147 219547 275175
rect 219575 275147 219609 275175
rect 219637 275147 219671 275175
rect 219699 275147 219747 275175
rect 219437 275113 219747 275147
rect 219437 275085 219485 275113
rect 219513 275085 219547 275113
rect 219575 275085 219609 275113
rect 219637 275085 219671 275113
rect 219699 275085 219747 275113
rect 219437 275051 219747 275085
rect 219437 275023 219485 275051
rect 219513 275023 219547 275051
rect 219575 275023 219609 275051
rect 219637 275023 219671 275051
rect 219699 275023 219747 275051
rect 219437 274989 219747 275023
rect 219437 274961 219485 274989
rect 219513 274961 219547 274989
rect 219575 274961 219609 274989
rect 219637 274961 219671 274989
rect 219699 274961 219747 274989
rect 219437 266175 219747 274961
rect 219437 266147 219485 266175
rect 219513 266147 219547 266175
rect 219575 266147 219609 266175
rect 219637 266147 219671 266175
rect 219699 266147 219747 266175
rect 219437 266113 219747 266147
rect 219437 266085 219485 266113
rect 219513 266085 219547 266113
rect 219575 266085 219609 266113
rect 219637 266085 219671 266113
rect 219699 266085 219747 266113
rect 219437 266051 219747 266085
rect 219437 266023 219485 266051
rect 219513 266023 219547 266051
rect 219575 266023 219609 266051
rect 219637 266023 219671 266051
rect 219699 266023 219747 266051
rect 219437 265989 219747 266023
rect 219437 265961 219485 265989
rect 219513 265961 219547 265989
rect 219575 265961 219609 265989
rect 219637 265961 219671 265989
rect 219699 265961 219747 265989
rect 219437 257175 219747 265961
rect 219437 257147 219485 257175
rect 219513 257147 219547 257175
rect 219575 257147 219609 257175
rect 219637 257147 219671 257175
rect 219699 257147 219747 257175
rect 219437 257113 219747 257147
rect 219437 257085 219485 257113
rect 219513 257085 219547 257113
rect 219575 257085 219609 257113
rect 219637 257085 219671 257113
rect 219699 257085 219747 257113
rect 219437 257051 219747 257085
rect 219437 257023 219485 257051
rect 219513 257023 219547 257051
rect 219575 257023 219609 257051
rect 219637 257023 219671 257051
rect 219699 257023 219747 257051
rect 219437 256989 219747 257023
rect 219437 256961 219485 256989
rect 219513 256961 219547 256989
rect 219575 256961 219609 256989
rect 219637 256961 219671 256989
rect 219699 256961 219747 256989
rect 219437 248175 219747 256961
rect 219437 248147 219485 248175
rect 219513 248147 219547 248175
rect 219575 248147 219609 248175
rect 219637 248147 219671 248175
rect 219699 248147 219747 248175
rect 219437 248113 219747 248147
rect 219437 248085 219485 248113
rect 219513 248085 219547 248113
rect 219575 248085 219609 248113
rect 219637 248085 219671 248113
rect 219699 248085 219747 248113
rect 219437 248051 219747 248085
rect 219437 248023 219485 248051
rect 219513 248023 219547 248051
rect 219575 248023 219609 248051
rect 219637 248023 219671 248051
rect 219699 248023 219747 248051
rect 219437 247989 219747 248023
rect 219437 247961 219485 247989
rect 219513 247961 219547 247989
rect 219575 247961 219609 247989
rect 219637 247961 219671 247989
rect 219699 247961 219747 247989
rect 219437 239175 219747 247961
rect 219437 239147 219485 239175
rect 219513 239147 219547 239175
rect 219575 239147 219609 239175
rect 219637 239147 219671 239175
rect 219699 239147 219747 239175
rect 219437 239113 219747 239147
rect 219437 239085 219485 239113
rect 219513 239085 219547 239113
rect 219575 239085 219609 239113
rect 219637 239085 219671 239113
rect 219699 239085 219747 239113
rect 219437 239051 219747 239085
rect 219437 239023 219485 239051
rect 219513 239023 219547 239051
rect 219575 239023 219609 239051
rect 219637 239023 219671 239051
rect 219699 239023 219747 239051
rect 219437 238989 219747 239023
rect 219437 238961 219485 238989
rect 219513 238961 219547 238989
rect 219575 238961 219609 238989
rect 219637 238961 219671 238989
rect 219699 238961 219747 238989
rect 219437 230175 219747 238961
rect 219437 230147 219485 230175
rect 219513 230147 219547 230175
rect 219575 230147 219609 230175
rect 219637 230147 219671 230175
rect 219699 230147 219747 230175
rect 219437 230113 219747 230147
rect 219437 230085 219485 230113
rect 219513 230085 219547 230113
rect 219575 230085 219609 230113
rect 219637 230085 219671 230113
rect 219699 230085 219747 230113
rect 219437 230051 219747 230085
rect 219437 230023 219485 230051
rect 219513 230023 219547 230051
rect 219575 230023 219609 230051
rect 219637 230023 219671 230051
rect 219699 230023 219747 230051
rect 219437 229989 219747 230023
rect 219437 229961 219485 229989
rect 219513 229961 219547 229989
rect 219575 229961 219609 229989
rect 219637 229961 219671 229989
rect 219699 229961 219747 229989
rect 219437 221175 219747 229961
rect 219437 221147 219485 221175
rect 219513 221147 219547 221175
rect 219575 221147 219609 221175
rect 219637 221147 219671 221175
rect 219699 221147 219747 221175
rect 219437 221113 219747 221147
rect 219437 221085 219485 221113
rect 219513 221085 219547 221113
rect 219575 221085 219609 221113
rect 219637 221085 219671 221113
rect 219699 221085 219747 221113
rect 219437 221051 219747 221085
rect 219437 221023 219485 221051
rect 219513 221023 219547 221051
rect 219575 221023 219609 221051
rect 219637 221023 219671 221051
rect 219699 221023 219747 221051
rect 219437 220989 219747 221023
rect 219437 220961 219485 220989
rect 219513 220961 219547 220989
rect 219575 220961 219609 220989
rect 219637 220961 219671 220989
rect 219699 220961 219747 220989
rect 219437 212175 219747 220961
rect 219437 212147 219485 212175
rect 219513 212147 219547 212175
rect 219575 212147 219609 212175
rect 219637 212147 219671 212175
rect 219699 212147 219747 212175
rect 219437 212113 219747 212147
rect 219437 212085 219485 212113
rect 219513 212085 219547 212113
rect 219575 212085 219609 212113
rect 219637 212085 219671 212113
rect 219699 212085 219747 212113
rect 219437 212051 219747 212085
rect 219437 212023 219485 212051
rect 219513 212023 219547 212051
rect 219575 212023 219609 212051
rect 219637 212023 219671 212051
rect 219699 212023 219747 212051
rect 219437 211989 219747 212023
rect 219437 211961 219485 211989
rect 219513 211961 219547 211989
rect 219575 211961 219609 211989
rect 219637 211961 219671 211989
rect 219699 211961 219747 211989
rect 219437 203175 219747 211961
rect 219437 203147 219485 203175
rect 219513 203147 219547 203175
rect 219575 203147 219609 203175
rect 219637 203147 219671 203175
rect 219699 203147 219747 203175
rect 219437 203113 219747 203147
rect 219437 203085 219485 203113
rect 219513 203085 219547 203113
rect 219575 203085 219609 203113
rect 219637 203085 219671 203113
rect 219699 203085 219747 203113
rect 219437 203051 219747 203085
rect 219437 203023 219485 203051
rect 219513 203023 219547 203051
rect 219575 203023 219609 203051
rect 219637 203023 219671 203051
rect 219699 203023 219747 203051
rect 219437 202989 219747 203023
rect 219437 202961 219485 202989
rect 219513 202961 219547 202989
rect 219575 202961 219609 202989
rect 219637 202961 219671 202989
rect 219699 202961 219747 202989
rect 219437 194175 219747 202961
rect 219437 194147 219485 194175
rect 219513 194147 219547 194175
rect 219575 194147 219609 194175
rect 219637 194147 219671 194175
rect 219699 194147 219747 194175
rect 219437 194113 219747 194147
rect 219437 194085 219485 194113
rect 219513 194085 219547 194113
rect 219575 194085 219609 194113
rect 219637 194085 219671 194113
rect 219699 194085 219747 194113
rect 219437 194051 219747 194085
rect 219437 194023 219485 194051
rect 219513 194023 219547 194051
rect 219575 194023 219609 194051
rect 219637 194023 219671 194051
rect 219699 194023 219747 194051
rect 219437 193989 219747 194023
rect 219437 193961 219485 193989
rect 219513 193961 219547 193989
rect 219575 193961 219609 193989
rect 219637 193961 219671 193989
rect 219699 193961 219747 193989
rect 219437 185175 219747 193961
rect 219437 185147 219485 185175
rect 219513 185147 219547 185175
rect 219575 185147 219609 185175
rect 219637 185147 219671 185175
rect 219699 185147 219747 185175
rect 219437 185113 219747 185147
rect 219437 185085 219485 185113
rect 219513 185085 219547 185113
rect 219575 185085 219609 185113
rect 219637 185085 219671 185113
rect 219699 185085 219747 185113
rect 219437 185051 219747 185085
rect 219437 185023 219485 185051
rect 219513 185023 219547 185051
rect 219575 185023 219609 185051
rect 219637 185023 219671 185051
rect 219699 185023 219747 185051
rect 219437 184989 219747 185023
rect 219437 184961 219485 184989
rect 219513 184961 219547 184989
rect 219575 184961 219609 184989
rect 219637 184961 219671 184989
rect 219699 184961 219747 184989
rect 219437 176175 219747 184961
rect 219437 176147 219485 176175
rect 219513 176147 219547 176175
rect 219575 176147 219609 176175
rect 219637 176147 219671 176175
rect 219699 176147 219747 176175
rect 219437 176113 219747 176147
rect 219437 176085 219485 176113
rect 219513 176085 219547 176113
rect 219575 176085 219609 176113
rect 219637 176085 219671 176113
rect 219699 176085 219747 176113
rect 219437 176051 219747 176085
rect 219437 176023 219485 176051
rect 219513 176023 219547 176051
rect 219575 176023 219609 176051
rect 219637 176023 219671 176051
rect 219699 176023 219747 176051
rect 219437 175989 219747 176023
rect 219437 175961 219485 175989
rect 219513 175961 219547 175989
rect 219575 175961 219609 175989
rect 219637 175961 219671 175989
rect 219699 175961 219747 175989
rect 219437 167175 219747 175961
rect 219437 167147 219485 167175
rect 219513 167147 219547 167175
rect 219575 167147 219609 167175
rect 219637 167147 219671 167175
rect 219699 167147 219747 167175
rect 219437 167113 219747 167147
rect 219437 167085 219485 167113
rect 219513 167085 219547 167113
rect 219575 167085 219609 167113
rect 219637 167085 219671 167113
rect 219699 167085 219747 167113
rect 219437 167051 219747 167085
rect 219437 167023 219485 167051
rect 219513 167023 219547 167051
rect 219575 167023 219609 167051
rect 219637 167023 219671 167051
rect 219699 167023 219747 167051
rect 219437 166989 219747 167023
rect 219437 166961 219485 166989
rect 219513 166961 219547 166989
rect 219575 166961 219609 166989
rect 219637 166961 219671 166989
rect 219699 166961 219747 166989
rect 219437 158175 219747 166961
rect 219437 158147 219485 158175
rect 219513 158147 219547 158175
rect 219575 158147 219609 158175
rect 219637 158147 219671 158175
rect 219699 158147 219747 158175
rect 219437 158113 219747 158147
rect 219437 158085 219485 158113
rect 219513 158085 219547 158113
rect 219575 158085 219609 158113
rect 219637 158085 219671 158113
rect 219699 158085 219747 158113
rect 219437 158051 219747 158085
rect 219437 158023 219485 158051
rect 219513 158023 219547 158051
rect 219575 158023 219609 158051
rect 219637 158023 219671 158051
rect 219699 158023 219747 158051
rect 219437 157989 219747 158023
rect 219437 157961 219485 157989
rect 219513 157961 219547 157989
rect 219575 157961 219609 157989
rect 219637 157961 219671 157989
rect 219699 157961 219747 157989
rect 219437 149175 219747 157961
rect 219437 149147 219485 149175
rect 219513 149147 219547 149175
rect 219575 149147 219609 149175
rect 219637 149147 219671 149175
rect 219699 149147 219747 149175
rect 219437 149113 219747 149147
rect 219437 149085 219485 149113
rect 219513 149085 219547 149113
rect 219575 149085 219609 149113
rect 219637 149085 219671 149113
rect 219699 149085 219747 149113
rect 219437 149051 219747 149085
rect 219437 149023 219485 149051
rect 219513 149023 219547 149051
rect 219575 149023 219609 149051
rect 219637 149023 219671 149051
rect 219699 149023 219747 149051
rect 219437 148989 219747 149023
rect 219437 148961 219485 148989
rect 219513 148961 219547 148989
rect 219575 148961 219609 148989
rect 219637 148961 219671 148989
rect 219699 148961 219747 148989
rect 219437 140175 219747 148961
rect 219437 140147 219485 140175
rect 219513 140147 219547 140175
rect 219575 140147 219609 140175
rect 219637 140147 219671 140175
rect 219699 140147 219747 140175
rect 219437 140113 219747 140147
rect 219437 140085 219485 140113
rect 219513 140085 219547 140113
rect 219575 140085 219609 140113
rect 219637 140085 219671 140113
rect 219699 140085 219747 140113
rect 219437 140051 219747 140085
rect 219437 140023 219485 140051
rect 219513 140023 219547 140051
rect 219575 140023 219609 140051
rect 219637 140023 219671 140051
rect 219699 140023 219747 140051
rect 219437 139989 219747 140023
rect 219437 139961 219485 139989
rect 219513 139961 219547 139989
rect 219575 139961 219609 139989
rect 219637 139961 219671 139989
rect 219699 139961 219747 139989
rect 219437 131175 219747 139961
rect 219437 131147 219485 131175
rect 219513 131147 219547 131175
rect 219575 131147 219609 131175
rect 219637 131147 219671 131175
rect 219699 131147 219747 131175
rect 219437 131113 219747 131147
rect 219437 131085 219485 131113
rect 219513 131085 219547 131113
rect 219575 131085 219609 131113
rect 219637 131085 219671 131113
rect 219699 131085 219747 131113
rect 219437 131051 219747 131085
rect 219437 131023 219485 131051
rect 219513 131023 219547 131051
rect 219575 131023 219609 131051
rect 219637 131023 219671 131051
rect 219699 131023 219747 131051
rect 219437 130989 219747 131023
rect 219437 130961 219485 130989
rect 219513 130961 219547 130989
rect 219575 130961 219609 130989
rect 219637 130961 219671 130989
rect 219699 130961 219747 130989
rect 219437 122175 219747 130961
rect 219437 122147 219485 122175
rect 219513 122147 219547 122175
rect 219575 122147 219609 122175
rect 219637 122147 219671 122175
rect 219699 122147 219747 122175
rect 219437 122113 219747 122147
rect 219437 122085 219485 122113
rect 219513 122085 219547 122113
rect 219575 122085 219609 122113
rect 219637 122085 219671 122113
rect 219699 122085 219747 122113
rect 219437 122051 219747 122085
rect 219437 122023 219485 122051
rect 219513 122023 219547 122051
rect 219575 122023 219609 122051
rect 219637 122023 219671 122051
rect 219699 122023 219747 122051
rect 219437 121989 219747 122023
rect 219437 121961 219485 121989
rect 219513 121961 219547 121989
rect 219575 121961 219609 121989
rect 219637 121961 219671 121989
rect 219699 121961 219747 121989
rect 219437 113175 219747 121961
rect 219437 113147 219485 113175
rect 219513 113147 219547 113175
rect 219575 113147 219609 113175
rect 219637 113147 219671 113175
rect 219699 113147 219747 113175
rect 219437 113113 219747 113147
rect 219437 113085 219485 113113
rect 219513 113085 219547 113113
rect 219575 113085 219609 113113
rect 219637 113085 219671 113113
rect 219699 113085 219747 113113
rect 219437 113051 219747 113085
rect 219437 113023 219485 113051
rect 219513 113023 219547 113051
rect 219575 113023 219609 113051
rect 219637 113023 219671 113051
rect 219699 113023 219747 113051
rect 219437 112989 219747 113023
rect 219437 112961 219485 112989
rect 219513 112961 219547 112989
rect 219575 112961 219609 112989
rect 219637 112961 219671 112989
rect 219699 112961 219747 112989
rect 219437 104175 219747 112961
rect 219437 104147 219485 104175
rect 219513 104147 219547 104175
rect 219575 104147 219609 104175
rect 219637 104147 219671 104175
rect 219699 104147 219747 104175
rect 219437 104113 219747 104147
rect 219437 104085 219485 104113
rect 219513 104085 219547 104113
rect 219575 104085 219609 104113
rect 219637 104085 219671 104113
rect 219699 104085 219747 104113
rect 219437 104051 219747 104085
rect 219437 104023 219485 104051
rect 219513 104023 219547 104051
rect 219575 104023 219609 104051
rect 219637 104023 219671 104051
rect 219699 104023 219747 104051
rect 219437 103989 219747 104023
rect 219437 103961 219485 103989
rect 219513 103961 219547 103989
rect 219575 103961 219609 103989
rect 219637 103961 219671 103989
rect 219699 103961 219747 103989
rect 219437 95175 219747 103961
rect 219437 95147 219485 95175
rect 219513 95147 219547 95175
rect 219575 95147 219609 95175
rect 219637 95147 219671 95175
rect 219699 95147 219747 95175
rect 219437 95113 219747 95147
rect 219437 95085 219485 95113
rect 219513 95085 219547 95113
rect 219575 95085 219609 95113
rect 219637 95085 219671 95113
rect 219699 95085 219747 95113
rect 219437 95051 219747 95085
rect 219437 95023 219485 95051
rect 219513 95023 219547 95051
rect 219575 95023 219609 95051
rect 219637 95023 219671 95051
rect 219699 95023 219747 95051
rect 219437 94989 219747 95023
rect 219437 94961 219485 94989
rect 219513 94961 219547 94989
rect 219575 94961 219609 94989
rect 219637 94961 219671 94989
rect 219699 94961 219747 94989
rect 219437 86175 219747 94961
rect 219437 86147 219485 86175
rect 219513 86147 219547 86175
rect 219575 86147 219609 86175
rect 219637 86147 219671 86175
rect 219699 86147 219747 86175
rect 219437 86113 219747 86147
rect 219437 86085 219485 86113
rect 219513 86085 219547 86113
rect 219575 86085 219609 86113
rect 219637 86085 219671 86113
rect 219699 86085 219747 86113
rect 219437 86051 219747 86085
rect 219437 86023 219485 86051
rect 219513 86023 219547 86051
rect 219575 86023 219609 86051
rect 219637 86023 219671 86051
rect 219699 86023 219747 86051
rect 219437 85989 219747 86023
rect 219437 85961 219485 85989
rect 219513 85961 219547 85989
rect 219575 85961 219609 85989
rect 219637 85961 219671 85989
rect 219699 85961 219747 85989
rect 219437 77175 219747 85961
rect 219437 77147 219485 77175
rect 219513 77147 219547 77175
rect 219575 77147 219609 77175
rect 219637 77147 219671 77175
rect 219699 77147 219747 77175
rect 219437 77113 219747 77147
rect 219437 77085 219485 77113
rect 219513 77085 219547 77113
rect 219575 77085 219609 77113
rect 219637 77085 219671 77113
rect 219699 77085 219747 77113
rect 219437 77051 219747 77085
rect 219437 77023 219485 77051
rect 219513 77023 219547 77051
rect 219575 77023 219609 77051
rect 219637 77023 219671 77051
rect 219699 77023 219747 77051
rect 219437 76989 219747 77023
rect 219437 76961 219485 76989
rect 219513 76961 219547 76989
rect 219575 76961 219609 76989
rect 219637 76961 219671 76989
rect 219699 76961 219747 76989
rect 219437 68175 219747 76961
rect 219437 68147 219485 68175
rect 219513 68147 219547 68175
rect 219575 68147 219609 68175
rect 219637 68147 219671 68175
rect 219699 68147 219747 68175
rect 219437 68113 219747 68147
rect 219437 68085 219485 68113
rect 219513 68085 219547 68113
rect 219575 68085 219609 68113
rect 219637 68085 219671 68113
rect 219699 68085 219747 68113
rect 219437 68051 219747 68085
rect 219437 68023 219485 68051
rect 219513 68023 219547 68051
rect 219575 68023 219609 68051
rect 219637 68023 219671 68051
rect 219699 68023 219747 68051
rect 219437 67989 219747 68023
rect 219437 67961 219485 67989
rect 219513 67961 219547 67989
rect 219575 67961 219609 67989
rect 219637 67961 219671 67989
rect 219699 67961 219747 67989
rect 219437 59175 219747 67961
rect 219437 59147 219485 59175
rect 219513 59147 219547 59175
rect 219575 59147 219609 59175
rect 219637 59147 219671 59175
rect 219699 59147 219747 59175
rect 219437 59113 219747 59147
rect 219437 59085 219485 59113
rect 219513 59085 219547 59113
rect 219575 59085 219609 59113
rect 219637 59085 219671 59113
rect 219699 59085 219747 59113
rect 219437 59051 219747 59085
rect 219437 59023 219485 59051
rect 219513 59023 219547 59051
rect 219575 59023 219609 59051
rect 219637 59023 219671 59051
rect 219699 59023 219747 59051
rect 219437 58989 219747 59023
rect 219437 58961 219485 58989
rect 219513 58961 219547 58989
rect 219575 58961 219609 58989
rect 219637 58961 219671 58989
rect 219699 58961 219747 58989
rect 219437 50175 219747 58961
rect 219437 50147 219485 50175
rect 219513 50147 219547 50175
rect 219575 50147 219609 50175
rect 219637 50147 219671 50175
rect 219699 50147 219747 50175
rect 219437 50113 219747 50147
rect 219437 50085 219485 50113
rect 219513 50085 219547 50113
rect 219575 50085 219609 50113
rect 219637 50085 219671 50113
rect 219699 50085 219747 50113
rect 219437 50051 219747 50085
rect 219437 50023 219485 50051
rect 219513 50023 219547 50051
rect 219575 50023 219609 50051
rect 219637 50023 219671 50051
rect 219699 50023 219747 50051
rect 219437 49989 219747 50023
rect 219437 49961 219485 49989
rect 219513 49961 219547 49989
rect 219575 49961 219609 49989
rect 219637 49961 219671 49989
rect 219699 49961 219747 49989
rect 219437 41175 219747 49961
rect 219437 41147 219485 41175
rect 219513 41147 219547 41175
rect 219575 41147 219609 41175
rect 219637 41147 219671 41175
rect 219699 41147 219747 41175
rect 219437 41113 219747 41147
rect 219437 41085 219485 41113
rect 219513 41085 219547 41113
rect 219575 41085 219609 41113
rect 219637 41085 219671 41113
rect 219699 41085 219747 41113
rect 219437 41051 219747 41085
rect 219437 41023 219485 41051
rect 219513 41023 219547 41051
rect 219575 41023 219609 41051
rect 219637 41023 219671 41051
rect 219699 41023 219747 41051
rect 219437 40989 219747 41023
rect 219437 40961 219485 40989
rect 219513 40961 219547 40989
rect 219575 40961 219609 40989
rect 219637 40961 219671 40989
rect 219699 40961 219747 40989
rect 219437 32175 219747 40961
rect 219437 32147 219485 32175
rect 219513 32147 219547 32175
rect 219575 32147 219609 32175
rect 219637 32147 219671 32175
rect 219699 32147 219747 32175
rect 219437 32113 219747 32147
rect 219437 32085 219485 32113
rect 219513 32085 219547 32113
rect 219575 32085 219609 32113
rect 219637 32085 219671 32113
rect 219699 32085 219747 32113
rect 219437 32051 219747 32085
rect 219437 32023 219485 32051
rect 219513 32023 219547 32051
rect 219575 32023 219609 32051
rect 219637 32023 219671 32051
rect 219699 32023 219747 32051
rect 219437 31989 219747 32023
rect 219437 31961 219485 31989
rect 219513 31961 219547 31989
rect 219575 31961 219609 31989
rect 219637 31961 219671 31989
rect 219699 31961 219747 31989
rect 219437 23175 219747 31961
rect 219437 23147 219485 23175
rect 219513 23147 219547 23175
rect 219575 23147 219609 23175
rect 219637 23147 219671 23175
rect 219699 23147 219747 23175
rect 219437 23113 219747 23147
rect 219437 23085 219485 23113
rect 219513 23085 219547 23113
rect 219575 23085 219609 23113
rect 219637 23085 219671 23113
rect 219699 23085 219747 23113
rect 219437 23051 219747 23085
rect 219437 23023 219485 23051
rect 219513 23023 219547 23051
rect 219575 23023 219609 23051
rect 219637 23023 219671 23051
rect 219699 23023 219747 23051
rect 219437 22989 219747 23023
rect 219437 22961 219485 22989
rect 219513 22961 219547 22989
rect 219575 22961 219609 22989
rect 219637 22961 219671 22989
rect 219699 22961 219747 22989
rect 219437 14175 219747 22961
rect 219437 14147 219485 14175
rect 219513 14147 219547 14175
rect 219575 14147 219609 14175
rect 219637 14147 219671 14175
rect 219699 14147 219747 14175
rect 219437 14113 219747 14147
rect 219437 14085 219485 14113
rect 219513 14085 219547 14113
rect 219575 14085 219609 14113
rect 219637 14085 219671 14113
rect 219699 14085 219747 14113
rect 219437 14051 219747 14085
rect 219437 14023 219485 14051
rect 219513 14023 219547 14051
rect 219575 14023 219609 14051
rect 219637 14023 219671 14051
rect 219699 14023 219747 14051
rect 219437 13989 219747 14023
rect 219437 13961 219485 13989
rect 219513 13961 219547 13989
rect 219575 13961 219609 13989
rect 219637 13961 219671 13989
rect 219699 13961 219747 13989
rect 219437 5175 219747 13961
rect 219437 5147 219485 5175
rect 219513 5147 219547 5175
rect 219575 5147 219609 5175
rect 219637 5147 219671 5175
rect 219699 5147 219747 5175
rect 219437 5113 219747 5147
rect 219437 5085 219485 5113
rect 219513 5085 219547 5113
rect 219575 5085 219609 5113
rect 219637 5085 219671 5113
rect 219699 5085 219747 5113
rect 219437 5051 219747 5085
rect 219437 5023 219485 5051
rect 219513 5023 219547 5051
rect 219575 5023 219609 5051
rect 219637 5023 219671 5051
rect 219699 5023 219747 5051
rect 219437 4989 219747 5023
rect 219437 4961 219485 4989
rect 219513 4961 219547 4989
rect 219575 4961 219609 4989
rect 219637 4961 219671 4989
rect 219699 4961 219747 4989
rect 219437 -560 219747 4961
rect 219437 -588 219485 -560
rect 219513 -588 219547 -560
rect 219575 -588 219609 -560
rect 219637 -588 219671 -560
rect 219699 -588 219747 -560
rect 219437 -622 219747 -588
rect 219437 -650 219485 -622
rect 219513 -650 219547 -622
rect 219575 -650 219609 -622
rect 219637 -650 219671 -622
rect 219699 -650 219747 -622
rect 219437 -684 219747 -650
rect 219437 -712 219485 -684
rect 219513 -712 219547 -684
rect 219575 -712 219609 -684
rect 219637 -712 219671 -684
rect 219699 -712 219747 -684
rect 219437 -746 219747 -712
rect 219437 -774 219485 -746
rect 219513 -774 219547 -746
rect 219575 -774 219609 -746
rect 219637 -774 219671 -746
rect 219699 -774 219747 -746
rect 219437 -822 219747 -774
rect 226577 298606 226887 299134
rect 226577 298578 226625 298606
rect 226653 298578 226687 298606
rect 226715 298578 226749 298606
rect 226777 298578 226811 298606
rect 226839 298578 226887 298606
rect 226577 298544 226887 298578
rect 226577 298516 226625 298544
rect 226653 298516 226687 298544
rect 226715 298516 226749 298544
rect 226777 298516 226811 298544
rect 226839 298516 226887 298544
rect 226577 298482 226887 298516
rect 226577 298454 226625 298482
rect 226653 298454 226687 298482
rect 226715 298454 226749 298482
rect 226777 298454 226811 298482
rect 226839 298454 226887 298482
rect 226577 298420 226887 298454
rect 226577 298392 226625 298420
rect 226653 298392 226687 298420
rect 226715 298392 226749 298420
rect 226777 298392 226811 298420
rect 226839 298392 226887 298420
rect 226577 290175 226887 298392
rect 226577 290147 226625 290175
rect 226653 290147 226687 290175
rect 226715 290147 226749 290175
rect 226777 290147 226811 290175
rect 226839 290147 226887 290175
rect 226577 290113 226887 290147
rect 226577 290085 226625 290113
rect 226653 290085 226687 290113
rect 226715 290085 226749 290113
rect 226777 290085 226811 290113
rect 226839 290085 226887 290113
rect 226577 290051 226887 290085
rect 226577 290023 226625 290051
rect 226653 290023 226687 290051
rect 226715 290023 226749 290051
rect 226777 290023 226811 290051
rect 226839 290023 226887 290051
rect 226577 289989 226887 290023
rect 226577 289961 226625 289989
rect 226653 289961 226687 289989
rect 226715 289961 226749 289989
rect 226777 289961 226811 289989
rect 226839 289961 226887 289989
rect 226577 281175 226887 289961
rect 226577 281147 226625 281175
rect 226653 281147 226687 281175
rect 226715 281147 226749 281175
rect 226777 281147 226811 281175
rect 226839 281147 226887 281175
rect 226577 281113 226887 281147
rect 226577 281085 226625 281113
rect 226653 281085 226687 281113
rect 226715 281085 226749 281113
rect 226777 281085 226811 281113
rect 226839 281085 226887 281113
rect 226577 281051 226887 281085
rect 226577 281023 226625 281051
rect 226653 281023 226687 281051
rect 226715 281023 226749 281051
rect 226777 281023 226811 281051
rect 226839 281023 226887 281051
rect 226577 280989 226887 281023
rect 226577 280961 226625 280989
rect 226653 280961 226687 280989
rect 226715 280961 226749 280989
rect 226777 280961 226811 280989
rect 226839 280961 226887 280989
rect 226577 272175 226887 280961
rect 226577 272147 226625 272175
rect 226653 272147 226687 272175
rect 226715 272147 226749 272175
rect 226777 272147 226811 272175
rect 226839 272147 226887 272175
rect 226577 272113 226887 272147
rect 226577 272085 226625 272113
rect 226653 272085 226687 272113
rect 226715 272085 226749 272113
rect 226777 272085 226811 272113
rect 226839 272085 226887 272113
rect 226577 272051 226887 272085
rect 226577 272023 226625 272051
rect 226653 272023 226687 272051
rect 226715 272023 226749 272051
rect 226777 272023 226811 272051
rect 226839 272023 226887 272051
rect 226577 271989 226887 272023
rect 226577 271961 226625 271989
rect 226653 271961 226687 271989
rect 226715 271961 226749 271989
rect 226777 271961 226811 271989
rect 226839 271961 226887 271989
rect 226577 263175 226887 271961
rect 226577 263147 226625 263175
rect 226653 263147 226687 263175
rect 226715 263147 226749 263175
rect 226777 263147 226811 263175
rect 226839 263147 226887 263175
rect 226577 263113 226887 263147
rect 226577 263085 226625 263113
rect 226653 263085 226687 263113
rect 226715 263085 226749 263113
rect 226777 263085 226811 263113
rect 226839 263085 226887 263113
rect 226577 263051 226887 263085
rect 226577 263023 226625 263051
rect 226653 263023 226687 263051
rect 226715 263023 226749 263051
rect 226777 263023 226811 263051
rect 226839 263023 226887 263051
rect 226577 262989 226887 263023
rect 226577 262961 226625 262989
rect 226653 262961 226687 262989
rect 226715 262961 226749 262989
rect 226777 262961 226811 262989
rect 226839 262961 226887 262989
rect 226577 254175 226887 262961
rect 226577 254147 226625 254175
rect 226653 254147 226687 254175
rect 226715 254147 226749 254175
rect 226777 254147 226811 254175
rect 226839 254147 226887 254175
rect 226577 254113 226887 254147
rect 226577 254085 226625 254113
rect 226653 254085 226687 254113
rect 226715 254085 226749 254113
rect 226777 254085 226811 254113
rect 226839 254085 226887 254113
rect 226577 254051 226887 254085
rect 226577 254023 226625 254051
rect 226653 254023 226687 254051
rect 226715 254023 226749 254051
rect 226777 254023 226811 254051
rect 226839 254023 226887 254051
rect 226577 253989 226887 254023
rect 226577 253961 226625 253989
rect 226653 253961 226687 253989
rect 226715 253961 226749 253989
rect 226777 253961 226811 253989
rect 226839 253961 226887 253989
rect 226577 245175 226887 253961
rect 226577 245147 226625 245175
rect 226653 245147 226687 245175
rect 226715 245147 226749 245175
rect 226777 245147 226811 245175
rect 226839 245147 226887 245175
rect 226577 245113 226887 245147
rect 226577 245085 226625 245113
rect 226653 245085 226687 245113
rect 226715 245085 226749 245113
rect 226777 245085 226811 245113
rect 226839 245085 226887 245113
rect 226577 245051 226887 245085
rect 226577 245023 226625 245051
rect 226653 245023 226687 245051
rect 226715 245023 226749 245051
rect 226777 245023 226811 245051
rect 226839 245023 226887 245051
rect 226577 244989 226887 245023
rect 226577 244961 226625 244989
rect 226653 244961 226687 244989
rect 226715 244961 226749 244989
rect 226777 244961 226811 244989
rect 226839 244961 226887 244989
rect 226577 236175 226887 244961
rect 226577 236147 226625 236175
rect 226653 236147 226687 236175
rect 226715 236147 226749 236175
rect 226777 236147 226811 236175
rect 226839 236147 226887 236175
rect 226577 236113 226887 236147
rect 226577 236085 226625 236113
rect 226653 236085 226687 236113
rect 226715 236085 226749 236113
rect 226777 236085 226811 236113
rect 226839 236085 226887 236113
rect 226577 236051 226887 236085
rect 226577 236023 226625 236051
rect 226653 236023 226687 236051
rect 226715 236023 226749 236051
rect 226777 236023 226811 236051
rect 226839 236023 226887 236051
rect 226577 235989 226887 236023
rect 226577 235961 226625 235989
rect 226653 235961 226687 235989
rect 226715 235961 226749 235989
rect 226777 235961 226811 235989
rect 226839 235961 226887 235989
rect 226577 227175 226887 235961
rect 226577 227147 226625 227175
rect 226653 227147 226687 227175
rect 226715 227147 226749 227175
rect 226777 227147 226811 227175
rect 226839 227147 226887 227175
rect 226577 227113 226887 227147
rect 226577 227085 226625 227113
rect 226653 227085 226687 227113
rect 226715 227085 226749 227113
rect 226777 227085 226811 227113
rect 226839 227085 226887 227113
rect 226577 227051 226887 227085
rect 226577 227023 226625 227051
rect 226653 227023 226687 227051
rect 226715 227023 226749 227051
rect 226777 227023 226811 227051
rect 226839 227023 226887 227051
rect 226577 226989 226887 227023
rect 226577 226961 226625 226989
rect 226653 226961 226687 226989
rect 226715 226961 226749 226989
rect 226777 226961 226811 226989
rect 226839 226961 226887 226989
rect 226577 218175 226887 226961
rect 226577 218147 226625 218175
rect 226653 218147 226687 218175
rect 226715 218147 226749 218175
rect 226777 218147 226811 218175
rect 226839 218147 226887 218175
rect 226577 218113 226887 218147
rect 226577 218085 226625 218113
rect 226653 218085 226687 218113
rect 226715 218085 226749 218113
rect 226777 218085 226811 218113
rect 226839 218085 226887 218113
rect 226577 218051 226887 218085
rect 226577 218023 226625 218051
rect 226653 218023 226687 218051
rect 226715 218023 226749 218051
rect 226777 218023 226811 218051
rect 226839 218023 226887 218051
rect 226577 217989 226887 218023
rect 226577 217961 226625 217989
rect 226653 217961 226687 217989
rect 226715 217961 226749 217989
rect 226777 217961 226811 217989
rect 226839 217961 226887 217989
rect 226577 209175 226887 217961
rect 226577 209147 226625 209175
rect 226653 209147 226687 209175
rect 226715 209147 226749 209175
rect 226777 209147 226811 209175
rect 226839 209147 226887 209175
rect 226577 209113 226887 209147
rect 226577 209085 226625 209113
rect 226653 209085 226687 209113
rect 226715 209085 226749 209113
rect 226777 209085 226811 209113
rect 226839 209085 226887 209113
rect 226577 209051 226887 209085
rect 226577 209023 226625 209051
rect 226653 209023 226687 209051
rect 226715 209023 226749 209051
rect 226777 209023 226811 209051
rect 226839 209023 226887 209051
rect 226577 208989 226887 209023
rect 226577 208961 226625 208989
rect 226653 208961 226687 208989
rect 226715 208961 226749 208989
rect 226777 208961 226811 208989
rect 226839 208961 226887 208989
rect 226577 200175 226887 208961
rect 226577 200147 226625 200175
rect 226653 200147 226687 200175
rect 226715 200147 226749 200175
rect 226777 200147 226811 200175
rect 226839 200147 226887 200175
rect 226577 200113 226887 200147
rect 226577 200085 226625 200113
rect 226653 200085 226687 200113
rect 226715 200085 226749 200113
rect 226777 200085 226811 200113
rect 226839 200085 226887 200113
rect 226577 200051 226887 200085
rect 226577 200023 226625 200051
rect 226653 200023 226687 200051
rect 226715 200023 226749 200051
rect 226777 200023 226811 200051
rect 226839 200023 226887 200051
rect 226577 199989 226887 200023
rect 226577 199961 226625 199989
rect 226653 199961 226687 199989
rect 226715 199961 226749 199989
rect 226777 199961 226811 199989
rect 226839 199961 226887 199989
rect 226577 191175 226887 199961
rect 226577 191147 226625 191175
rect 226653 191147 226687 191175
rect 226715 191147 226749 191175
rect 226777 191147 226811 191175
rect 226839 191147 226887 191175
rect 226577 191113 226887 191147
rect 226577 191085 226625 191113
rect 226653 191085 226687 191113
rect 226715 191085 226749 191113
rect 226777 191085 226811 191113
rect 226839 191085 226887 191113
rect 226577 191051 226887 191085
rect 226577 191023 226625 191051
rect 226653 191023 226687 191051
rect 226715 191023 226749 191051
rect 226777 191023 226811 191051
rect 226839 191023 226887 191051
rect 226577 190989 226887 191023
rect 226577 190961 226625 190989
rect 226653 190961 226687 190989
rect 226715 190961 226749 190989
rect 226777 190961 226811 190989
rect 226839 190961 226887 190989
rect 226577 182175 226887 190961
rect 226577 182147 226625 182175
rect 226653 182147 226687 182175
rect 226715 182147 226749 182175
rect 226777 182147 226811 182175
rect 226839 182147 226887 182175
rect 226577 182113 226887 182147
rect 226577 182085 226625 182113
rect 226653 182085 226687 182113
rect 226715 182085 226749 182113
rect 226777 182085 226811 182113
rect 226839 182085 226887 182113
rect 226577 182051 226887 182085
rect 226577 182023 226625 182051
rect 226653 182023 226687 182051
rect 226715 182023 226749 182051
rect 226777 182023 226811 182051
rect 226839 182023 226887 182051
rect 226577 181989 226887 182023
rect 226577 181961 226625 181989
rect 226653 181961 226687 181989
rect 226715 181961 226749 181989
rect 226777 181961 226811 181989
rect 226839 181961 226887 181989
rect 226577 173175 226887 181961
rect 226577 173147 226625 173175
rect 226653 173147 226687 173175
rect 226715 173147 226749 173175
rect 226777 173147 226811 173175
rect 226839 173147 226887 173175
rect 226577 173113 226887 173147
rect 226577 173085 226625 173113
rect 226653 173085 226687 173113
rect 226715 173085 226749 173113
rect 226777 173085 226811 173113
rect 226839 173085 226887 173113
rect 226577 173051 226887 173085
rect 226577 173023 226625 173051
rect 226653 173023 226687 173051
rect 226715 173023 226749 173051
rect 226777 173023 226811 173051
rect 226839 173023 226887 173051
rect 226577 172989 226887 173023
rect 226577 172961 226625 172989
rect 226653 172961 226687 172989
rect 226715 172961 226749 172989
rect 226777 172961 226811 172989
rect 226839 172961 226887 172989
rect 226577 164175 226887 172961
rect 226577 164147 226625 164175
rect 226653 164147 226687 164175
rect 226715 164147 226749 164175
rect 226777 164147 226811 164175
rect 226839 164147 226887 164175
rect 226577 164113 226887 164147
rect 226577 164085 226625 164113
rect 226653 164085 226687 164113
rect 226715 164085 226749 164113
rect 226777 164085 226811 164113
rect 226839 164085 226887 164113
rect 226577 164051 226887 164085
rect 226577 164023 226625 164051
rect 226653 164023 226687 164051
rect 226715 164023 226749 164051
rect 226777 164023 226811 164051
rect 226839 164023 226887 164051
rect 226577 163989 226887 164023
rect 226577 163961 226625 163989
rect 226653 163961 226687 163989
rect 226715 163961 226749 163989
rect 226777 163961 226811 163989
rect 226839 163961 226887 163989
rect 226577 155175 226887 163961
rect 226577 155147 226625 155175
rect 226653 155147 226687 155175
rect 226715 155147 226749 155175
rect 226777 155147 226811 155175
rect 226839 155147 226887 155175
rect 226577 155113 226887 155147
rect 226577 155085 226625 155113
rect 226653 155085 226687 155113
rect 226715 155085 226749 155113
rect 226777 155085 226811 155113
rect 226839 155085 226887 155113
rect 226577 155051 226887 155085
rect 226577 155023 226625 155051
rect 226653 155023 226687 155051
rect 226715 155023 226749 155051
rect 226777 155023 226811 155051
rect 226839 155023 226887 155051
rect 226577 154989 226887 155023
rect 226577 154961 226625 154989
rect 226653 154961 226687 154989
rect 226715 154961 226749 154989
rect 226777 154961 226811 154989
rect 226839 154961 226887 154989
rect 226577 146175 226887 154961
rect 226577 146147 226625 146175
rect 226653 146147 226687 146175
rect 226715 146147 226749 146175
rect 226777 146147 226811 146175
rect 226839 146147 226887 146175
rect 226577 146113 226887 146147
rect 226577 146085 226625 146113
rect 226653 146085 226687 146113
rect 226715 146085 226749 146113
rect 226777 146085 226811 146113
rect 226839 146085 226887 146113
rect 226577 146051 226887 146085
rect 226577 146023 226625 146051
rect 226653 146023 226687 146051
rect 226715 146023 226749 146051
rect 226777 146023 226811 146051
rect 226839 146023 226887 146051
rect 226577 145989 226887 146023
rect 226577 145961 226625 145989
rect 226653 145961 226687 145989
rect 226715 145961 226749 145989
rect 226777 145961 226811 145989
rect 226839 145961 226887 145989
rect 226577 137175 226887 145961
rect 226577 137147 226625 137175
rect 226653 137147 226687 137175
rect 226715 137147 226749 137175
rect 226777 137147 226811 137175
rect 226839 137147 226887 137175
rect 226577 137113 226887 137147
rect 226577 137085 226625 137113
rect 226653 137085 226687 137113
rect 226715 137085 226749 137113
rect 226777 137085 226811 137113
rect 226839 137085 226887 137113
rect 226577 137051 226887 137085
rect 226577 137023 226625 137051
rect 226653 137023 226687 137051
rect 226715 137023 226749 137051
rect 226777 137023 226811 137051
rect 226839 137023 226887 137051
rect 226577 136989 226887 137023
rect 226577 136961 226625 136989
rect 226653 136961 226687 136989
rect 226715 136961 226749 136989
rect 226777 136961 226811 136989
rect 226839 136961 226887 136989
rect 226577 128175 226887 136961
rect 226577 128147 226625 128175
rect 226653 128147 226687 128175
rect 226715 128147 226749 128175
rect 226777 128147 226811 128175
rect 226839 128147 226887 128175
rect 226577 128113 226887 128147
rect 226577 128085 226625 128113
rect 226653 128085 226687 128113
rect 226715 128085 226749 128113
rect 226777 128085 226811 128113
rect 226839 128085 226887 128113
rect 226577 128051 226887 128085
rect 226577 128023 226625 128051
rect 226653 128023 226687 128051
rect 226715 128023 226749 128051
rect 226777 128023 226811 128051
rect 226839 128023 226887 128051
rect 226577 127989 226887 128023
rect 226577 127961 226625 127989
rect 226653 127961 226687 127989
rect 226715 127961 226749 127989
rect 226777 127961 226811 127989
rect 226839 127961 226887 127989
rect 226577 119175 226887 127961
rect 226577 119147 226625 119175
rect 226653 119147 226687 119175
rect 226715 119147 226749 119175
rect 226777 119147 226811 119175
rect 226839 119147 226887 119175
rect 226577 119113 226887 119147
rect 226577 119085 226625 119113
rect 226653 119085 226687 119113
rect 226715 119085 226749 119113
rect 226777 119085 226811 119113
rect 226839 119085 226887 119113
rect 226577 119051 226887 119085
rect 226577 119023 226625 119051
rect 226653 119023 226687 119051
rect 226715 119023 226749 119051
rect 226777 119023 226811 119051
rect 226839 119023 226887 119051
rect 226577 118989 226887 119023
rect 226577 118961 226625 118989
rect 226653 118961 226687 118989
rect 226715 118961 226749 118989
rect 226777 118961 226811 118989
rect 226839 118961 226887 118989
rect 226577 110175 226887 118961
rect 226577 110147 226625 110175
rect 226653 110147 226687 110175
rect 226715 110147 226749 110175
rect 226777 110147 226811 110175
rect 226839 110147 226887 110175
rect 226577 110113 226887 110147
rect 226577 110085 226625 110113
rect 226653 110085 226687 110113
rect 226715 110085 226749 110113
rect 226777 110085 226811 110113
rect 226839 110085 226887 110113
rect 226577 110051 226887 110085
rect 226577 110023 226625 110051
rect 226653 110023 226687 110051
rect 226715 110023 226749 110051
rect 226777 110023 226811 110051
rect 226839 110023 226887 110051
rect 226577 109989 226887 110023
rect 226577 109961 226625 109989
rect 226653 109961 226687 109989
rect 226715 109961 226749 109989
rect 226777 109961 226811 109989
rect 226839 109961 226887 109989
rect 226577 101175 226887 109961
rect 226577 101147 226625 101175
rect 226653 101147 226687 101175
rect 226715 101147 226749 101175
rect 226777 101147 226811 101175
rect 226839 101147 226887 101175
rect 226577 101113 226887 101147
rect 226577 101085 226625 101113
rect 226653 101085 226687 101113
rect 226715 101085 226749 101113
rect 226777 101085 226811 101113
rect 226839 101085 226887 101113
rect 226577 101051 226887 101085
rect 226577 101023 226625 101051
rect 226653 101023 226687 101051
rect 226715 101023 226749 101051
rect 226777 101023 226811 101051
rect 226839 101023 226887 101051
rect 226577 100989 226887 101023
rect 226577 100961 226625 100989
rect 226653 100961 226687 100989
rect 226715 100961 226749 100989
rect 226777 100961 226811 100989
rect 226839 100961 226887 100989
rect 226577 92175 226887 100961
rect 226577 92147 226625 92175
rect 226653 92147 226687 92175
rect 226715 92147 226749 92175
rect 226777 92147 226811 92175
rect 226839 92147 226887 92175
rect 226577 92113 226887 92147
rect 226577 92085 226625 92113
rect 226653 92085 226687 92113
rect 226715 92085 226749 92113
rect 226777 92085 226811 92113
rect 226839 92085 226887 92113
rect 226577 92051 226887 92085
rect 226577 92023 226625 92051
rect 226653 92023 226687 92051
rect 226715 92023 226749 92051
rect 226777 92023 226811 92051
rect 226839 92023 226887 92051
rect 226577 91989 226887 92023
rect 226577 91961 226625 91989
rect 226653 91961 226687 91989
rect 226715 91961 226749 91989
rect 226777 91961 226811 91989
rect 226839 91961 226887 91989
rect 226577 83175 226887 91961
rect 226577 83147 226625 83175
rect 226653 83147 226687 83175
rect 226715 83147 226749 83175
rect 226777 83147 226811 83175
rect 226839 83147 226887 83175
rect 226577 83113 226887 83147
rect 226577 83085 226625 83113
rect 226653 83085 226687 83113
rect 226715 83085 226749 83113
rect 226777 83085 226811 83113
rect 226839 83085 226887 83113
rect 226577 83051 226887 83085
rect 226577 83023 226625 83051
rect 226653 83023 226687 83051
rect 226715 83023 226749 83051
rect 226777 83023 226811 83051
rect 226839 83023 226887 83051
rect 226577 82989 226887 83023
rect 226577 82961 226625 82989
rect 226653 82961 226687 82989
rect 226715 82961 226749 82989
rect 226777 82961 226811 82989
rect 226839 82961 226887 82989
rect 226577 74175 226887 82961
rect 226577 74147 226625 74175
rect 226653 74147 226687 74175
rect 226715 74147 226749 74175
rect 226777 74147 226811 74175
rect 226839 74147 226887 74175
rect 226577 74113 226887 74147
rect 226577 74085 226625 74113
rect 226653 74085 226687 74113
rect 226715 74085 226749 74113
rect 226777 74085 226811 74113
rect 226839 74085 226887 74113
rect 226577 74051 226887 74085
rect 226577 74023 226625 74051
rect 226653 74023 226687 74051
rect 226715 74023 226749 74051
rect 226777 74023 226811 74051
rect 226839 74023 226887 74051
rect 226577 73989 226887 74023
rect 226577 73961 226625 73989
rect 226653 73961 226687 73989
rect 226715 73961 226749 73989
rect 226777 73961 226811 73989
rect 226839 73961 226887 73989
rect 226577 65175 226887 73961
rect 226577 65147 226625 65175
rect 226653 65147 226687 65175
rect 226715 65147 226749 65175
rect 226777 65147 226811 65175
rect 226839 65147 226887 65175
rect 226577 65113 226887 65147
rect 226577 65085 226625 65113
rect 226653 65085 226687 65113
rect 226715 65085 226749 65113
rect 226777 65085 226811 65113
rect 226839 65085 226887 65113
rect 226577 65051 226887 65085
rect 226577 65023 226625 65051
rect 226653 65023 226687 65051
rect 226715 65023 226749 65051
rect 226777 65023 226811 65051
rect 226839 65023 226887 65051
rect 226577 64989 226887 65023
rect 226577 64961 226625 64989
rect 226653 64961 226687 64989
rect 226715 64961 226749 64989
rect 226777 64961 226811 64989
rect 226839 64961 226887 64989
rect 226577 56175 226887 64961
rect 226577 56147 226625 56175
rect 226653 56147 226687 56175
rect 226715 56147 226749 56175
rect 226777 56147 226811 56175
rect 226839 56147 226887 56175
rect 226577 56113 226887 56147
rect 226577 56085 226625 56113
rect 226653 56085 226687 56113
rect 226715 56085 226749 56113
rect 226777 56085 226811 56113
rect 226839 56085 226887 56113
rect 226577 56051 226887 56085
rect 226577 56023 226625 56051
rect 226653 56023 226687 56051
rect 226715 56023 226749 56051
rect 226777 56023 226811 56051
rect 226839 56023 226887 56051
rect 226577 55989 226887 56023
rect 226577 55961 226625 55989
rect 226653 55961 226687 55989
rect 226715 55961 226749 55989
rect 226777 55961 226811 55989
rect 226839 55961 226887 55989
rect 226577 47175 226887 55961
rect 226577 47147 226625 47175
rect 226653 47147 226687 47175
rect 226715 47147 226749 47175
rect 226777 47147 226811 47175
rect 226839 47147 226887 47175
rect 226577 47113 226887 47147
rect 226577 47085 226625 47113
rect 226653 47085 226687 47113
rect 226715 47085 226749 47113
rect 226777 47085 226811 47113
rect 226839 47085 226887 47113
rect 226577 47051 226887 47085
rect 226577 47023 226625 47051
rect 226653 47023 226687 47051
rect 226715 47023 226749 47051
rect 226777 47023 226811 47051
rect 226839 47023 226887 47051
rect 226577 46989 226887 47023
rect 226577 46961 226625 46989
rect 226653 46961 226687 46989
rect 226715 46961 226749 46989
rect 226777 46961 226811 46989
rect 226839 46961 226887 46989
rect 226577 38175 226887 46961
rect 226577 38147 226625 38175
rect 226653 38147 226687 38175
rect 226715 38147 226749 38175
rect 226777 38147 226811 38175
rect 226839 38147 226887 38175
rect 226577 38113 226887 38147
rect 226577 38085 226625 38113
rect 226653 38085 226687 38113
rect 226715 38085 226749 38113
rect 226777 38085 226811 38113
rect 226839 38085 226887 38113
rect 226577 38051 226887 38085
rect 226577 38023 226625 38051
rect 226653 38023 226687 38051
rect 226715 38023 226749 38051
rect 226777 38023 226811 38051
rect 226839 38023 226887 38051
rect 226577 37989 226887 38023
rect 226577 37961 226625 37989
rect 226653 37961 226687 37989
rect 226715 37961 226749 37989
rect 226777 37961 226811 37989
rect 226839 37961 226887 37989
rect 226577 29175 226887 37961
rect 226577 29147 226625 29175
rect 226653 29147 226687 29175
rect 226715 29147 226749 29175
rect 226777 29147 226811 29175
rect 226839 29147 226887 29175
rect 226577 29113 226887 29147
rect 226577 29085 226625 29113
rect 226653 29085 226687 29113
rect 226715 29085 226749 29113
rect 226777 29085 226811 29113
rect 226839 29085 226887 29113
rect 226577 29051 226887 29085
rect 226577 29023 226625 29051
rect 226653 29023 226687 29051
rect 226715 29023 226749 29051
rect 226777 29023 226811 29051
rect 226839 29023 226887 29051
rect 226577 28989 226887 29023
rect 226577 28961 226625 28989
rect 226653 28961 226687 28989
rect 226715 28961 226749 28989
rect 226777 28961 226811 28989
rect 226839 28961 226887 28989
rect 226577 20175 226887 28961
rect 226577 20147 226625 20175
rect 226653 20147 226687 20175
rect 226715 20147 226749 20175
rect 226777 20147 226811 20175
rect 226839 20147 226887 20175
rect 226577 20113 226887 20147
rect 226577 20085 226625 20113
rect 226653 20085 226687 20113
rect 226715 20085 226749 20113
rect 226777 20085 226811 20113
rect 226839 20085 226887 20113
rect 226577 20051 226887 20085
rect 226577 20023 226625 20051
rect 226653 20023 226687 20051
rect 226715 20023 226749 20051
rect 226777 20023 226811 20051
rect 226839 20023 226887 20051
rect 226577 19989 226887 20023
rect 226577 19961 226625 19989
rect 226653 19961 226687 19989
rect 226715 19961 226749 19989
rect 226777 19961 226811 19989
rect 226839 19961 226887 19989
rect 226577 11175 226887 19961
rect 226577 11147 226625 11175
rect 226653 11147 226687 11175
rect 226715 11147 226749 11175
rect 226777 11147 226811 11175
rect 226839 11147 226887 11175
rect 226577 11113 226887 11147
rect 226577 11085 226625 11113
rect 226653 11085 226687 11113
rect 226715 11085 226749 11113
rect 226777 11085 226811 11113
rect 226839 11085 226887 11113
rect 226577 11051 226887 11085
rect 226577 11023 226625 11051
rect 226653 11023 226687 11051
rect 226715 11023 226749 11051
rect 226777 11023 226811 11051
rect 226839 11023 226887 11051
rect 226577 10989 226887 11023
rect 226577 10961 226625 10989
rect 226653 10961 226687 10989
rect 226715 10961 226749 10989
rect 226777 10961 226811 10989
rect 226839 10961 226887 10989
rect 226577 2175 226887 10961
rect 226577 2147 226625 2175
rect 226653 2147 226687 2175
rect 226715 2147 226749 2175
rect 226777 2147 226811 2175
rect 226839 2147 226887 2175
rect 226577 2113 226887 2147
rect 226577 2085 226625 2113
rect 226653 2085 226687 2113
rect 226715 2085 226749 2113
rect 226777 2085 226811 2113
rect 226839 2085 226887 2113
rect 226577 2051 226887 2085
rect 226577 2023 226625 2051
rect 226653 2023 226687 2051
rect 226715 2023 226749 2051
rect 226777 2023 226811 2051
rect 226839 2023 226887 2051
rect 226577 1989 226887 2023
rect 226577 1961 226625 1989
rect 226653 1961 226687 1989
rect 226715 1961 226749 1989
rect 226777 1961 226811 1989
rect 226839 1961 226887 1989
rect 226577 -80 226887 1961
rect 226577 -108 226625 -80
rect 226653 -108 226687 -80
rect 226715 -108 226749 -80
rect 226777 -108 226811 -80
rect 226839 -108 226887 -80
rect 226577 -142 226887 -108
rect 226577 -170 226625 -142
rect 226653 -170 226687 -142
rect 226715 -170 226749 -142
rect 226777 -170 226811 -142
rect 226839 -170 226887 -142
rect 226577 -204 226887 -170
rect 226577 -232 226625 -204
rect 226653 -232 226687 -204
rect 226715 -232 226749 -204
rect 226777 -232 226811 -204
rect 226839 -232 226887 -204
rect 226577 -266 226887 -232
rect 226577 -294 226625 -266
rect 226653 -294 226687 -266
rect 226715 -294 226749 -266
rect 226777 -294 226811 -266
rect 226839 -294 226887 -266
rect 226577 -822 226887 -294
rect 228437 299086 228747 299134
rect 228437 299058 228485 299086
rect 228513 299058 228547 299086
rect 228575 299058 228609 299086
rect 228637 299058 228671 299086
rect 228699 299058 228747 299086
rect 228437 299024 228747 299058
rect 228437 298996 228485 299024
rect 228513 298996 228547 299024
rect 228575 298996 228609 299024
rect 228637 298996 228671 299024
rect 228699 298996 228747 299024
rect 228437 298962 228747 298996
rect 228437 298934 228485 298962
rect 228513 298934 228547 298962
rect 228575 298934 228609 298962
rect 228637 298934 228671 298962
rect 228699 298934 228747 298962
rect 228437 298900 228747 298934
rect 228437 298872 228485 298900
rect 228513 298872 228547 298900
rect 228575 298872 228609 298900
rect 228637 298872 228671 298900
rect 228699 298872 228747 298900
rect 228437 293175 228747 298872
rect 228437 293147 228485 293175
rect 228513 293147 228547 293175
rect 228575 293147 228609 293175
rect 228637 293147 228671 293175
rect 228699 293147 228747 293175
rect 228437 293113 228747 293147
rect 228437 293085 228485 293113
rect 228513 293085 228547 293113
rect 228575 293085 228609 293113
rect 228637 293085 228671 293113
rect 228699 293085 228747 293113
rect 228437 293051 228747 293085
rect 228437 293023 228485 293051
rect 228513 293023 228547 293051
rect 228575 293023 228609 293051
rect 228637 293023 228671 293051
rect 228699 293023 228747 293051
rect 228437 292989 228747 293023
rect 228437 292961 228485 292989
rect 228513 292961 228547 292989
rect 228575 292961 228609 292989
rect 228637 292961 228671 292989
rect 228699 292961 228747 292989
rect 228437 284175 228747 292961
rect 228437 284147 228485 284175
rect 228513 284147 228547 284175
rect 228575 284147 228609 284175
rect 228637 284147 228671 284175
rect 228699 284147 228747 284175
rect 228437 284113 228747 284147
rect 228437 284085 228485 284113
rect 228513 284085 228547 284113
rect 228575 284085 228609 284113
rect 228637 284085 228671 284113
rect 228699 284085 228747 284113
rect 228437 284051 228747 284085
rect 228437 284023 228485 284051
rect 228513 284023 228547 284051
rect 228575 284023 228609 284051
rect 228637 284023 228671 284051
rect 228699 284023 228747 284051
rect 228437 283989 228747 284023
rect 228437 283961 228485 283989
rect 228513 283961 228547 283989
rect 228575 283961 228609 283989
rect 228637 283961 228671 283989
rect 228699 283961 228747 283989
rect 228437 275175 228747 283961
rect 228437 275147 228485 275175
rect 228513 275147 228547 275175
rect 228575 275147 228609 275175
rect 228637 275147 228671 275175
rect 228699 275147 228747 275175
rect 228437 275113 228747 275147
rect 228437 275085 228485 275113
rect 228513 275085 228547 275113
rect 228575 275085 228609 275113
rect 228637 275085 228671 275113
rect 228699 275085 228747 275113
rect 228437 275051 228747 275085
rect 228437 275023 228485 275051
rect 228513 275023 228547 275051
rect 228575 275023 228609 275051
rect 228637 275023 228671 275051
rect 228699 275023 228747 275051
rect 228437 274989 228747 275023
rect 228437 274961 228485 274989
rect 228513 274961 228547 274989
rect 228575 274961 228609 274989
rect 228637 274961 228671 274989
rect 228699 274961 228747 274989
rect 228437 266175 228747 274961
rect 228437 266147 228485 266175
rect 228513 266147 228547 266175
rect 228575 266147 228609 266175
rect 228637 266147 228671 266175
rect 228699 266147 228747 266175
rect 228437 266113 228747 266147
rect 228437 266085 228485 266113
rect 228513 266085 228547 266113
rect 228575 266085 228609 266113
rect 228637 266085 228671 266113
rect 228699 266085 228747 266113
rect 228437 266051 228747 266085
rect 228437 266023 228485 266051
rect 228513 266023 228547 266051
rect 228575 266023 228609 266051
rect 228637 266023 228671 266051
rect 228699 266023 228747 266051
rect 228437 265989 228747 266023
rect 228437 265961 228485 265989
rect 228513 265961 228547 265989
rect 228575 265961 228609 265989
rect 228637 265961 228671 265989
rect 228699 265961 228747 265989
rect 228437 257175 228747 265961
rect 228437 257147 228485 257175
rect 228513 257147 228547 257175
rect 228575 257147 228609 257175
rect 228637 257147 228671 257175
rect 228699 257147 228747 257175
rect 228437 257113 228747 257147
rect 228437 257085 228485 257113
rect 228513 257085 228547 257113
rect 228575 257085 228609 257113
rect 228637 257085 228671 257113
rect 228699 257085 228747 257113
rect 228437 257051 228747 257085
rect 228437 257023 228485 257051
rect 228513 257023 228547 257051
rect 228575 257023 228609 257051
rect 228637 257023 228671 257051
rect 228699 257023 228747 257051
rect 228437 256989 228747 257023
rect 228437 256961 228485 256989
rect 228513 256961 228547 256989
rect 228575 256961 228609 256989
rect 228637 256961 228671 256989
rect 228699 256961 228747 256989
rect 228437 248175 228747 256961
rect 228437 248147 228485 248175
rect 228513 248147 228547 248175
rect 228575 248147 228609 248175
rect 228637 248147 228671 248175
rect 228699 248147 228747 248175
rect 228437 248113 228747 248147
rect 228437 248085 228485 248113
rect 228513 248085 228547 248113
rect 228575 248085 228609 248113
rect 228637 248085 228671 248113
rect 228699 248085 228747 248113
rect 228437 248051 228747 248085
rect 228437 248023 228485 248051
rect 228513 248023 228547 248051
rect 228575 248023 228609 248051
rect 228637 248023 228671 248051
rect 228699 248023 228747 248051
rect 228437 247989 228747 248023
rect 228437 247961 228485 247989
rect 228513 247961 228547 247989
rect 228575 247961 228609 247989
rect 228637 247961 228671 247989
rect 228699 247961 228747 247989
rect 228437 239175 228747 247961
rect 228437 239147 228485 239175
rect 228513 239147 228547 239175
rect 228575 239147 228609 239175
rect 228637 239147 228671 239175
rect 228699 239147 228747 239175
rect 228437 239113 228747 239147
rect 228437 239085 228485 239113
rect 228513 239085 228547 239113
rect 228575 239085 228609 239113
rect 228637 239085 228671 239113
rect 228699 239085 228747 239113
rect 228437 239051 228747 239085
rect 228437 239023 228485 239051
rect 228513 239023 228547 239051
rect 228575 239023 228609 239051
rect 228637 239023 228671 239051
rect 228699 239023 228747 239051
rect 228437 238989 228747 239023
rect 228437 238961 228485 238989
rect 228513 238961 228547 238989
rect 228575 238961 228609 238989
rect 228637 238961 228671 238989
rect 228699 238961 228747 238989
rect 228437 230175 228747 238961
rect 228437 230147 228485 230175
rect 228513 230147 228547 230175
rect 228575 230147 228609 230175
rect 228637 230147 228671 230175
rect 228699 230147 228747 230175
rect 228437 230113 228747 230147
rect 228437 230085 228485 230113
rect 228513 230085 228547 230113
rect 228575 230085 228609 230113
rect 228637 230085 228671 230113
rect 228699 230085 228747 230113
rect 228437 230051 228747 230085
rect 228437 230023 228485 230051
rect 228513 230023 228547 230051
rect 228575 230023 228609 230051
rect 228637 230023 228671 230051
rect 228699 230023 228747 230051
rect 228437 229989 228747 230023
rect 228437 229961 228485 229989
rect 228513 229961 228547 229989
rect 228575 229961 228609 229989
rect 228637 229961 228671 229989
rect 228699 229961 228747 229989
rect 228437 221175 228747 229961
rect 228437 221147 228485 221175
rect 228513 221147 228547 221175
rect 228575 221147 228609 221175
rect 228637 221147 228671 221175
rect 228699 221147 228747 221175
rect 228437 221113 228747 221147
rect 228437 221085 228485 221113
rect 228513 221085 228547 221113
rect 228575 221085 228609 221113
rect 228637 221085 228671 221113
rect 228699 221085 228747 221113
rect 228437 221051 228747 221085
rect 228437 221023 228485 221051
rect 228513 221023 228547 221051
rect 228575 221023 228609 221051
rect 228637 221023 228671 221051
rect 228699 221023 228747 221051
rect 228437 220989 228747 221023
rect 228437 220961 228485 220989
rect 228513 220961 228547 220989
rect 228575 220961 228609 220989
rect 228637 220961 228671 220989
rect 228699 220961 228747 220989
rect 228437 212175 228747 220961
rect 228437 212147 228485 212175
rect 228513 212147 228547 212175
rect 228575 212147 228609 212175
rect 228637 212147 228671 212175
rect 228699 212147 228747 212175
rect 228437 212113 228747 212147
rect 228437 212085 228485 212113
rect 228513 212085 228547 212113
rect 228575 212085 228609 212113
rect 228637 212085 228671 212113
rect 228699 212085 228747 212113
rect 228437 212051 228747 212085
rect 228437 212023 228485 212051
rect 228513 212023 228547 212051
rect 228575 212023 228609 212051
rect 228637 212023 228671 212051
rect 228699 212023 228747 212051
rect 228437 211989 228747 212023
rect 228437 211961 228485 211989
rect 228513 211961 228547 211989
rect 228575 211961 228609 211989
rect 228637 211961 228671 211989
rect 228699 211961 228747 211989
rect 228437 203175 228747 211961
rect 228437 203147 228485 203175
rect 228513 203147 228547 203175
rect 228575 203147 228609 203175
rect 228637 203147 228671 203175
rect 228699 203147 228747 203175
rect 228437 203113 228747 203147
rect 228437 203085 228485 203113
rect 228513 203085 228547 203113
rect 228575 203085 228609 203113
rect 228637 203085 228671 203113
rect 228699 203085 228747 203113
rect 228437 203051 228747 203085
rect 228437 203023 228485 203051
rect 228513 203023 228547 203051
rect 228575 203023 228609 203051
rect 228637 203023 228671 203051
rect 228699 203023 228747 203051
rect 228437 202989 228747 203023
rect 228437 202961 228485 202989
rect 228513 202961 228547 202989
rect 228575 202961 228609 202989
rect 228637 202961 228671 202989
rect 228699 202961 228747 202989
rect 228437 194175 228747 202961
rect 228437 194147 228485 194175
rect 228513 194147 228547 194175
rect 228575 194147 228609 194175
rect 228637 194147 228671 194175
rect 228699 194147 228747 194175
rect 228437 194113 228747 194147
rect 228437 194085 228485 194113
rect 228513 194085 228547 194113
rect 228575 194085 228609 194113
rect 228637 194085 228671 194113
rect 228699 194085 228747 194113
rect 228437 194051 228747 194085
rect 228437 194023 228485 194051
rect 228513 194023 228547 194051
rect 228575 194023 228609 194051
rect 228637 194023 228671 194051
rect 228699 194023 228747 194051
rect 228437 193989 228747 194023
rect 228437 193961 228485 193989
rect 228513 193961 228547 193989
rect 228575 193961 228609 193989
rect 228637 193961 228671 193989
rect 228699 193961 228747 193989
rect 228437 185175 228747 193961
rect 228437 185147 228485 185175
rect 228513 185147 228547 185175
rect 228575 185147 228609 185175
rect 228637 185147 228671 185175
rect 228699 185147 228747 185175
rect 228437 185113 228747 185147
rect 228437 185085 228485 185113
rect 228513 185085 228547 185113
rect 228575 185085 228609 185113
rect 228637 185085 228671 185113
rect 228699 185085 228747 185113
rect 228437 185051 228747 185085
rect 228437 185023 228485 185051
rect 228513 185023 228547 185051
rect 228575 185023 228609 185051
rect 228637 185023 228671 185051
rect 228699 185023 228747 185051
rect 228437 184989 228747 185023
rect 228437 184961 228485 184989
rect 228513 184961 228547 184989
rect 228575 184961 228609 184989
rect 228637 184961 228671 184989
rect 228699 184961 228747 184989
rect 228437 176175 228747 184961
rect 228437 176147 228485 176175
rect 228513 176147 228547 176175
rect 228575 176147 228609 176175
rect 228637 176147 228671 176175
rect 228699 176147 228747 176175
rect 228437 176113 228747 176147
rect 228437 176085 228485 176113
rect 228513 176085 228547 176113
rect 228575 176085 228609 176113
rect 228637 176085 228671 176113
rect 228699 176085 228747 176113
rect 228437 176051 228747 176085
rect 228437 176023 228485 176051
rect 228513 176023 228547 176051
rect 228575 176023 228609 176051
rect 228637 176023 228671 176051
rect 228699 176023 228747 176051
rect 228437 175989 228747 176023
rect 228437 175961 228485 175989
rect 228513 175961 228547 175989
rect 228575 175961 228609 175989
rect 228637 175961 228671 175989
rect 228699 175961 228747 175989
rect 228437 167175 228747 175961
rect 228437 167147 228485 167175
rect 228513 167147 228547 167175
rect 228575 167147 228609 167175
rect 228637 167147 228671 167175
rect 228699 167147 228747 167175
rect 228437 167113 228747 167147
rect 228437 167085 228485 167113
rect 228513 167085 228547 167113
rect 228575 167085 228609 167113
rect 228637 167085 228671 167113
rect 228699 167085 228747 167113
rect 228437 167051 228747 167085
rect 228437 167023 228485 167051
rect 228513 167023 228547 167051
rect 228575 167023 228609 167051
rect 228637 167023 228671 167051
rect 228699 167023 228747 167051
rect 228437 166989 228747 167023
rect 228437 166961 228485 166989
rect 228513 166961 228547 166989
rect 228575 166961 228609 166989
rect 228637 166961 228671 166989
rect 228699 166961 228747 166989
rect 228437 158175 228747 166961
rect 228437 158147 228485 158175
rect 228513 158147 228547 158175
rect 228575 158147 228609 158175
rect 228637 158147 228671 158175
rect 228699 158147 228747 158175
rect 228437 158113 228747 158147
rect 228437 158085 228485 158113
rect 228513 158085 228547 158113
rect 228575 158085 228609 158113
rect 228637 158085 228671 158113
rect 228699 158085 228747 158113
rect 228437 158051 228747 158085
rect 228437 158023 228485 158051
rect 228513 158023 228547 158051
rect 228575 158023 228609 158051
rect 228637 158023 228671 158051
rect 228699 158023 228747 158051
rect 228437 157989 228747 158023
rect 228437 157961 228485 157989
rect 228513 157961 228547 157989
rect 228575 157961 228609 157989
rect 228637 157961 228671 157989
rect 228699 157961 228747 157989
rect 228437 149175 228747 157961
rect 228437 149147 228485 149175
rect 228513 149147 228547 149175
rect 228575 149147 228609 149175
rect 228637 149147 228671 149175
rect 228699 149147 228747 149175
rect 228437 149113 228747 149147
rect 228437 149085 228485 149113
rect 228513 149085 228547 149113
rect 228575 149085 228609 149113
rect 228637 149085 228671 149113
rect 228699 149085 228747 149113
rect 228437 149051 228747 149085
rect 228437 149023 228485 149051
rect 228513 149023 228547 149051
rect 228575 149023 228609 149051
rect 228637 149023 228671 149051
rect 228699 149023 228747 149051
rect 228437 148989 228747 149023
rect 228437 148961 228485 148989
rect 228513 148961 228547 148989
rect 228575 148961 228609 148989
rect 228637 148961 228671 148989
rect 228699 148961 228747 148989
rect 228437 140175 228747 148961
rect 228437 140147 228485 140175
rect 228513 140147 228547 140175
rect 228575 140147 228609 140175
rect 228637 140147 228671 140175
rect 228699 140147 228747 140175
rect 228437 140113 228747 140147
rect 228437 140085 228485 140113
rect 228513 140085 228547 140113
rect 228575 140085 228609 140113
rect 228637 140085 228671 140113
rect 228699 140085 228747 140113
rect 228437 140051 228747 140085
rect 228437 140023 228485 140051
rect 228513 140023 228547 140051
rect 228575 140023 228609 140051
rect 228637 140023 228671 140051
rect 228699 140023 228747 140051
rect 228437 139989 228747 140023
rect 228437 139961 228485 139989
rect 228513 139961 228547 139989
rect 228575 139961 228609 139989
rect 228637 139961 228671 139989
rect 228699 139961 228747 139989
rect 228437 131175 228747 139961
rect 228437 131147 228485 131175
rect 228513 131147 228547 131175
rect 228575 131147 228609 131175
rect 228637 131147 228671 131175
rect 228699 131147 228747 131175
rect 228437 131113 228747 131147
rect 228437 131085 228485 131113
rect 228513 131085 228547 131113
rect 228575 131085 228609 131113
rect 228637 131085 228671 131113
rect 228699 131085 228747 131113
rect 228437 131051 228747 131085
rect 228437 131023 228485 131051
rect 228513 131023 228547 131051
rect 228575 131023 228609 131051
rect 228637 131023 228671 131051
rect 228699 131023 228747 131051
rect 228437 130989 228747 131023
rect 228437 130961 228485 130989
rect 228513 130961 228547 130989
rect 228575 130961 228609 130989
rect 228637 130961 228671 130989
rect 228699 130961 228747 130989
rect 228437 122175 228747 130961
rect 228437 122147 228485 122175
rect 228513 122147 228547 122175
rect 228575 122147 228609 122175
rect 228637 122147 228671 122175
rect 228699 122147 228747 122175
rect 228437 122113 228747 122147
rect 228437 122085 228485 122113
rect 228513 122085 228547 122113
rect 228575 122085 228609 122113
rect 228637 122085 228671 122113
rect 228699 122085 228747 122113
rect 228437 122051 228747 122085
rect 228437 122023 228485 122051
rect 228513 122023 228547 122051
rect 228575 122023 228609 122051
rect 228637 122023 228671 122051
rect 228699 122023 228747 122051
rect 228437 121989 228747 122023
rect 228437 121961 228485 121989
rect 228513 121961 228547 121989
rect 228575 121961 228609 121989
rect 228637 121961 228671 121989
rect 228699 121961 228747 121989
rect 228437 113175 228747 121961
rect 228437 113147 228485 113175
rect 228513 113147 228547 113175
rect 228575 113147 228609 113175
rect 228637 113147 228671 113175
rect 228699 113147 228747 113175
rect 228437 113113 228747 113147
rect 228437 113085 228485 113113
rect 228513 113085 228547 113113
rect 228575 113085 228609 113113
rect 228637 113085 228671 113113
rect 228699 113085 228747 113113
rect 228437 113051 228747 113085
rect 228437 113023 228485 113051
rect 228513 113023 228547 113051
rect 228575 113023 228609 113051
rect 228637 113023 228671 113051
rect 228699 113023 228747 113051
rect 228437 112989 228747 113023
rect 228437 112961 228485 112989
rect 228513 112961 228547 112989
rect 228575 112961 228609 112989
rect 228637 112961 228671 112989
rect 228699 112961 228747 112989
rect 228437 104175 228747 112961
rect 228437 104147 228485 104175
rect 228513 104147 228547 104175
rect 228575 104147 228609 104175
rect 228637 104147 228671 104175
rect 228699 104147 228747 104175
rect 228437 104113 228747 104147
rect 228437 104085 228485 104113
rect 228513 104085 228547 104113
rect 228575 104085 228609 104113
rect 228637 104085 228671 104113
rect 228699 104085 228747 104113
rect 228437 104051 228747 104085
rect 228437 104023 228485 104051
rect 228513 104023 228547 104051
rect 228575 104023 228609 104051
rect 228637 104023 228671 104051
rect 228699 104023 228747 104051
rect 228437 103989 228747 104023
rect 228437 103961 228485 103989
rect 228513 103961 228547 103989
rect 228575 103961 228609 103989
rect 228637 103961 228671 103989
rect 228699 103961 228747 103989
rect 228437 95175 228747 103961
rect 228437 95147 228485 95175
rect 228513 95147 228547 95175
rect 228575 95147 228609 95175
rect 228637 95147 228671 95175
rect 228699 95147 228747 95175
rect 228437 95113 228747 95147
rect 228437 95085 228485 95113
rect 228513 95085 228547 95113
rect 228575 95085 228609 95113
rect 228637 95085 228671 95113
rect 228699 95085 228747 95113
rect 228437 95051 228747 95085
rect 228437 95023 228485 95051
rect 228513 95023 228547 95051
rect 228575 95023 228609 95051
rect 228637 95023 228671 95051
rect 228699 95023 228747 95051
rect 228437 94989 228747 95023
rect 228437 94961 228485 94989
rect 228513 94961 228547 94989
rect 228575 94961 228609 94989
rect 228637 94961 228671 94989
rect 228699 94961 228747 94989
rect 228437 86175 228747 94961
rect 228437 86147 228485 86175
rect 228513 86147 228547 86175
rect 228575 86147 228609 86175
rect 228637 86147 228671 86175
rect 228699 86147 228747 86175
rect 228437 86113 228747 86147
rect 228437 86085 228485 86113
rect 228513 86085 228547 86113
rect 228575 86085 228609 86113
rect 228637 86085 228671 86113
rect 228699 86085 228747 86113
rect 228437 86051 228747 86085
rect 228437 86023 228485 86051
rect 228513 86023 228547 86051
rect 228575 86023 228609 86051
rect 228637 86023 228671 86051
rect 228699 86023 228747 86051
rect 228437 85989 228747 86023
rect 228437 85961 228485 85989
rect 228513 85961 228547 85989
rect 228575 85961 228609 85989
rect 228637 85961 228671 85989
rect 228699 85961 228747 85989
rect 228437 77175 228747 85961
rect 228437 77147 228485 77175
rect 228513 77147 228547 77175
rect 228575 77147 228609 77175
rect 228637 77147 228671 77175
rect 228699 77147 228747 77175
rect 228437 77113 228747 77147
rect 228437 77085 228485 77113
rect 228513 77085 228547 77113
rect 228575 77085 228609 77113
rect 228637 77085 228671 77113
rect 228699 77085 228747 77113
rect 228437 77051 228747 77085
rect 228437 77023 228485 77051
rect 228513 77023 228547 77051
rect 228575 77023 228609 77051
rect 228637 77023 228671 77051
rect 228699 77023 228747 77051
rect 228437 76989 228747 77023
rect 228437 76961 228485 76989
rect 228513 76961 228547 76989
rect 228575 76961 228609 76989
rect 228637 76961 228671 76989
rect 228699 76961 228747 76989
rect 228437 68175 228747 76961
rect 228437 68147 228485 68175
rect 228513 68147 228547 68175
rect 228575 68147 228609 68175
rect 228637 68147 228671 68175
rect 228699 68147 228747 68175
rect 228437 68113 228747 68147
rect 228437 68085 228485 68113
rect 228513 68085 228547 68113
rect 228575 68085 228609 68113
rect 228637 68085 228671 68113
rect 228699 68085 228747 68113
rect 228437 68051 228747 68085
rect 228437 68023 228485 68051
rect 228513 68023 228547 68051
rect 228575 68023 228609 68051
rect 228637 68023 228671 68051
rect 228699 68023 228747 68051
rect 228437 67989 228747 68023
rect 228437 67961 228485 67989
rect 228513 67961 228547 67989
rect 228575 67961 228609 67989
rect 228637 67961 228671 67989
rect 228699 67961 228747 67989
rect 228437 59175 228747 67961
rect 228437 59147 228485 59175
rect 228513 59147 228547 59175
rect 228575 59147 228609 59175
rect 228637 59147 228671 59175
rect 228699 59147 228747 59175
rect 228437 59113 228747 59147
rect 228437 59085 228485 59113
rect 228513 59085 228547 59113
rect 228575 59085 228609 59113
rect 228637 59085 228671 59113
rect 228699 59085 228747 59113
rect 228437 59051 228747 59085
rect 228437 59023 228485 59051
rect 228513 59023 228547 59051
rect 228575 59023 228609 59051
rect 228637 59023 228671 59051
rect 228699 59023 228747 59051
rect 228437 58989 228747 59023
rect 228437 58961 228485 58989
rect 228513 58961 228547 58989
rect 228575 58961 228609 58989
rect 228637 58961 228671 58989
rect 228699 58961 228747 58989
rect 228437 50175 228747 58961
rect 228437 50147 228485 50175
rect 228513 50147 228547 50175
rect 228575 50147 228609 50175
rect 228637 50147 228671 50175
rect 228699 50147 228747 50175
rect 228437 50113 228747 50147
rect 228437 50085 228485 50113
rect 228513 50085 228547 50113
rect 228575 50085 228609 50113
rect 228637 50085 228671 50113
rect 228699 50085 228747 50113
rect 228437 50051 228747 50085
rect 228437 50023 228485 50051
rect 228513 50023 228547 50051
rect 228575 50023 228609 50051
rect 228637 50023 228671 50051
rect 228699 50023 228747 50051
rect 228437 49989 228747 50023
rect 228437 49961 228485 49989
rect 228513 49961 228547 49989
rect 228575 49961 228609 49989
rect 228637 49961 228671 49989
rect 228699 49961 228747 49989
rect 228437 41175 228747 49961
rect 228437 41147 228485 41175
rect 228513 41147 228547 41175
rect 228575 41147 228609 41175
rect 228637 41147 228671 41175
rect 228699 41147 228747 41175
rect 228437 41113 228747 41147
rect 228437 41085 228485 41113
rect 228513 41085 228547 41113
rect 228575 41085 228609 41113
rect 228637 41085 228671 41113
rect 228699 41085 228747 41113
rect 228437 41051 228747 41085
rect 228437 41023 228485 41051
rect 228513 41023 228547 41051
rect 228575 41023 228609 41051
rect 228637 41023 228671 41051
rect 228699 41023 228747 41051
rect 228437 40989 228747 41023
rect 228437 40961 228485 40989
rect 228513 40961 228547 40989
rect 228575 40961 228609 40989
rect 228637 40961 228671 40989
rect 228699 40961 228747 40989
rect 228437 32175 228747 40961
rect 228437 32147 228485 32175
rect 228513 32147 228547 32175
rect 228575 32147 228609 32175
rect 228637 32147 228671 32175
rect 228699 32147 228747 32175
rect 228437 32113 228747 32147
rect 228437 32085 228485 32113
rect 228513 32085 228547 32113
rect 228575 32085 228609 32113
rect 228637 32085 228671 32113
rect 228699 32085 228747 32113
rect 228437 32051 228747 32085
rect 228437 32023 228485 32051
rect 228513 32023 228547 32051
rect 228575 32023 228609 32051
rect 228637 32023 228671 32051
rect 228699 32023 228747 32051
rect 228437 31989 228747 32023
rect 228437 31961 228485 31989
rect 228513 31961 228547 31989
rect 228575 31961 228609 31989
rect 228637 31961 228671 31989
rect 228699 31961 228747 31989
rect 228437 23175 228747 31961
rect 228437 23147 228485 23175
rect 228513 23147 228547 23175
rect 228575 23147 228609 23175
rect 228637 23147 228671 23175
rect 228699 23147 228747 23175
rect 228437 23113 228747 23147
rect 228437 23085 228485 23113
rect 228513 23085 228547 23113
rect 228575 23085 228609 23113
rect 228637 23085 228671 23113
rect 228699 23085 228747 23113
rect 228437 23051 228747 23085
rect 228437 23023 228485 23051
rect 228513 23023 228547 23051
rect 228575 23023 228609 23051
rect 228637 23023 228671 23051
rect 228699 23023 228747 23051
rect 228437 22989 228747 23023
rect 228437 22961 228485 22989
rect 228513 22961 228547 22989
rect 228575 22961 228609 22989
rect 228637 22961 228671 22989
rect 228699 22961 228747 22989
rect 228437 14175 228747 22961
rect 228437 14147 228485 14175
rect 228513 14147 228547 14175
rect 228575 14147 228609 14175
rect 228637 14147 228671 14175
rect 228699 14147 228747 14175
rect 228437 14113 228747 14147
rect 228437 14085 228485 14113
rect 228513 14085 228547 14113
rect 228575 14085 228609 14113
rect 228637 14085 228671 14113
rect 228699 14085 228747 14113
rect 228437 14051 228747 14085
rect 228437 14023 228485 14051
rect 228513 14023 228547 14051
rect 228575 14023 228609 14051
rect 228637 14023 228671 14051
rect 228699 14023 228747 14051
rect 228437 13989 228747 14023
rect 228437 13961 228485 13989
rect 228513 13961 228547 13989
rect 228575 13961 228609 13989
rect 228637 13961 228671 13989
rect 228699 13961 228747 13989
rect 228437 5175 228747 13961
rect 228437 5147 228485 5175
rect 228513 5147 228547 5175
rect 228575 5147 228609 5175
rect 228637 5147 228671 5175
rect 228699 5147 228747 5175
rect 228437 5113 228747 5147
rect 228437 5085 228485 5113
rect 228513 5085 228547 5113
rect 228575 5085 228609 5113
rect 228637 5085 228671 5113
rect 228699 5085 228747 5113
rect 228437 5051 228747 5085
rect 228437 5023 228485 5051
rect 228513 5023 228547 5051
rect 228575 5023 228609 5051
rect 228637 5023 228671 5051
rect 228699 5023 228747 5051
rect 228437 4989 228747 5023
rect 228437 4961 228485 4989
rect 228513 4961 228547 4989
rect 228575 4961 228609 4989
rect 228637 4961 228671 4989
rect 228699 4961 228747 4989
rect 228437 -560 228747 4961
rect 228437 -588 228485 -560
rect 228513 -588 228547 -560
rect 228575 -588 228609 -560
rect 228637 -588 228671 -560
rect 228699 -588 228747 -560
rect 228437 -622 228747 -588
rect 228437 -650 228485 -622
rect 228513 -650 228547 -622
rect 228575 -650 228609 -622
rect 228637 -650 228671 -622
rect 228699 -650 228747 -622
rect 228437 -684 228747 -650
rect 228437 -712 228485 -684
rect 228513 -712 228547 -684
rect 228575 -712 228609 -684
rect 228637 -712 228671 -684
rect 228699 -712 228747 -684
rect 228437 -746 228747 -712
rect 228437 -774 228485 -746
rect 228513 -774 228547 -746
rect 228575 -774 228609 -746
rect 228637 -774 228671 -746
rect 228699 -774 228747 -746
rect 228437 -822 228747 -774
rect 235577 298606 235887 299134
rect 235577 298578 235625 298606
rect 235653 298578 235687 298606
rect 235715 298578 235749 298606
rect 235777 298578 235811 298606
rect 235839 298578 235887 298606
rect 235577 298544 235887 298578
rect 235577 298516 235625 298544
rect 235653 298516 235687 298544
rect 235715 298516 235749 298544
rect 235777 298516 235811 298544
rect 235839 298516 235887 298544
rect 235577 298482 235887 298516
rect 235577 298454 235625 298482
rect 235653 298454 235687 298482
rect 235715 298454 235749 298482
rect 235777 298454 235811 298482
rect 235839 298454 235887 298482
rect 235577 298420 235887 298454
rect 235577 298392 235625 298420
rect 235653 298392 235687 298420
rect 235715 298392 235749 298420
rect 235777 298392 235811 298420
rect 235839 298392 235887 298420
rect 235577 290175 235887 298392
rect 235577 290147 235625 290175
rect 235653 290147 235687 290175
rect 235715 290147 235749 290175
rect 235777 290147 235811 290175
rect 235839 290147 235887 290175
rect 235577 290113 235887 290147
rect 235577 290085 235625 290113
rect 235653 290085 235687 290113
rect 235715 290085 235749 290113
rect 235777 290085 235811 290113
rect 235839 290085 235887 290113
rect 235577 290051 235887 290085
rect 235577 290023 235625 290051
rect 235653 290023 235687 290051
rect 235715 290023 235749 290051
rect 235777 290023 235811 290051
rect 235839 290023 235887 290051
rect 235577 289989 235887 290023
rect 235577 289961 235625 289989
rect 235653 289961 235687 289989
rect 235715 289961 235749 289989
rect 235777 289961 235811 289989
rect 235839 289961 235887 289989
rect 235577 281175 235887 289961
rect 235577 281147 235625 281175
rect 235653 281147 235687 281175
rect 235715 281147 235749 281175
rect 235777 281147 235811 281175
rect 235839 281147 235887 281175
rect 235577 281113 235887 281147
rect 235577 281085 235625 281113
rect 235653 281085 235687 281113
rect 235715 281085 235749 281113
rect 235777 281085 235811 281113
rect 235839 281085 235887 281113
rect 235577 281051 235887 281085
rect 235577 281023 235625 281051
rect 235653 281023 235687 281051
rect 235715 281023 235749 281051
rect 235777 281023 235811 281051
rect 235839 281023 235887 281051
rect 235577 280989 235887 281023
rect 235577 280961 235625 280989
rect 235653 280961 235687 280989
rect 235715 280961 235749 280989
rect 235777 280961 235811 280989
rect 235839 280961 235887 280989
rect 235577 272175 235887 280961
rect 235577 272147 235625 272175
rect 235653 272147 235687 272175
rect 235715 272147 235749 272175
rect 235777 272147 235811 272175
rect 235839 272147 235887 272175
rect 235577 272113 235887 272147
rect 235577 272085 235625 272113
rect 235653 272085 235687 272113
rect 235715 272085 235749 272113
rect 235777 272085 235811 272113
rect 235839 272085 235887 272113
rect 235577 272051 235887 272085
rect 235577 272023 235625 272051
rect 235653 272023 235687 272051
rect 235715 272023 235749 272051
rect 235777 272023 235811 272051
rect 235839 272023 235887 272051
rect 235577 271989 235887 272023
rect 235577 271961 235625 271989
rect 235653 271961 235687 271989
rect 235715 271961 235749 271989
rect 235777 271961 235811 271989
rect 235839 271961 235887 271989
rect 235577 263175 235887 271961
rect 235577 263147 235625 263175
rect 235653 263147 235687 263175
rect 235715 263147 235749 263175
rect 235777 263147 235811 263175
rect 235839 263147 235887 263175
rect 235577 263113 235887 263147
rect 235577 263085 235625 263113
rect 235653 263085 235687 263113
rect 235715 263085 235749 263113
rect 235777 263085 235811 263113
rect 235839 263085 235887 263113
rect 235577 263051 235887 263085
rect 235577 263023 235625 263051
rect 235653 263023 235687 263051
rect 235715 263023 235749 263051
rect 235777 263023 235811 263051
rect 235839 263023 235887 263051
rect 235577 262989 235887 263023
rect 235577 262961 235625 262989
rect 235653 262961 235687 262989
rect 235715 262961 235749 262989
rect 235777 262961 235811 262989
rect 235839 262961 235887 262989
rect 235577 254175 235887 262961
rect 235577 254147 235625 254175
rect 235653 254147 235687 254175
rect 235715 254147 235749 254175
rect 235777 254147 235811 254175
rect 235839 254147 235887 254175
rect 235577 254113 235887 254147
rect 235577 254085 235625 254113
rect 235653 254085 235687 254113
rect 235715 254085 235749 254113
rect 235777 254085 235811 254113
rect 235839 254085 235887 254113
rect 235577 254051 235887 254085
rect 235577 254023 235625 254051
rect 235653 254023 235687 254051
rect 235715 254023 235749 254051
rect 235777 254023 235811 254051
rect 235839 254023 235887 254051
rect 235577 253989 235887 254023
rect 235577 253961 235625 253989
rect 235653 253961 235687 253989
rect 235715 253961 235749 253989
rect 235777 253961 235811 253989
rect 235839 253961 235887 253989
rect 235577 245175 235887 253961
rect 235577 245147 235625 245175
rect 235653 245147 235687 245175
rect 235715 245147 235749 245175
rect 235777 245147 235811 245175
rect 235839 245147 235887 245175
rect 235577 245113 235887 245147
rect 235577 245085 235625 245113
rect 235653 245085 235687 245113
rect 235715 245085 235749 245113
rect 235777 245085 235811 245113
rect 235839 245085 235887 245113
rect 235577 245051 235887 245085
rect 235577 245023 235625 245051
rect 235653 245023 235687 245051
rect 235715 245023 235749 245051
rect 235777 245023 235811 245051
rect 235839 245023 235887 245051
rect 235577 244989 235887 245023
rect 235577 244961 235625 244989
rect 235653 244961 235687 244989
rect 235715 244961 235749 244989
rect 235777 244961 235811 244989
rect 235839 244961 235887 244989
rect 235577 236175 235887 244961
rect 235577 236147 235625 236175
rect 235653 236147 235687 236175
rect 235715 236147 235749 236175
rect 235777 236147 235811 236175
rect 235839 236147 235887 236175
rect 235577 236113 235887 236147
rect 235577 236085 235625 236113
rect 235653 236085 235687 236113
rect 235715 236085 235749 236113
rect 235777 236085 235811 236113
rect 235839 236085 235887 236113
rect 235577 236051 235887 236085
rect 235577 236023 235625 236051
rect 235653 236023 235687 236051
rect 235715 236023 235749 236051
rect 235777 236023 235811 236051
rect 235839 236023 235887 236051
rect 235577 235989 235887 236023
rect 235577 235961 235625 235989
rect 235653 235961 235687 235989
rect 235715 235961 235749 235989
rect 235777 235961 235811 235989
rect 235839 235961 235887 235989
rect 235577 227175 235887 235961
rect 235577 227147 235625 227175
rect 235653 227147 235687 227175
rect 235715 227147 235749 227175
rect 235777 227147 235811 227175
rect 235839 227147 235887 227175
rect 235577 227113 235887 227147
rect 235577 227085 235625 227113
rect 235653 227085 235687 227113
rect 235715 227085 235749 227113
rect 235777 227085 235811 227113
rect 235839 227085 235887 227113
rect 235577 227051 235887 227085
rect 235577 227023 235625 227051
rect 235653 227023 235687 227051
rect 235715 227023 235749 227051
rect 235777 227023 235811 227051
rect 235839 227023 235887 227051
rect 235577 226989 235887 227023
rect 235577 226961 235625 226989
rect 235653 226961 235687 226989
rect 235715 226961 235749 226989
rect 235777 226961 235811 226989
rect 235839 226961 235887 226989
rect 235577 218175 235887 226961
rect 235577 218147 235625 218175
rect 235653 218147 235687 218175
rect 235715 218147 235749 218175
rect 235777 218147 235811 218175
rect 235839 218147 235887 218175
rect 235577 218113 235887 218147
rect 235577 218085 235625 218113
rect 235653 218085 235687 218113
rect 235715 218085 235749 218113
rect 235777 218085 235811 218113
rect 235839 218085 235887 218113
rect 235577 218051 235887 218085
rect 235577 218023 235625 218051
rect 235653 218023 235687 218051
rect 235715 218023 235749 218051
rect 235777 218023 235811 218051
rect 235839 218023 235887 218051
rect 235577 217989 235887 218023
rect 235577 217961 235625 217989
rect 235653 217961 235687 217989
rect 235715 217961 235749 217989
rect 235777 217961 235811 217989
rect 235839 217961 235887 217989
rect 235577 209175 235887 217961
rect 235577 209147 235625 209175
rect 235653 209147 235687 209175
rect 235715 209147 235749 209175
rect 235777 209147 235811 209175
rect 235839 209147 235887 209175
rect 235577 209113 235887 209147
rect 235577 209085 235625 209113
rect 235653 209085 235687 209113
rect 235715 209085 235749 209113
rect 235777 209085 235811 209113
rect 235839 209085 235887 209113
rect 235577 209051 235887 209085
rect 235577 209023 235625 209051
rect 235653 209023 235687 209051
rect 235715 209023 235749 209051
rect 235777 209023 235811 209051
rect 235839 209023 235887 209051
rect 235577 208989 235887 209023
rect 235577 208961 235625 208989
rect 235653 208961 235687 208989
rect 235715 208961 235749 208989
rect 235777 208961 235811 208989
rect 235839 208961 235887 208989
rect 235577 200175 235887 208961
rect 235577 200147 235625 200175
rect 235653 200147 235687 200175
rect 235715 200147 235749 200175
rect 235777 200147 235811 200175
rect 235839 200147 235887 200175
rect 235577 200113 235887 200147
rect 235577 200085 235625 200113
rect 235653 200085 235687 200113
rect 235715 200085 235749 200113
rect 235777 200085 235811 200113
rect 235839 200085 235887 200113
rect 235577 200051 235887 200085
rect 235577 200023 235625 200051
rect 235653 200023 235687 200051
rect 235715 200023 235749 200051
rect 235777 200023 235811 200051
rect 235839 200023 235887 200051
rect 235577 199989 235887 200023
rect 235577 199961 235625 199989
rect 235653 199961 235687 199989
rect 235715 199961 235749 199989
rect 235777 199961 235811 199989
rect 235839 199961 235887 199989
rect 235577 191175 235887 199961
rect 235577 191147 235625 191175
rect 235653 191147 235687 191175
rect 235715 191147 235749 191175
rect 235777 191147 235811 191175
rect 235839 191147 235887 191175
rect 235577 191113 235887 191147
rect 235577 191085 235625 191113
rect 235653 191085 235687 191113
rect 235715 191085 235749 191113
rect 235777 191085 235811 191113
rect 235839 191085 235887 191113
rect 235577 191051 235887 191085
rect 235577 191023 235625 191051
rect 235653 191023 235687 191051
rect 235715 191023 235749 191051
rect 235777 191023 235811 191051
rect 235839 191023 235887 191051
rect 235577 190989 235887 191023
rect 235577 190961 235625 190989
rect 235653 190961 235687 190989
rect 235715 190961 235749 190989
rect 235777 190961 235811 190989
rect 235839 190961 235887 190989
rect 235577 182175 235887 190961
rect 235577 182147 235625 182175
rect 235653 182147 235687 182175
rect 235715 182147 235749 182175
rect 235777 182147 235811 182175
rect 235839 182147 235887 182175
rect 235577 182113 235887 182147
rect 235577 182085 235625 182113
rect 235653 182085 235687 182113
rect 235715 182085 235749 182113
rect 235777 182085 235811 182113
rect 235839 182085 235887 182113
rect 235577 182051 235887 182085
rect 235577 182023 235625 182051
rect 235653 182023 235687 182051
rect 235715 182023 235749 182051
rect 235777 182023 235811 182051
rect 235839 182023 235887 182051
rect 235577 181989 235887 182023
rect 235577 181961 235625 181989
rect 235653 181961 235687 181989
rect 235715 181961 235749 181989
rect 235777 181961 235811 181989
rect 235839 181961 235887 181989
rect 235577 173175 235887 181961
rect 235577 173147 235625 173175
rect 235653 173147 235687 173175
rect 235715 173147 235749 173175
rect 235777 173147 235811 173175
rect 235839 173147 235887 173175
rect 235577 173113 235887 173147
rect 235577 173085 235625 173113
rect 235653 173085 235687 173113
rect 235715 173085 235749 173113
rect 235777 173085 235811 173113
rect 235839 173085 235887 173113
rect 235577 173051 235887 173085
rect 235577 173023 235625 173051
rect 235653 173023 235687 173051
rect 235715 173023 235749 173051
rect 235777 173023 235811 173051
rect 235839 173023 235887 173051
rect 235577 172989 235887 173023
rect 235577 172961 235625 172989
rect 235653 172961 235687 172989
rect 235715 172961 235749 172989
rect 235777 172961 235811 172989
rect 235839 172961 235887 172989
rect 235577 164175 235887 172961
rect 235577 164147 235625 164175
rect 235653 164147 235687 164175
rect 235715 164147 235749 164175
rect 235777 164147 235811 164175
rect 235839 164147 235887 164175
rect 235577 164113 235887 164147
rect 235577 164085 235625 164113
rect 235653 164085 235687 164113
rect 235715 164085 235749 164113
rect 235777 164085 235811 164113
rect 235839 164085 235887 164113
rect 235577 164051 235887 164085
rect 235577 164023 235625 164051
rect 235653 164023 235687 164051
rect 235715 164023 235749 164051
rect 235777 164023 235811 164051
rect 235839 164023 235887 164051
rect 235577 163989 235887 164023
rect 235577 163961 235625 163989
rect 235653 163961 235687 163989
rect 235715 163961 235749 163989
rect 235777 163961 235811 163989
rect 235839 163961 235887 163989
rect 235577 155175 235887 163961
rect 235577 155147 235625 155175
rect 235653 155147 235687 155175
rect 235715 155147 235749 155175
rect 235777 155147 235811 155175
rect 235839 155147 235887 155175
rect 235577 155113 235887 155147
rect 235577 155085 235625 155113
rect 235653 155085 235687 155113
rect 235715 155085 235749 155113
rect 235777 155085 235811 155113
rect 235839 155085 235887 155113
rect 235577 155051 235887 155085
rect 235577 155023 235625 155051
rect 235653 155023 235687 155051
rect 235715 155023 235749 155051
rect 235777 155023 235811 155051
rect 235839 155023 235887 155051
rect 235577 154989 235887 155023
rect 235577 154961 235625 154989
rect 235653 154961 235687 154989
rect 235715 154961 235749 154989
rect 235777 154961 235811 154989
rect 235839 154961 235887 154989
rect 235577 146175 235887 154961
rect 235577 146147 235625 146175
rect 235653 146147 235687 146175
rect 235715 146147 235749 146175
rect 235777 146147 235811 146175
rect 235839 146147 235887 146175
rect 235577 146113 235887 146147
rect 235577 146085 235625 146113
rect 235653 146085 235687 146113
rect 235715 146085 235749 146113
rect 235777 146085 235811 146113
rect 235839 146085 235887 146113
rect 235577 146051 235887 146085
rect 235577 146023 235625 146051
rect 235653 146023 235687 146051
rect 235715 146023 235749 146051
rect 235777 146023 235811 146051
rect 235839 146023 235887 146051
rect 235577 145989 235887 146023
rect 235577 145961 235625 145989
rect 235653 145961 235687 145989
rect 235715 145961 235749 145989
rect 235777 145961 235811 145989
rect 235839 145961 235887 145989
rect 235577 137175 235887 145961
rect 235577 137147 235625 137175
rect 235653 137147 235687 137175
rect 235715 137147 235749 137175
rect 235777 137147 235811 137175
rect 235839 137147 235887 137175
rect 235577 137113 235887 137147
rect 235577 137085 235625 137113
rect 235653 137085 235687 137113
rect 235715 137085 235749 137113
rect 235777 137085 235811 137113
rect 235839 137085 235887 137113
rect 235577 137051 235887 137085
rect 235577 137023 235625 137051
rect 235653 137023 235687 137051
rect 235715 137023 235749 137051
rect 235777 137023 235811 137051
rect 235839 137023 235887 137051
rect 235577 136989 235887 137023
rect 235577 136961 235625 136989
rect 235653 136961 235687 136989
rect 235715 136961 235749 136989
rect 235777 136961 235811 136989
rect 235839 136961 235887 136989
rect 235577 128175 235887 136961
rect 235577 128147 235625 128175
rect 235653 128147 235687 128175
rect 235715 128147 235749 128175
rect 235777 128147 235811 128175
rect 235839 128147 235887 128175
rect 235577 128113 235887 128147
rect 235577 128085 235625 128113
rect 235653 128085 235687 128113
rect 235715 128085 235749 128113
rect 235777 128085 235811 128113
rect 235839 128085 235887 128113
rect 235577 128051 235887 128085
rect 235577 128023 235625 128051
rect 235653 128023 235687 128051
rect 235715 128023 235749 128051
rect 235777 128023 235811 128051
rect 235839 128023 235887 128051
rect 235577 127989 235887 128023
rect 235577 127961 235625 127989
rect 235653 127961 235687 127989
rect 235715 127961 235749 127989
rect 235777 127961 235811 127989
rect 235839 127961 235887 127989
rect 235577 119175 235887 127961
rect 235577 119147 235625 119175
rect 235653 119147 235687 119175
rect 235715 119147 235749 119175
rect 235777 119147 235811 119175
rect 235839 119147 235887 119175
rect 235577 119113 235887 119147
rect 235577 119085 235625 119113
rect 235653 119085 235687 119113
rect 235715 119085 235749 119113
rect 235777 119085 235811 119113
rect 235839 119085 235887 119113
rect 235577 119051 235887 119085
rect 235577 119023 235625 119051
rect 235653 119023 235687 119051
rect 235715 119023 235749 119051
rect 235777 119023 235811 119051
rect 235839 119023 235887 119051
rect 235577 118989 235887 119023
rect 235577 118961 235625 118989
rect 235653 118961 235687 118989
rect 235715 118961 235749 118989
rect 235777 118961 235811 118989
rect 235839 118961 235887 118989
rect 235577 110175 235887 118961
rect 235577 110147 235625 110175
rect 235653 110147 235687 110175
rect 235715 110147 235749 110175
rect 235777 110147 235811 110175
rect 235839 110147 235887 110175
rect 235577 110113 235887 110147
rect 235577 110085 235625 110113
rect 235653 110085 235687 110113
rect 235715 110085 235749 110113
rect 235777 110085 235811 110113
rect 235839 110085 235887 110113
rect 235577 110051 235887 110085
rect 235577 110023 235625 110051
rect 235653 110023 235687 110051
rect 235715 110023 235749 110051
rect 235777 110023 235811 110051
rect 235839 110023 235887 110051
rect 235577 109989 235887 110023
rect 235577 109961 235625 109989
rect 235653 109961 235687 109989
rect 235715 109961 235749 109989
rect 235777 109961 235811 109989
rect 235839 109961 235887 109989
rect 235577 101175 235887 109961
rect 235577 101147 235625 101175
rect 235653 101147 235687 101175
rect 235715 101147 235749 101175
rect 235777 101147 235811 101175
rect 235839 101147 235887 101175
rect 235577 101113 235887 101147
rect 235577 101085 235625 101113
rect 235653 101085 235687 101113
rect 235715 101085 235749 101113
rect 235777 101085 235811 101113
rect 235839 101085 235887 101113
rect 235577 101051 235887 101085
rect 235577 101023 235625 101051
rect 235653 101023 235687 101051
rect 235715 101023 235749 101051
rect 235777 101023 235811 101051
rect 235839 101023 235887 101051
rect 235577 100989 235887 101023
rect 235577 100961 235625 100989
rect 235653 100961 235687 100989
rect 235715 100961 235749 100989
rect 235777 100961 235811 100989
rect 235839 100961 235887 100989
rect 235577 92175 235887 100961
rect 235577 92147 235625 92175
rect 235653 92147 235687 92175
rect 235715 92147 235749 92175
rect 235777 92147 235811 92175
rect 235839 92147 235887 92175
rect 235577 92113 235887 92147
rect 235577 92085 235625 92113
rect 235653 92085 235687 92113
rect 235715 92085 235749 92113
rect 235777 92085 235811 92113
rect 235839 92085 235887 92113
rect 235577 92051 235887 92085
rect 235577 92023 235625 92051
rect 235653 92023 235687 92051
rect 235715 92023 235749 92051
rect 235777 92023 235811 92051
rect 235839 92023 235887 92051
rect 235577 91989 235887 92023
rect 235577 91961 235625 91989
rect 235653 91961 235687 91989
rect 235715 91961 235749 91989
rect 235777 91961 235811 91989
rect 235839 91961 235887 91989
rect 235577 83175 235887 91961
rect 235577 83147 235625 83175
rect 235653 83147 235687 83175
rect 235715 83147 235749 83175
rect 235777 83147 235811 83175
rect 235839 83147 235887 83175
rect 235577 83113 235887 83147
rect 235577 83085 235625 83113
rect 235653 83085 235687 83113
rect 235715 83085 235749 83113
rect 235777 83085 235811 83113
rect 235839 83085 235887 83113
rect 235577 83051 235887 83085
rect 235577 83023 235625 83051
rect 235653 83023 235687 83051
rect 235715 83023 235749 83051
rect 235777 83023 235811 83051
rect 235839 83023 235887 83051
rect 235577 82989 235887 83023
rect 235577 82961 235625 82989
rect 235653 82961 235687 82989
rect 235715 82961 235749 82989
rect 235777 82961 235811 82989
rect 235839 82961 235887 82989
rect 235577 74175 235887 82961
rect 235577 74147 235625 74175
rect 235653 74147 235687 74175
rect 235715 74147 235749 74175
rect 235777 74147 235811 74175
rect 235839 74147 235887 74175
rect 235577 74113 235887 74147
rect 235577 74085 235625 74113
rect 235653 74085 235687 74113
rect 235715 74085 235749 74113
rect 235777 74085 235811 74113
rect 235839 74085 235887 74113
rect 235577 74051 235887 74085
rect 235577 74023 235625 74051
rect 235653 74023 235687 74051
rect 235715 74023 235749 74051
rect 235777 74023 235811 74051
rect 235839 74023 235887 74051
rect 235577 73989 235887 74023
rect 235577 73961 235625 73989
rect 235653 73961 235687 73989
rect 235715 73961 235749 73989
rect 235777 73961 235811 73989
rect 235839 73961 235887 73989
rect 235577 65175 235887 73961
rect 235577 65147 235625 65175
rect 235653 65147 235687 65175
rect 235715 65147 235749 65175
rect 235777 65147 235811 65175
rect 235839 65147 235887 65175
rect 235577 65113 235887 65147
rect 235577 65085 235625 65113
rect 235653 65085 235687 65113
rect 235715 65085 235749 65113
rect 235777 65085 235811 65113
rect 235839 65085 235887 65113
rect 235577 65051 235887 65085
rect 235577 65023 235625 65051
rect 235653 65023 235687 65051
rect 235715 65023 235749 65051
rect 235777 65023 235811 65051
rect 235839 65023 235887 65051
rect 235577 64989 235887 65023
rect 235577 64961 235625 64989
rect 235653 64961 235687 64989
rect 235715 64961 235749 64989
rect 235777 64961 235811 64989
rect 235839 64961 235887 64989
rect 235577 56175 235887 64961
rect 235577 56147 235625 56175
rect 235653 56147 235687 56175
rect 235715 56147 235749 56175
rect 235777 56147 235811 56175
rect 235839 56147 235887 56175
rect 235577 56113 235887 56147
rect 235577 56085 235625 56113
rect 235653 56085 235687 56113
rect 235715 56085 235749 56113
rect 235777 56085 235811 56113
rect 235839 56085 235887 56113
rect 235577 56051 235887 56085
rect 235577 56023 235625 56051
rect 235653 56023 235687 56051
rect 235715 56023 235749 56051
rect 235777 56023 235811 56051
rect 235839 56023 235887 56051
rect 235577 55989 235887 56023
rect 235577 55961 235625 55989
rect 235653 55961 235687 55989
rect 235715 55961 235749 55989
rect 235777 55961 235811 55989
rect 235839 55961 235887 55989
rect 235577 47175 235887 55961
rect 235577 47147 235625 47175
rect 235653 47147 235687 47175
rect 235715 47147 235749 47175
rect 235777 47147 235811 47175
rect 235839 47147 235887 47175
rect 235577 47113 235887 47147
rect 235577 47085 235625 47113
rect 235653 47085 235687 47113
rect 235715 47085 235749 47113
rect 235777 47085 235811 47113
rect 235839 47085 235887 47113
rect 235577 47051 235887 47085
rect 235577 47023 235625 47051
rect 235653 47023 235687 47051
rect 235715 47023 235749 47051
rect 235777 47023 235811 47051
rect 235839 47023 235887 47051
rect 235577 46989 235887 47023
rect 235577 46961 235625 46989
rect 235653 46961 235687 46989
rect 235715 46961 235749 46989
rect 235777 46961 235811 46989
rect 235839 46961 235887 46989
rect 235577 38175 235887 46961
rect 235577 38147 235625 38175
rect 235653 38147 235687 38175
rect 235715 38147 235749 38175
rect 235777 38147 235811 38175
rect 235839 38147 235887 38175
rect 235577 38113 235887 38147
rect 235577 38085 235625 38113
rect 235653 38085 235687 38113
rect 235715 38085 235749 38113
rect 235777 38085 235811 38113
rect 235839 38085 235887 38113
rect 235577 38051 235887 38085
rect 235577 38023 235625 38051
rect 235653 38023 235687 38051
rect 235715 38023 235749 38051
rect 235777 38023 235811 38051
rect 235839 38023 235887 38051
rect 235577 37989 235887 38023
rect 235577 37961 235625 37989
rect 235653 37961 235687 37989
rect 235715 37961 235749 37989
rect 235777 37961 235811 37989
rect 235839 37961 235887 37989
rect 235577 29175 235887 37961
rect 235577 29147 235625 29175
rect 235653 29147 235687 29175
rect 235715 29147 235749 29175
rect 235777 29147 235811 29175
rect 235839 29147 235887 29175
rect 235577 29113 235887 29147
rect 235577 29085 235625 29113
rect 235653 29085 235687 29113
rect 235715 29085 235749 29113
rect 235777 29085 235811 29113
rect 235839 29085 235887 29113
rect 235577 29051 235887 29085
rect 235577 29023 235625 29051
rect 235653 29023 235687 29051
rect 235715 29023 235749 29051
rect 235777 29023 235811 29051
rect 235839 29023 235887 29051
rect 235577 28989 235887 29023
rect 235577 28961 235625 28989
rect 235653 28961 235687 28989
rect 235715 28961 235749 28989
rect 235777 28961 235811 28989
rect 235839 28961 235887 28989
rect 235577 20175 235887 28961
rect 235577 20147 235625 20175
rect 235653 20147 235687 20175
rect 235715 20147 235749 20175
rect 235777 20147 235811 20175
rect 235839 20147 235887 20175
rect 235577 20113 235887 20147
rect 235577 20085 235625 20113
rect 235653 20085 235687 20113
rect 235715 20085 235749 20113
rect 235777 20085 235811 20113
rect 235839 20085 235887 20113
rect 235577 20051 235887 20085
rect 235577 20023 235625 20051
rect 235653 20023 235687 20051
rect 235715 20023 235749 20051
rect 235777 20023 235811 20051
rect 235839 20023 235887 20051
rect 235577 19989 235887 20023
rect 235577 19961 235625 19989
rect 235653 19961 235687 19989
rect 235715 19961 235749 19989
rect 235777 19961 235811 19989
rect 235839 19961 235887 19989
rect 235577 11175 235887 19961
rect 235577 11147 235625 11175
rect 235653 11147 235687 11175
rect 235715 11147 235749 11175
rect 235777 11147 235811 11175
rect 235839 11147 235887 11175
rect 235577 11113 235887 11147
rect 235577 11085 235625 11113
rect 235653 11085 235687 11113
rect 235715 11085 235749 11113
rect 235777 11085 235811 11113
rect 235839 11085 235887 11113
rect 235577 11051 235887 11085
rect 235577 11023 235625 11051
rect 235653 11023 235687 11051
rect 235715 11023 235749 11051
rect 235777 11023 235811 11051
rect 235839 11023 235887 11051
rect 235577 10989 235887 11023
rect 235577 10961 235625 10989
rect 235653 10961 235687 10989
rect 235715 10961 235749 10989
rect 235777 10961 235811 10989
rect 235839 10961 235887 10989
rect 235577 2175 235887 10961
rect 235577 2147 235625 2175
rect 235653 2147 235687 2175
rect 235715 2147 235749 2175
rect 235777 2147 235811 2175
rect 235839 2147 235887 2175
rect 235577 2113 235887 2147
rect 235577 2085 235625 2113
rect 235653 2085 235687 2113
rect 235715 2085 235749 2113
rect 235777 2085 235811 2113
rect 235839 2085 235887 2113
rect 235577 2051 235887 2085
rect 235577 2023 235625 2051
rect 235653 2023 235687 2051
rect 235715 2023 235749 2051
rect 235777 2023 235811 2051
rect 235839 2023 235887 2051
rect 235577 1989 235887 2023
rect 235577 1961 235625 1989
rect 235653 1961 235687 1989
rect 235715 1961 235749 1989
rect 235777 1961 235811 1989
rect 235839 1961 235887 1989
rect 235577 -80 235887 1961
rect 235577 -108 235625 -80
rect 235653 -108 235687 -80
rect 235715 -108 235749 -80
rect 235777 -108 235811 -80
rect 235839 -108 235887 -80
rect 235577 -142 235887 -108
rect 235577 -170 235625 -142
rect 235653 -170 235687 -142
rect 235715 -170 235749 -142
rect 235777 -170 235811 -142
rect 235839 -170 235887 -142
rect 235577 -204 235887 -170
rect 235577 -232 235625 -204
rect 235653 -232 235687 -204
rect 235715 -232 235749 -204
rect 235777 -232 235811 -204
rect 235839 -232 235887 -204
rect 235577 -266 235887 -232
rect 235577 -294 235625 -266
rect 235653 -294 235687 -266
rect 235715 -294 235749 -266
rect 235777 -294 235811 -266
rect 235839 -294 235887 -266
rect 235577 -822 235887 -294
rect 237437 299086 237747 299134
rect 237437 299058 237485 299086
rect 237513 299058 237547 299086
rect 237575 299058 237609 299086
rect 237637 299058 237671 299086
rect 237699 299058 237747 299086
rect 237437 299024 237747 299058
rect 237437 298996 237485 299024
rect 237513 298996 237547 299024
rect 237575 298996 237609 299024
rect 237637 298996 237671 299024
rect 237699 298996 237747 299024
rect 237437 298962 237747 298996
rect 237437 298934 237485 298962
rect 237513 298934 237547 298962
rect 237575 298934 237609 298962
rect 237637 298934 237671 298962
rect 237699 298934 237747 298962
rect 237437 298900 237747 298934
rect 237437 298872 237485 298900
rect 237513 298872 237547 298900
rect 237575 298872 237609 298900
rect 237637 298872 237671 298900
rect 237699 298872 237747 298900
rect 237437 293175 237747 298872
rect 237437 293147 237485 293175
rect 237513 293147 237547 293175
rect 237575 293147 237609 293175
rect 237637 293147 237671 293175
rect 237699 293147 237747 293175
rect 237437 293113 237747 293147
rect 237437 293085 237485 293113
rect 237513 293085 237547 293113
rect 237575 293085 237609 293113
rect 237637 293085 237671 293113
rect 237699 293085 237747 293113
rect 237437 293051 237747 293085
rect 237437 293023 237485 293051
rect 237513 293023 237547 293051
rect 237575 293023 237609 293051
rect 237637 293023 237671 293051
rect 237699 293023 237747 293051
rect 237437 292989 237747 293023
rect 237437 292961 237485 292989
rect 237513 292961 237547 292989
rect 237575 292961 237609 292989
rect 237637 292961 237671 292989
rect 237699 292961 237747 292989
rect 237437 284175 237747 292961
rect 237437 284147 237485 284175
rect 237513 284147 237547 284175
rect 237575 284147 237609 284175
rect 237637 284147 237671 284175
rect 237699 284147 237747 284175
rect 237437 284113 237747 284147
rect 237437 284085 237485 284113
rect 237513 284085 237547 284113
rect 237575 284085 237609 284113
rect 237637 284085 237671 284113
rect 237699 284085 237747 284113
rect 237437 284051 237747 284085
rect 237437 284023 237485 284051
rect 237513 284023 237547 284051
rect 237575 284023 237609 284051
rect 237637 284023 237671 284051
rect 237699 284023 237747 284051
rect 237437 283989 237747 284023
rect 237437 283961 237485 283989
rect 237513 283961 237547 283989
rect 237575 283961 237609 283989
rect 237637 283961 237671 283989
rect 237699 283961 237747 283989
rect 237437 275175 237747 283961
rect 237437 275147 237485 275175
rect 237513 275147 237547 275175
rect 237575 275147 237609 275175
rect 237637 275147 237671 275175
rect 237699 275147 237747 275175
rect 237437 275113 237747 275147
rect 237437 275085 237485 275113
rect 237513 275085 237547 275113
rect 237575 275085 237609 275113
rect 237637 275085 237671 275113
rect 237699 275085 237747 275113
rect 237437 275051 237747 275085
rect 237437 275023 237485 275051
rect 237513 275023 237547 275051
rect 237575 275023 237609 275051
rect 237637 275023 237671 275051
rect 237699 275023 237747 275051
rect 237437 274989 237747 275023
rect 237437 274961 237485 274989
rect 237513 274961 237547 274989
rect 237575 274961 237609 274989
rect 237637 274961 237671 274989
rect 237699 274961 237747 274989
rect 237437 266175 237747 274961
rect 237437 266147 237485 266175
rect 237513 266147 237547 266175
rect 237575 266147 237609 266175
rect 237637 266147 237671 266175
rect 237699 266147 237747 266175
rect 237437 266113 237747 266147
rect 237437 266085 237485 266113
rect 237513 266085 237547 266113
rect 237575 266085 237609 266113
rect 237637 266085 237671 266113
rect 237699 266085 237747 266113
rect 237437 266051 237747 266085
rect 237437 266023 237485 266051
rect 237513 266023 237547 266051
rect 237575 266023 237609 266051
rect 237637 266023 237671 266051
rect 237699 266023 237747 266051
rect 237437 265989 237747 266023
rect 237437 265961 237485 265989
rect 237513 265961 237547 265989
rect 237575 265961 237609 265989
rect 237637 265961 237671 265989
rect 237699 265961 237747 265989
rect 237437 257175 237747 265961
rect 237437 257147 237485 257175
rect 237513 257147 237547 257175
rect 237575 257147 237609 257175
rect 237637 257147 237671 257175
rect 237699 257147 237747 257175
rect 237437 257113 237747 257147
rect 237437 257085 237485 257113
rect 237513 257085 237547 257113
rect 237575 257085 237609 257113
rect 237637 257085 237671 257113
rect 237699 257085 237747 257113
rect 237437 257051 237747 257085
rect 237437 257023 237485 257051
rect 237513 257023 237547 257051
rect 237575 257023 237609 257051
rect 237637 257023 237671 257051
rect 237699 257023 237747 257051
rect 237437 256989 237747 257023
rect 237437 256961 237485 256989
rect 237513 256961 237547 256989
rect 237575 256961 237609 256989
rect 237637 256961 237671 256989
rect 237699 256961 237747 256989
rect 237437 248175 237747 256961
rect 237437 248147 237485 248175
rect 237513 248147 237547 248175
rect 237575 248147 237609 248175
rect 237637 248147 237671 248175
rect 237699 248147 237747 248175
rect 237437 248113 237747 248147
rect 237437 248085 237485 248113
rect 237513 248085 237547 248113
rect 237575 248085 237609 248113
rect 237637 248085 237671 248113
rect 237699 248085 237747 248113
rect 237437 248051 237747 248085
rect 237437 248023 237485 248051
rect 237513 248023 237547 248051
rect 237575 248023 237609 248051
rect 237637 248023 237671 248051
rect 237699 248023 237747 248051
rect 237437 247989 237747 248023
rect 237437 247961 237485 247989
rect 237513 247961 237547 247989
rect 237575 247961 237609 247989
rect 237637 247961 237671 247989
rect 237699 247961 237747 247989
rect 237437 239175 237747 247961
rect 237437 239147 237485 239175
rect 237513 239147 237547 239175
rect 237575 239147 237609 239175
rect 237637 239147 237671 239175
rect 237699 239147 237747 239175
rect 237437 239113 237747 239147
rect 237437 239085 237485 239113
rect 237513 239085 237547 239113
rect 237575 239085 237609 239113
rect 237637 239085 237671 239113
rect 237699 239085 237747 239113
rect 237437 239051 237747 239085
rect 237437 239023 237485 239051
rect 237513 239023 237547 239051
rect 237575 239023 237609 239051
rect 237637 239023 237671 239051
rect 237699 239023 237747 239051
rect 237437 238989 237747 239023
rect 237437 238961 237485 238989
rect 237513 238961 237547 238989
rect 237575 238961 237609 238989
rect 237637 238961 237671 238989
rect 237699 238961 237747 238989
rect 237437 230175 237747 238961
rect 237437 230147 237485 230175
rect 237513 230147 237547 230175
rect 237575 230147 237609 230175
rect 237637 230147 237671 230175
rect 237699 230147 237747 230175
rect 237437 230113 237747 230147
rect 237437 230085 237485 230113
rect 237513 230085 237547 230113
rect 237575 230085 237609 230113
rect 237637 230085 237671 230113
rect 237699 230085 237747 230113
rect 237437 230051 237747 230085
rect 237437 230023 237485 230051
rect 237513 230023 237547 230051
rect 237575 230023 237609 230051
rect 237637 230023 237671 230051
rect 237699 230023 237747 230051
rect 237437 229989 237747 230023
rect 237437 229961 237485 229989
rect 237513 229961 237547 229989
rect 237575 229961 237609 229989
rect 237637 229961 237671 229989
rect 237699 229961 237747 229989
rect 237437 221175 237747 229961
rect 237437 221147 237485 221175
rect 237513 221147 237547 221175
rect 237575 221147 237609 221175
rect 237637 221147 237671 221175
rect 237699 221147 237747 221175
rect 237437 221113 237747 221147
rect 237437 221085 237485 221113
rect 237513 221085 237547 221113
rect 237575 221085 237609 221113
rect 237637 221085 237671 221113
rect 237699 221085 237747 221113
rect 237437 221051 237747 221085
rect 237437 221023 237485 221051
rect 237513 221023 237547 221051
rect 237575 221023 237609 221051
rect 237637 221023 237671 221051
rect 237699 221023 237747 221051
rect 237437 220989 237747 221023
rect 237437 220961 237485 220989
rect 237513 220961 237547 220989
rect 237575 220961 237609 220989
rect 237637 220961 237671 220989
rect 237699 220961 237747 220989
rect 237437 212175 237747 220961
rect 237437 212147 237485 212175
rect 237513 212147 237547 212175
rect 237575 212147 237609 212175
rect 237637 212147 237671 212175
rect 237699 212147 237747 212175
rect 237437 212113 237747 212147
rect 237437 212085 237485 212113
rect 237513 212085 237547 212113
rect 237575 212085 237609 212113
rect 237637 212085 237671 212113
rect 237699 212085 237747 212113
rect 237437 212051 237747 212085
rect 237437 212023 237485 212051
rect 237513 212023 237547 212051
rect 237575 212023 237609 212051
rect 237637 212023 237671 212051
rect 237699 212023 237747 212051
rect 237437 211989 237747 212023
rect 237437 211961 237485 211989
rect 237513 211961 237547 211989
rect 237575 211961 237609 211989
rect 237637 211961 237671 211989
rect 237699 211961 237747 211989
rect 237437 203175 237747 211961
rect 237437 203147 237485 203175
rect 237513 203147 237547 203175
rect 237575 203147 237609 203175
rect 237637 203147 237671 203175
rect 237699 203147 237747 203175
rect 237437 203113 237747 203147
rect 237437 203085 237485 203113
rect 237513 203085 237547 203113
rect 237575 203085 237609 203113
rect 237637 203085 237671 203113
rect 237699 203085 237747 203113
rect 237437 203051 237747 203085
rect 237437 203023 237485 203051
rect 237513 203023 237547 203051
rect 237575 203023 237609 203051
rect 237637 203023 237671 203051
rect 237699 203023 237747 203051
rect 237437 202989 237747 203023
rect 237437 202961 237485 202989
rect 237513 202961 237547 202989
rect 237575 202961 237609 202989
rect 237637 202961 237671 202989
rect 237699 202961 237747 202989
rect 237437 194175 237747 202961
rect 237437 194147 237485 194175
rect 237513 194147 237547 194175
rect 237575 194147 237609 194175
rect 237637 194147 237671 194175
rect 237699 194147 237747 194175
rect 237437 194113 237747 194147
rect 237437 194085 237485 194113
rect 237513 194085 237547 194113
rect 237575 194085 237609 194113
rect 237637 194085 237671 194113
rect 237699 194085 237747 194113
rect 237437 194051 237747 194085
rect 237437 194023 237485 194051
rect 237513 194023 237547 194051
rect 237575 194023 237609 194051
rect 237637 194023 237671 194051
rect 237699 194023 237747 194051
rect 237437 193989 237747 194023
rect 237437 193961 237485 193989
rect 237513 193961 237547 193989
rect 237575 193961 237609 193989
rect 237637 193961 237671 193989
rect 237699 193961 237747 193989
rect 237437 185175 237747 193961
rect 237437 185147 237485 185175
rect 237513 185147 237547 185175
rect 237575 185147 237609 185175
rect 237637 185147 237671 185175
rect 237699 185147 237747 185175
rect 237437 185113 237747 185147
rect 237437 185085 237485 185113
rect 237513 185085 237547 185113
rect 237575 185085 237609 185113
rect 237637 185085 237671 185113
rect 237699 185085 237747 185113
rect 237437 185051 237747 185085
rect 237437 185023 237485 185051
rect 237513 185023 237547 185051
rect 237575 185023 237609 185051
rect 237637 185023 237671 185051
rect 237699 185023 237747 185051
rect 237437 184989 237747 185023
rect 237437 184961 237485 184989
rect 237513 184961 237547 184989
rect 237575 184961 237609 184989
rect 237637 184961 237671 184989
rect 237699 184961 237747 184989
rect 237437 176175 237747 184961
rect 237437 176147 237485 176175
rect 237513 176147 237547 176175
rect 237575 176147 237609 176175
rect 237637 176147 237671 176175
rect 237699 176147 237747 176175
rect 237437 176113 237747 176147
rect 237437 176085 237485 176113
rect 237513 176085 237547 176113
rect 237575 176085 237609 176113
rect 237637 176085 237671 176113
rect 237699 176085 237747 176113
rect 237437 176051 237747 176085
rect 237437 176023 237485 176051
rect 237513 176023 237547 176051
rect 237575 176023 237609 176051
rect 237637 176023 237671 176051
rect 237699 176023 237747 176051
rect 237437 175989 237747 176023
rect 237437 175961 237485 175989
rect 237513 175961 237547 175989
rect 237575 175961 237609 175989
rect 237637 175961 237671 175989
rect 237699 175961 237747 175989
rect 237437 167175 237747 175961
rect 237437 167147 237485 167175
rect 237513 167147 237547 167175
rect 237575 167147 237609 167175
rect 237637 167147 237671 167175
rect 237699 167147 237747 167175
rect 237437 167113 237747 167147
rect 237437 167085 237485 167113
rect 237513 167085 237547 167113
rect 237575 167085 237609 167113
rect 237637 167085 237671 167113
rect 237699 167085 237747 167113
rect 237437 167051 237747 167085
rect 237437 167023 237485 167051
rect 237513 167023 237547 167051
rect 237575 167023 237609 167051
rect 237637 167023 237671 167051
rect 237699 167023 237747 167051
rect 237437 166989 237747 167023
rect 237437 166961 237485 166989
rect 237513 166961 237547 166989
rect 237575 166961 237609 166989
rect 237637 166961 237671 166989
rect 237699 166961 237747 166989
rect 237437 158175 237747 166961
rect 237437 158147 237485 158175
rect 237513 158147 237547 158175
rect 237575 158147 237609 158175
rect 237637 158147 237671 158175
rect 237699 158147 237747 158175
rect 237437 158113 237747 158147
rect 237437 158085 237485 158113
rect 237513 158085 237547 158113
rect 237575 158085 237609 158113
rect 237637 158085 237671 158113
rect 237699 158085 237747 158113
rect 237437 158051 237747 158085
rect 237437 158023 237485 158051
rect 237513 158023 237547 158051
rect 237575 158023 237609 158051
rect 237637 158023 237671 158051
rect 237699 158023 237747 158051
rect 237437 157989 237747 158023
rect 237437 157961 237485 157989
rect 237513 157961 237547 157989
rect 237575 157961 237609 157989
rect 237637 157961 237671 157989
rect 237699 157961 237747 157989
rect 237437 149175 237747 157961
rect 237437 149147 237485 149175
rect 237513 149147 237547 149175
rect 237575 149147 237609 149175
rect 237637 149147 237671 149175
rect 237699 149147 237747 149175
rect 237437 149113 237747 149147
rect 237437 149085 237485 149113
rect 237513 149085 237547 149113
rect 237575 149085 237609 149113
rect 237637 149085 237671 149113
rect 237699 149085 237747 149113
rect 237437 149051 237747 149085
rect 237437 149023 237485 149051
rect 237513 149023 237547 149051
rect 237575 149023 237609 149051
rect 237637 149023 237671 149051
rect 237699 149023 237747 149051
rect 237437 148989 237747 149023
rect 237437 148961 237485 148989
rect 237513 148961 237547 148989
rect 237575 148961 237609 148989
rect 237637 148961 237671 148989
rect 237699 148961 237747 148989
rect 237437 140175 237747 148961
rect 237437 140147 237485 140175
rect 237513 140147 237547 140175
rect 237575 140147 237609 140175
rect 237637 140147 237671 140175
rect 237699 140147 237747 140175
rect 237437 140113 237747 140147
rect 237437 140085 237485 140113
rect 237513 140085 237547 140113
rect 237575 140085 237609 140113
rect 237637 140085 237671 140113
rect 237699 140085 237747 140113
rect 237437 140051 237747 140085
rect 237437 140023 237485 140051
rect 237513 140023 237547 140051
rect 237575 140023 237609 140051
rect 237637 140023 237671 140051
rect 237699 140023 237747 140051
rect 237437 139989 237747 140023
rect 237437 139961 237485 139989
rect 237513 139961 237547 139989
rect 237575 139961 237609 139989
rect 237637 139961 237671 139989
rect 237699 139961 237747 139989
rect 237437 131175 237747 139961
rect 237437 131147 237485 131175
rect 237513 131147 237547 131175
rect 237575 131147 237609 131175
rect 237637 131147 237671 131175
rect 237699 131147 237747 131175
rect 237437 131113 237747 131147
rect 237437 131085 237485 131113
rect 237513 131085 237547 131113
rect 237575 131085 237609 131113
rect 237637 131085 237671 131113
rect 237699 131085 237747 131113
rect 237437 131051 237747 131085
rect 237437 131023 237485 131051
rect 237513 131023 237547 131051
rect 237575 131023 237609 131051
rect 237637 131023 237671 131051
rect 237699 131023 237747 131051
rect 237437 130989 237747 131023
rect 237437 130961 237485 130989
rect 237513 130961 237547 130989
rect 237575 130961 237609 130989
rect 237637 130961 237671 130989
rect 237699 130961 237747 130989
rect 237437 122175 237747 130961
rect 237437 122147 237485 122175
rect 237513 122147 237547 122175
rect 237575 122147 237609 122175
rect 237637 122147 237671 122175
rect 237699 122147 237747 122175
rect 237437 122113 237747 122147
rect 237437 122085 237485 122113
rect 237513 122085 237547 122113
rect 237575 122085 237609 122113
rect 237637 122085 237671 122113
rect 237699 122085 237747 122113
rect 237437 122051 237747 122085
rect 237437 122023 237485 122051
rect 237513 122023 237547 122051
rect 237575 122023 237609 122051
rect 237637 122023 237671 122051
rect 237699 122023 237747 122051
rect 237437 121989 237747 122023
rect 237437 121961 237485 121989
rect 237513 121961 237547 121989
rect 237575 121961 237609 121989
rect 237637 121961 237671 121989
rect 237699 121961 237747 121989
rect 237437 113175 237747 121961
rect 237437 113147 237485 113175
rect 237513 113147 237547 113175
rect 237575 113147 237609 113175
rect 237637 113147 237671 113175
rect 237699 113147 237747 113175
rect 237437 113113 237747 113147
rect 237437 113085 237485 113113
rect 237513 113085 237547 113113
rect 237575 113085 237609 113113
rect 237637 113085 237671 113113
rect 237699 113085 237747 113113
rect 237437 113051 237747 113085
rect 237437 113023 237485 113051
rect 237513 113023 237547 113051
rect 237575 113023 237609 113051
rect 237637 113023 237671 113051
rect 237699 113023 237747 113051
rect 237437 112989 237747 113023
rect 237437 112961 237485 112989
rect 237513 112961 237547 112989
rect 237575 112961 237609 112989
rect 237637 112961 237671 112989
rect 237699 112961 237747 112989
rect 237437 104175 237747 112961
rect 237437 104147 237485 104175
rect 237513 104147 237547 104175
rect 237575 104147 237609 104175
rect 237637 104147 237671 104175
rect 237699 104147 237747 104175
rect 237437 104113 237747 104147
rect 237437 104085 237485 104113
rect 237513 104085 237547 104113
rect 237575 104085 237609 104113
rect 237637 104085 237671 104113
rect 237699 104085 237747 104113
rect 237437 104051 237747 104085
rect 237437 104023 237485 104051
rect 237513 104023 237547 104051
rect 237575 104023 237609 104051
rect 237637 104023 237671 104051
rect 237699 104023 237747 104051
rect 237437 103989 237747 104023
rect 237437 103961 237485 103989
rect 237513 103961 237547 103989
rect 237575 103961 237609 103989
rect 237637 103961 237671 103989
rect 237699 103961 237747 103989
rect 237437 95175 237747 103961
rect 237437 95147 237485 95175
rect 237513 95147 237547 95175
rect 237575 95147 237609 95175
rect 237637 95147 237671 95175
rect 237699 95147 237747 95175
rect 237437 95113 237747 95147
rect 237437 95085 237485 95113
rect 237513 95085 237547 95113
rect 237575 95085 237609 95113
rect 237637 95085 237671 95113
rect 237699 95085 237747 95113
rect 237437 95051 237747 95085
rect 237437 95023 237485 95051
rect 237513 95023 237547 95051
rect 237575 95023 237609 95051
rect 237637 95023 237671 95051
rect 237699 95023 237747 95051
rect 237437 94989 237747 95023
rect 237437 94961 237485 94989
rect 237513 94961 237547 94989
rect 237575 94961 237609 94989
rect 237637 94961 237671 94989
rect 237699 94961 237747 94989
rect 237437 86175 237747 94961
rect 237437 86147 237485 86175
rect 237513 86147 237547 86175
rect 237575 86147 237609 86175
rect 237637 86147 237671 86175
rect 237699 86147 237747 86175
rect 237437 86113 237747 86147
rect 237437 86085 237485 86113
rect 237513 86085 237547 86113
rect 237575 86085 237609 86113
rect 237637 86085 237671 86113
rect 237699 86085 237747 86113
rect 237437 86051 237747 86085
rect 237437 86023 237485 86051
rect 237513 86023 237547 86051
rect 237575 86023 237609 86051
rect 237637 86023 237671 86051
rect 237699 86023 237747 86051
rect 237437 85989 237747 86023
rect 237437 85961 237485 85989
rect 237513 85961 237547 85989
rect 237575 85961 237609 85989
rect 237637 85961 237671 85989
rect 237699 85961 237747 85989
rect 237437 77175 237747 85961
rect 237437 77147 237485 77175
rect 237513 77147 237547 77175
rect 237575 77147 237609 77175
rect 237637 77147 237671 77175
rect 237699 77147 237747 77175
rect 237437 77113 237747 77147
rect 237437 77085 237485 77113
rect 237513 77085 237547 77113
rect 237575 77085 237609 77113
rect 237637 77085 237671 77113
rect 237699 77085 237747 77113
rect 237437 77051 237747 77085
rect 237437 77023 237485 77051
rect 237513 77023 237547 77051
rect 237575 77023 237609 77051
rect 237637 77023 237671 77051
rect 237699 77023 237747 77051
rect 237437 76989 237747 77023
rect 237437 76961 237485 76989
rect 237513 76961 237547 76989
rect 237575 76961 237609 76989
rect 237637 76961 237671 76989
rect 237699 76961 237747 76989
rect 237437 68175 237747 76961
rect 237437 68147 237485 68175
rect 237513 68147 237547 68175
rect 237575 68147 237609 68175
rect 237637 68147 237671 68175
rect 237699 68147 237747 68175
rect 237437 68113 237747 68147
rect 237437 68085 237485 68113
rect 237513 68085 237547 68113
rect 237575 68085 237609 68113
rect 237637 68085 237671 68113
rect 237699 68085 237747 68113
rect 237437 68051 237747 68085
rect 237437 68023 237485 68051
rect 237513 68023 237547 68051
rect 237575 68023 237609 68051
rect 237637 68023 237671 68051
rect 237699 68023 237747 68051
rect 237437 67989 237747 68023
rect 237437 67961 237485 67989
rect 237513 67961 237547 67989
rect 237575 67961 237609 67989
rect 237637 67961 237671 67989
rect 237699 67961 237747 67989
rect 237437 59175 237747 67961
rect 237437 59147 237485 59175
rect 237513 59147 237547 59175
rect 237575 59147 237609 59175
rect 237637 59147 237671 59175
rect 237699 59147 237747 59175
rect 237437 59113 237747 59147
rect 237437 59085 237485 59113
rect 237513 59085 237547 59113
rect 237575 59085 237609 59113
rect 237637 59085 237671 59113
rect 237699 59085 237747 59113
rect 237437 59051 237747 59085
rect 237437 59023 237485 59051
rect 237513 59023 237547 59051
rect 237575 59023 237609 59051
rect 237637 59023 237671 59051
rect 237699 59023 237747 59051
rect 237437 58989 237747 59023
rect 237437 58961 237485 58989
rect 237513 58961 237547 58989
rect 237575 58961 237609 58989
rect 237637 58961 237671 58989
rect 237699 58961 237747 58989
rect 237437 50175 237747 58961
rect 237437 50147 237485 50175
rect 237513 50147 237547 50175
rect 237575 50147 237609 50175
rect 237637 50147 237671 50175
rect 237699 50147 237747 50175
rect 237437 50113 237747 50147
rect 237437 50085 237485 50113
rect 237513 50085 237547 50113
rect 237575 50085 237609 50113
rect 237637 50085 237671 50113
rect 237699 50085 237747 50113
rect 237437 50051 237747 50085
rect 237437 50023 237485 50051
rect 237513 50023 237547 50051
rect 237575 50023 237609 50051
rect 237637 50023 237671 50051
rect 237699 50023 237747 50051
rect 237437 49989 237747 50023
rect 237437 49961 237485 49989
rect 237513 49961 237547 49989
rect 237575 49961 237609 49989
rect 237637 49961 237671 49989
rect 237699 49961 237747 49989
rect 237437 41175 237747 49961
rect 237437 41147 237485 41175
rect 237513 41147 237547 41175
rect 237575 41147 237609 41175
rect 237637 41147 237671 41175
rect 237699 41147 237747 41175
rect 237437 41113 237747 41147
rect 237437 41085 237485 41113
rect 237513 41085 237547 41113
rect 237575 41085 237609 41113
rect 237637 41085 237671 41113
rect 237699 41085 237747 41113
rect 237437 41051 237747 41085
rect 237437 41023 237485 41051
rect 237513 41023 237547 41051
rect 237575 41023 237609 41051
rect 237637 41023 237671 41051
rect 237699 41023 237747 41051
rect 237437 40989 237747 41023
rect 237437 40961 237485 40989
rect 237513 40961 237547 40989
rect 237575 40961 237609 40989
rect 237637 40961 237671 40989
rect 237699 40961 237747 40989
rect 237437 32175 237747 40961
rect 237437 32147 237485 32175
rect 237513 32147 237547 32175
rect 237575 32147 237609 32175
rect 237637 32147 237671 32175
rect 237699 32147 237747 32175
rect 237437 32113 237747 32147
rect 237437 32085 237485 32113
rect 237513 32085 237547 32113
rect 237575 32085 237609 32113
rect 237637 32085 237671 32113
rect 237699 32085 237747 32113
rect 237437 32051 237747 32085
rect 237437 32023 237485 32051
rect 237513 32023 237547 32051
rect 237575 32023 237609 32051
rect 237637 32023 237671 32051
rect 237699 32023 237747 32051
rect 237437 31989 237747 32023
rect 237437 31961 237485 31989
rect 237513 31961 237547 31989
rect 237575 31961 237609 31989
rect 237637 31961 237671 31989
rect 237699 31961 237747 31989
rect 237437 23175 237747 31961
rect 237437 23147 237485 23175
rect 237513 23147 237547 23175
rect 237575 23147 237609 23175
rect 237637 23147 237671 23175
rect 237699 23147 237747 23175
rect 237437 23113 237747 23147
rect 237437 23085 237485 23113
rect 237513 23085 237547 23113
rect 237575 23085 237609 23113
rect 237637 23085 237671 23113
rect 237699 23085 237747 23113
rect 237437 23051 237747 23085
rect 237437 23023 237485 23051
rect 237513 23023 237547 23051
rect 237575 23023 237609 23051
rect 237637 23023 237671 23051
rect 237699 23023 237747 23051
rect 237437 22989 237747 23023
rect 237437 22961 237485 22989
rect 237513 22961 237547 22989
rect 237575 22961 237609 22989
rect 237637 22961 237671 22989
rect 237699 22961 237747 22989
rect 237437 14175 237747 22961
rect 237437 14147 237485 14175
rect 237513 14147 237547 14175
rect 237575 14147 237609 14175
rect 237637 14147 237671 14175
rect 237699 14147 237747 14175
rect 237437 14113 237747 14147
rect 237437 14085 237485 14113
rect 237513 14085 237547 14113
rect 237575 14085 237609 14113
rect 237637 14085 237671 14113
rect 237699 14085 237747 14113
rect 237437 14051 237747 14085
rect 237437 14023 237485 14051
rect 237513 14023 237547 14051
rect 237575 14023 237609 14051
rect 237637 14023 237671 14051
rect 237699 14023 237747 14051
rect 237437 13989 237747 14023
rect 237437 13961 237485 13989
rect 237513 13961 237547 13989
rect 237575 13961 237609 13989
rect 237637 13961 237671 13989
rect 237699 13961 237747 13989
rect 237437 5175 237747 13961
rect 237437 5147 237485 5175
rect 237513 5147 237547 5175
rect 237575 5147 237609 5175
rect 237637 5147 237671 5175
rect 237699 5147 237747 5175
rect 237437 5113 237747 5147
rect 237437 5085 237485 5113
rect 237513 5085 237547 5113
rect 237575 5085 237609 5113
rect 237637 5085 237671 5113
rect 237699 5085 237747 5113
rect 237437 5051 237747 5085
rect 237437 5023 237485 5051
rect 237513 5023 237547 5051
rect 237575 5023 237609 5051
rect 237637 5023 237671 5051
rect 237699 5023 237747 5051
rect 237437 4989 237747 5023
rect 237437 4961 237485 4989
rect 237513 4961 237547 4989
rect 237575 4961 237609 4989
rect 237637 4961 237671 4989
rect 237699 4961 237747 4989
rect 237437 -560 237747 4961
rect 237437 -588 237485 -560
rect 237513 -588 237547 -560
rect 237575 -588 237609 -560
rect 237637 -588 237671 -560
rect 237699 -588 237747 -560
rect 237437 -622 237747 -588
rect 237437 -650 237485 -622
rect 237513 -650 237547 -622
rect 237575 -650 237609 -622
rect 237637 -650 237671 -622
rect 237699 -650 237747 -622
rect 237437 -684 237747 -650
rect 237437 -712 237485 -684
rect 237513 -712 237547 -684
rect 237575 -712 237609 -684
rect 237637 -712 237671 -684
rect 237699 -712 237747 -684
rect 237437 -746 237747 -712
rect 237437 -774 237485 -746
rect 237513 -774 237547 -746
rect 237575 -774 237609 -746
rect 237637 -774 237671 -746
rect 237699 -774 237747 -746
rect 237437 -822 237747 -774
rect 244577 298606 244887 299134
rect 244577 298578 244625 298606
rect 244653 298578 244687 298606
rect 244715 298578 244749 298606
rect 244777 298578 244811 298606
rect 244839 298578 244887 298606
rect 244577 298544 244887 298578
rect 244577 298516 244625 298544
rect 244653 298516 244687 298544
rect 244715 298516 244749 298544
rect 244777 298516 244811 298544
rect 244839 298516 244887 298544
rect 244577 298482 244887 298516
rect 244577 298454 244625 298482
rect 244653 298454 244687 298482
rect 244715 298454 244749 298482
rect 244777 298454 244811 298482
rect 244839 298454 244887 298482
rect 244577 298420 244887 298454
rect 244577 298392 244625 298420
rect 244653 298392 244687 298420
rect 244715 298392 244749 298420
rect 244777 298392 244811 298420
rect 244839 298392 244887 298420
rect 244577 290175 244887 298392
rect 244577 290147 244625 290175
rect 244653 290147 244687 290175
rect 244715 290147 244749 290175
rect 244777 290147 244811 290175
rect 244839 290147 244887 290175
rect 244577 290113 244887 290147
rect 244577 290085 244625 290113
rect 244653 290085 244687 290113
rect 244715 290085 244749 290113
rect 244777 290085 244811 290113
rect 244839 290085 244887 290113
rect 244577 290051 244887 290085
rect 244577 290023 244625 290051
rect 244653 290023 244687 290051
rect 244715 290023 244749 290051
rect 244777 290023 244811 290051
rect 244839 290023 244887 290051
rect 244577 289989 244887 290023
rect 244577 289961 244625 289989
rect 244653 289961 244687 289989
rect 244715 289961 244749 289989
rect 244777 289961 244811 289989
rect 244839 289961 244887 289989
rect 244577 281175 244887 289961
rect 244577 281147 244625 281175
rect 244653 281147 244687 281175
rect 244715 281147 244749 281175
rect 244777 281147 244811 281175
rect 244839 281147 244887 281175
rect 244577 281113 244887 281147
rect 244577 281085 244625 281113
rect 244653 281085 244687 281113
rect 244715 281085 244749 281113
rect 244777 281085 244811 281113
rect 244839 281085 244887 281113
rect 244577 281051 244887 281085
rect 244577 281023 244625 281051
rect 244653 281023 244687 281051
rect 244715 281023 244749 281051
rect 244777 281023 244811 281051
rect 244839 281023 244887 281051
rect 244577 280989 244887 281023
rect 244577 280961 244625 280989
rect 244653 280961 244687 280989
rect 244715 280961 244749 280989
rect 244777 280961 244811 280989
rect 244839 280961 244887 280989
rect 244577 272175 244887 280961
rect 244577 272147 244625 272175
rect 244653 272147 244687 272175
rect 244715 272147 244749 272175
rect 244777 272147 244811 272175
rect 244839 272147 244887 272175
rect 244577 272113 244887 272147
rect 244577 272085 244625 272113
rect 244653 272085 244687 272113
rect 244715 272085 244749 272113
rect 244777 272085 244811 272113
rect 244839 272085 244887 272113
rect 244577 272051 244887 272085
rect 244577 272023 244625 272051
rect 244653 272023 244687 272051
rect 244715 272023 244749 272051
rect 244777 272023 244811 272051
rect 244839 272023 244887 272051
rect 244577 271989 244887 272023
rect 244577 271961 244625 271989
rect 244653 271961 244687 271989
rect 244715 271961 244749 271989
rect 244777 271961 244811 271989
rect 244839 271961 244887 271989
rect 244577 263175 244887 271961
rect 244577 263147 244625 263175
rect 244653 263147 244687 263175
rect 244715 263147 244749 263175
rect 244777 263147 244811 263175
rect 244839 263147 244887 263175
rect 244577 263113 244887 263147
rect 244577 263085 244625 263113
rect 244653 263085 244687 263113
rect 244715 263085 244749 263113
rect 244777 263085 244811 263113
rect 244839 263085 244887 263113
rect 244577 263051 244887 263085
rect 244577 263023 244625 263051
rect 244653 263023 244687 263051
rect 244715 263023 244749 263051
rect 244777 263023 244811 263051
rect 244839 263023 244887 263051
rect 244577 262989 244887 263023
rect 244577 262961 244625 262989
rect 244653 262961 244687 262989
rect 244715 262961 244749 262989
rect 244777 262961 244811 262989
rect 244839 262961 244887 262989
rect 244577 254175 244887 262961
rect 244577 254147 244625 254175
rect 244653 254147 244687 254175
rect 244715 254147 244749 254175
rect 244777 254147 244811 254175
rect 244839 254147 244887 254175
rect 244577 254113 244887 254147
rect 244577 254085 244625 254113
rect 244653 254085 244687 254113
rect 244715 254085 244749 254113
rect 244777 254085 244811 254113
rect 244839 254085 244887 254113
rect 244577 254051 244887 254085
rect 244577 254023 244625 254051
rect 244653 254023 244687 254051
rect 244715 254023 244749 254051
rect 244777 254023 244811 254051
rect 244839 254023 244887 254051
rect 244577 253989 244887 254023
rect 244577 253961 244625 253989
rect 244653 253961 244687 253989
rect 244715 253961 244749 253989
rect 244777 253961 244811 253989
rect 244839 253961 244887 253989
rect 244577 245175 244887 253961
rect 244577 245147 244625 245175
rect 244653 245147 244687 245175
rect 244715 245147 244749 245175
rect 244777 245147 244811 245175
rect 244839 245147 244887 245175
rect 244577 245113 244887 245147
rect 244577 245085 244625 245113
rect 244653 245085 244687 245113
rect 244715 245085 244749 245113
rect 244777 245085 244811 245113
rect 244839 245085 244887 245113
rect 244577 245051 244887 245085
rect 244577 245023 244625 245051
rect 244653 245023 244687 245051
rect 244715 245023 244749 245051
rect 244777 245023 244811 245051
rect 244839 245023 244887 245051
rect 244577 244989 244887 245023
rect 244577 244961 244625 244989
rect 244653 244961 244687 244989
rect 244715 244961 244749 244989
rect 244777 244961 244811 244989
rect 244839 244961 244887 244989
rect 244577 236175 244887 244961
rect 244577 236147 244625 236175
rect 244653 236147 244687 236175
rect 244715 236147 244749 236175
rect 244777 236147 244811 236175
rect 244839 236147 244887 236175
rect 244577 236113 244887 236147
rect 244577 236085 244625 236113
rect 244653 236085 244687 236113
rect 244715 236085 244749 236113
rect 244777 236085 244811 236113
rect 244839 236085 244887 236113
rect 244577 236051 244887 236085
rect 244577 236023 244625 236051
rect 244653 236023 244687 236051
rect 244715 236023 244749 236051
rect 244777 236023 244811 236051
rect 244839 236023 244887 236051
rect 244577 235989 244887 236023
rect 244577 235961 244625 235989
rect 244653 235961 244687 235989
rect 244715 235961 244749 235989
rect 244777 235961 244811 235989
rect 244839 235961 244887 235989
rect 244577 227175 244887 235961
rect 244577 227147 244625 227175
rect 244653 227147 244687 227175
rect 244715 227147 244749 227175
rect 244777 227147 244811 227175
rect 244839 227147 244887 227175
rect 244577 227113 244887 227147
rect 244577 227085 244625 227113
rect 244653 227085 244687 227113
rect 244715 227085 244749 227113
rect 244777 227085 244811 227113
rect 244839 227085 244887 227113
rect 244577 227051 244887 227085
rect 244577 227023 244625 227051
rect 244653 227023 244687 227051
rect 244715 227023 244749 227051
rect 244777 227023 244811 227051
rect 244839 227023 244887 227051
rect 244577 226989 244887 227023
rect 244577 226961 244625 226989
rect 244653 226961 244687 226989
rect 244715 226961 244749 226989
rect 244777 226961 244811 226989
rect 244839 226961 244887 226989
rect 244577 218175 244887 226961
rect 244577 218147 244625 218175
rect 244653 218147 244687 218175
rect 244715 218147 244749 218175
rect 244777 218147 244811 218175
rect 244839 218147 244887 218175
rect 244577 218113 244887 218147
rect 244577 218085 244625 218113
rect 244653 218085 244687 218113
rect 244715 218085 244749 218113
rect 244777 218085 244811 218113
rect 244839 218085 244887 218113
rect 244577 218051 244887 218085
rect 244577 218023 244625 218051
rect 244653 218023 244687 218051
rect 244715 218023 244749 218051
rect 244777 218023 244811 218051
rect 244839 218023 244887 218051
rect 244577 217989 244887 218023
rect 244577 217961 244625 217989
rect 244653 217961 244687 217989
rect 244715 217961 244749 217989
rect 244777 217961 244811 217989
rect 244839 217961 244887 217989
rect 244577 209175 244887 217961
rect 244577 209147 244625 209175
rect 244653 209147 244687 209175
rect 244715 209147 244749 209175
rect 244777 209147 244811 209175
rect 244839 209147 244887 209175
rect 244577 209113 244887 209147
rect 244577 209085 244625 209113
rect 244653 209085 244687 209113
rect 244715 209085 244749 209113
rect 244777 209085 244811 209113
rect 244839 209085 244887 209113
rect 244577 209051 244887 209085
rect 244577 209023 244625 209051
rect 244653 209023 244687 209051
rect 244715 209023 244749 209051
rect 244777 209023 244811 209051
rect 244839 209023 244887 209051
rect 244577 208989 244887 209023
rect 244577 208961 244625 208989
rect 244653 208961 244687 208989
rect 244715 208961 244749 208989
rect 244777 208961 244811 208989
rect 244839 208961 244887 208989
rect 244577 200175 244887 208961
rect 244577 200147 244625 200175
rect 244653 200147 244687 200175
rect 244715 200147 244749 200175
rect 244777 200147 244811 200175
rect 244839 200147 244887 200175
rect 244577 200113 244887 200147
rect 244577 200085 244625 200113
rect 244653 200085 244687 200113
rect 244715 200085 244749 200113
rect 244777 200085 244811 200113
rect 244839 200085 244887 200113
rect 244577 200051 244887 200085
rect 244577 200023 244625 200051
rect 244653 200023 244687 200051
rect 244715 200023 244749 200051
rect 244777 200023 244811 200051
rect 244839 200023 244887 200051
rect 244577 199989 244887 200023
rect 244577 199961 244625 199989
rect 244653 199961 244687 199989
rect 244715 199961 244749 199989
rect 244777 199961 244811 199989
rect 244839 199961 244887 199989
rect 244577 191175 244887 199961
rect 244577 191147 244625 191175
rect 244653 191147 244687 191175
rect 244715 191147 244749 191175
rect 244777 191147 244811 191175
rect 244839 191147 244887 191175
rect 244577 191113 244887 191147
rect 244577 191085 244625 191113
rect 244653 191085 244687 191113
rect 244715 191085 244749 191113
rect 244777 191085 244811 191113
rect 244839 191085 244887 191113
rect 244577 191051 244887 191085
rect 244577 191023 244625 191051
rect 244653 191023 244687 191051
rect 244715 191023 244749 191051
rect 244777 191023 244811 191051
rect 244839 191023 244887 191051
rect 244577 190989 244887 191023
rect 244577 190961 244625 190989
rect 244653 190961 244687 190989
rect 244715 190961 244749 190989
rect 244777 190961 244811 190989
rect 244839 190961 244887 190989
rect 244577 182175 244887 190961
rect 244577 182147 244625 182175
rect 244653 182147 244687 182175
rect 244715 182147 244749 182175
rect 244777 182147 244811 182175
rect 244839 182147 244887 182175
rect 244577 182113 244887 182147
rect 244577 182085 244625 182113
rect 244653 182085 244687 182113
rect 244715 182085 244749 182113
rect 244777 182085 244811 182113
rect 244839 182085 244887 182113
rect 244577 182051 244887 182085
rect 244577 182023 244625 182051
rect 244653 182023 244687 182051
rect 244715 182023 244749 182051
rect 244777 182023 244811 182051
rect 244839 182023 244887 182051
rect 244577 181989 244887 182023
rect 244577 181961 244625 181989
rect 244653 181961 244687 181989
rect 244715 181961 244749 181989
rect 244777 181961 244811 181989
rect 244839 181961 244887 181989
rect 244577 173175 244887 181961
rect 244577 173147 244625 173175
rect 244653 173147 244687 173175
rect 244715 173147 244749 173175
rect 244777 173147 244811 173175
rect 244839 173147 244887 173175
rect 244577 173113 244887 173147
rect 244577 173085 244625 173113
rect 244653 173085 244687 173113
rect 244715 173085 244749 173113
rect 244777 173085 244811 173113
rect 244839 173085 244887 173113
rect 244577 173051 244887 173085
rect 244577 173023 244625 173051
rect 244653 173023 244687 173051
rect 244715 173023 244749 173051
rect 244777 173023 244811 173051
rect 244839 173023 244887 173051
rect 244577 172989 244887 173023
rect 244577 172961 244625 172989
rect 244653 172961 244687 172989
rect 244715 172961 244749 172989
rect 244777 172961 244811 172989
rect 244839 172961 244887 172989
rect 244577 164175 244887 172961
rect 244577 164147 244625 164175
rect 244653 164147 244687 164175
rect 244715 164147 244749 164175
rect 244777 164147 244811 164175
rect 244839 164147 244887 164175
rect 244577 164113 244887 164147
rect 244577 164085 244625 164113
rect 244653 164085 244687 164113
rect 244715 164085 244749 164113
rect 244777 164085 244811 164113
rect 244839 164085 244887 164113
rect 244577 164051 244887 164085
rect 244577 164023 244625 164051
rect 244653 164023 244687 164051
rect 244715 164023 244749 164051
rect 244777 164023 244811 164051
rect 244839 164023 244887 164051
rect 244577 163989 244887 164023
rect 244577 163961 244625 163989
rect 244653 163961 244687 163989
rect 244715 163961 244749 163989
rect 244777 163961 244811 163989
rect 244839 163961 244887 163989
rect 244577 155175 244887 163961
rect 244577 155147 244625 155175
rect 244653 155147 244687 155175
rect 244715 155147 244749 155175
rect 244777 155147 244811 155175
rect 244839 155147 244887 155175
rect 244577 155113 244887 155147
rect 244577 155085 244625 155113
rect 244653 155085 244687 155113
rect 244715 155085 244749 155113
rect 244777 155085 244811 155113
rect 244839 155085 244887 155113
rect 244577 155051 244887 155085
rect 244577 155023 244625 155051
rect 244653 155023 244687 155051
rect 244715 155023 244749 155051
rect 244777 155023 244811 155051
rect 244839 155023 244887 155051
rect 244577 154989 244887 155023
rect 244577 154961 244625 154989
rect 244653 154961 244687 154989
rect 244715 154961 244749 154989
rect 244777 154961 244811 154989
rect 244839 154961 244887 154989
rect 244577 146175 244887 154961
rect 244577 146147 244625 146175
rect 244653 146147 244687 146175
rect 244715 146147 244749 146175
rect 244777 146147 244811 146175
rect 244839 146147 244887 146175
rect 244577 146113 244887 146147
rect 244577 146085 244625 146113
rect 244653 146085 244687 146113
rect 244715 146085 244749 146113
rect 244777 146085 244811 146113
rect 244839 146085 244887 146113
rect 244577 146051 244887 146085
rect 244577 146023 244625 146051
rect 244653 146023 244687 146051
rect 244715 146023 244749 146051
rect 244777 146023 244811 146051
rect 244839 146023 244887 146051
rect 244577 145989 244887 146023
rect 244577 145961 244625 145989
rect 244653 145961 244687 145989
rect 244715 145961 244749 145989
rect 244777 145961 244811 145989
rect 244839 145961 244887 145989
rect 244577 137175 244887 145961
rect 244577 137147 244625 137175
rect 244653 137147 244687 137175
rect 244715 137147 244749 137175
rect 244777 137147 244811 137175
rect 244839 137147 244887 137175
rect 244577 137113 244887 137147
rect 244577 137085 244625 137113
rect 244653 137085 244687 137113
rect 244715 137085 244749 137113
rect 244777 137085 244811 137113
rect 244839 137085 244887 137113
rect 244577 137051 244887 137085
rect 244577 137023 244625 137051
rect 244653 137023 244687 137051
rect 244715 137023 244749 137051
rect 244777 137023 244811 137051
rect 244839 137023 244887 137051
rect 244577 136989 244887 137023
rect 244577 136961 244625 136989
rect 244653 136961 244687 136989
rect 244715 136961 244749 136989
rect 244777 136961 244811 136989
rect 244839 136961 244887 136989
rect 244577 128175 244887 136961
rect 244577 128147 244625 128175
rect 244653 128147 244687 128175
rect 244715 128147 244749 128175
rect 244777 128147 244811 128175
rect 244839 128147 244887 128175
rect 244577 128113 244887 128147
rect 244577 128085 244625 128113
rect 244653 128085 244687 128113
rect 244715 128085 244749 128113
rect 244777 128085 244811 128113
rect 244839 128085 244887 128113
rect 244577 128051 244887 128085
rect 244577 128023 244625 128051
rect 244653 128023 244687 128051
rect 244715 128023 244749 128051
rect 244777 128023 244811 128051
rect 244839 128023 244887 128051
rect 244577 127989 244887 128023
rect 244577 127961 244625 127989
rect 244653 127961 244687 127989
rect 244715 127961 244749 127989
rect 244777 127961 244811 127989
rect 244839 127961 244887 127989
rect 244577 119175 244887 127961
rect 244577 119147 244625 119175
rect 244653 119147 244687 119175
rect 244715 119147 244749 119175
rect 244777 119147 244811 119175
rect 244839 119147 244887 119175
rect 244577 119113 244887 119147
rect 244577 119085 244625 119113
rect 244653 119085 244687 119113
rect 244715 119085 244749 119113
rect 244777 119085 244811 119113
rect 244839 119085 244887 119113
rect 244577 119051 244887 119085
rect 244577 119023 244625 119051
rect 244653 119023 244687 119051
rect 244715 119023 244749 119051
rect 244777 119023 244811 119051
rect 244839 119023 244887 119051
rect 244577 118989 244887 119023
rect 244577 118961 244625 118989
rect 244653 118961 244687 118989
rect 244715 118961 244749 118989
rect 244777 118961 244811 118989
rect 244839 118961 244887 118989
rect 244577 110175 244887 118961
rect 244577 110147 244625 110175
rect 244653 110147 244687 110175
rect 244715 110147 244749 110175
rect 244777 110147 244811 110175
rect 244839 110147 244887 110175
rect 244577 110113 244887 110147
rect 244577 110085 244625 110113
rect 244653 110085 244687 110113
rect 244715 110085 244749 110113
rect 244777 110085 244811 110113
rect 244839 110085 244887 110113
rect 244577 110051 244887 110085
rect 244577 110023 244625 110051
rect 244653 110023 244687 110051
rect 244715 110023 244749 110051
rect 244777 110023 244811 110051
rect 244839 110023 244887 110051
rect 244577 109989 244887 110023
rect 244577 109961 244625 109989
rect 244653 109961 244687 109989
rect 244715 109961 244749 109989
rect 244777 109961 244811 109989
rect 244839 109961 244887 109989
rect 244577 101175 244887 109961
rect 244577 101147 244625 101175
rect 244653 101147 244687 101175
rect 244715 101147 244749 101175
rect 244777 101147 244811 101175
rect 244839 101147 244887 101175
rect 244577 101113 244887 101147
rect 244577 101085 244625 101113
rect 244653 101085 244687 101113
rect 244715 101085 244749 101113
rect 244777 101085 244811 101113
rect 244839 101085 244887 101113
rect 244577 101051 244887 101085
rect 244577 101023 244625 101051
rect 244653 101023 244687 101051
rect 244715 101023 244749 101051
rect 244777 101023 244811 101051
rect 244839 101023 244887 101051
rect 244577 100989 244887 101023
rect 244577 100961 244625 100989
rect 244653 100961 244687 100989
rect 244715 100961 244749 100989
rect 244777 100961 244811 100989
rect 244839 100961 244887 100989
rect 244577 92175 244887 100961
rect 244577 92147 244625 92175
rect 244653 92147 244687 92175
rect 244715 92147 244749 92175
rect 244777 92147 244811 92175
rect 244839 92147 244887 92175
rect 244577 92113 244887 92147
rect 244577 92085 244625 92113
rect 244653 92085 244687 92113
rect 244715 92085 244749 92113
rect 244777 92085 244811 92113
rect 244839 92085 244887 92113
rect 244577 92051 244887 92085
rect 244577 92023 244625 92051
rect 244653 92023 244687 92051
rect 244715 92023 244749 92051
rect 244777 92023 244811 92051
rect 244839 92023 244887 92051
rect 244577 91989 244887 92023
rect 244577 91961 244625 91989
rect 244653 91961 244687 91989
rect 244715 91961 244749 91989
rect 244777 91961 244811 91989
rect 244839 91961 244887 91989
rect 244577 83175 244887 91961
rect 244577 83147 244625 83175
rect 244653 83147 244687 83175
rect 244715 83147 244749 83175
rect 244777 83147 244811 83175
rect 244839 83147 244887 83175
rect 244577 83113 244887 83147
rect 244577 83085 244625 83113
rect 244653 83085 244687 83113
rect 244715 83085 244749 83113
rect 244777 83085 244811 83113
rect 244839 83085 244887 83113
rect 244577 83051 244887 83085
rect 244577 83023 244625 83051
rect 244653 83023 244687 83051
rect 244715 83023 244749 83051
rect 244777 83023 244811 83051
rect 244839 83023 244887 83051
rect 244577 82989 244887 83023
rect 244577 82961 244625 82989
rect 244653 82961 244687 82989
rect 244715 82961 244749 82989
rect 244777 82961 244811 82989
rect 244839 82961 244887 82989
rect 244577 74175 244887 82961
rect 244577 74147 244625 74175
rect 244653 74147 244687 74175
rect 244715 74147 244749 74175
rect 244777 74147 244811 74175
rect 244839 74147 244887 74175
rect 244577 74113 244887 74147
rect 244577 74085 244625 74113
rect 244653 74085 244687 74113
rect 244715 74085 244749 74113
rect 244777 74085 244811 74113
rect 244839 74085 244887 74113
rect 244577 74051 244887 74085
rect 244577 74023 244625 74051
rect 244653 74023 244687 74051
rect 244715 74023 244749 74051
rect 244777 74023 244811 74051
rect 244839 74023 244887 74051
rect 244577 73989 244887 74023
rect 244577 73961 244625 73989
rect 244653 73961 244687 73989
rect 244715 73961 244749 73989
rect 244777 73961 244811 73989
rect 244839 73961 244887 73989
rect 244577 65175 244887 73961
rect 244577 65147 244625 65175
rect 244653 65147 244687 65175
rect 244715 65147 244749 65175
rect 244777 65147 244811 65175
rect 244839 65147 244887 65175
rect 244577 65113 244887 65147
rect 244577 65085 244625 65113
rect 244653 65085 244687 65113
rect 244715 65085 244749 65113
rect 244777 65085 244811 65113
rect 244839 65085 244887 65113
rect 244577 65051 244887 65085
rect 244577 65023 244625 65051
rect 244653 65023 244687 65051
rect 244715 65023 244749 65051
rect 244777 65023 244811 65051
rect 244839 65023 244887 65051
rect 244577 64989 244887 65023
rect 244577 64961 244625 64989
rect 244653 64961 244687 64989
rect 244715 64961 244749 64989
rect 244777 64961 244811 64989
rect 244839 64961 244887 64989
rect 244577 56175 244887 64961
rect 244577 56147 244625 56175
rect 244653 56147 244687 56175
rect 244715 56147 244749 56175
rect 244777 56147 244811 56175
rect 244839 56147 244887 56175
rect 244577 56113 244887 56147
rect 244577 56085 244625 56113
rect 244653 56085 244687 56113
rect 244715 56085 244749 56113
rect 244777 56085 244811 56113
rect 244839 56085 244887 56113
rect 244577 56051 244887 56085
rect 244577 56023 244625 56051
rect 244653 56023 244687 56051
rect 244715 56023 244749 56051
rect 244777 56023 244811 56051
rect 244839 56023 244887 56051
rect 244577 55989 244887 56023
rect 244577 55961 244625 55989
rect 244653 55961 244687 55989
rect 244715 55961 244749 55989
rect 244777 55961 244811 55989
rect 244839 55961 244887 55989
rect 244577 47175 244887 55961
rect 244577 47147 244625 47175
rect 244653 47147 244687 47175
rect 244715 47147 244749 47175
rect 244777 47147 244811 47175
rect 244839 47147 244887 47175
rect 244577 47113 244887 47147
rect 244577 47085 244625 47113
rect 244653 47085 244687 47113
rect 244715 47085 244749 47113
rect 244777 47085 244811 47113
rect 244839 47085 244887 47113
rect 244577 47051 244887 47085
rect 244577 47023 244625 47051
rect 244653 47023 244687 47051
rect 244715 47023 244749 47051
rect 244777 47023 244811 47051
rect 244839 47023 244887 47051
rect 244577 46989 244887 47023
rect 244577 46961 244625 46989
rect 244653 46961 244687 46989
rect 244715 46961 244749 46989
rect 244777 46961 244811 46989
rect 244839 46961 244887 46989
rect 244577 38175 244887 46961
rect 244577 38147 244625 38175
rect 244653 38147 244687 38175
rect 244715 38147 244749 38175
rect 244777 38147 244811 38175
rect 244839 38147 244887 38175
rect 244577 38113 244887 38147
rect 244577 38085 244625 38113
rect 244653 38085 244687 38113
rect 244715 38085 244749 38113
rect 244777 38085 244811 38113
rect 244839 38085 244887 38113
rect 244577 38051 244887 38085
rect 244577 38023 244625 38051
rect 244653 38023 244687 38051
rect 244715 38023 244749 38051
rect 244777 38023 244811 38051
rect 244839 38023 244887 38051
rect 244577 37989 244887 38023
rect 244577 37961 244625 37989
rect 244653 37961 244687 37989
rect 244715 37961 244749 37989
rect 244777 37961 244811 37989
rect 244839 37961 244887 37989
rect 244577 29175 244887 37961
rect 244577 29147 244625 29175
rect 244653 29147 244687 29175
rect 244715 29147 244749 29175
rect 244777 29147 244811 29175
rect 244839 29147 244887 29175
rect 244577 29113 244887 29147
rect 244577 29085 244625 29113
rect 244653 29085 244687 29113
rect 244715 29085 244749 29113
rect 244777 29085 244811 29113
rect 244839 29085 244887 29113
rect 244577 29051 244887 29085
rect 244577 29023 244625 29051
rect 244653 29023 244687 29051
rect 244715 29023 244749 29051
rect 244777 29023 244811 29051
rect 244839 29023 244887 29051
rect 244577 28989 244887 29023
rect 244577 28961 244625 28989
rect 244653 28961 244687 28989
rect 244715 28961 244749 28989
rect 244777 28961 244811 28989
rect 244839 28961 244887 28989
rect 244577 20175 244887 28961
rect 244577 20147 244625 20175
rect 244653 20147 244687 20175
rect 244715 20147 244749 20175
rect 244777 20147 244811 20175
rect 244839 20147 244887 20175
rect 244577 20113 244887 20147
rect 244577 20085 244625 20113
rect 244653 20085 244687 20113
rect 244715 20085 244749 20113
rect 244777 20085 244811 20113
rect 244839 20085 244887 20113
rect 244577 20051 244887 20085
rect 244577 20023 244625 20051
rect 244653 20023 244687 20051
rect 244715 20023 244749 20051
rect 244777 20023 244811 20051
rect 244839 20023 244887 20051
rect 244577 19989 244887 20023
rect 244577 19961 244625 19989
rect 244653 19961 244687 19989
rect 244715 19961 244749 19989
rect 244777 19961 244811 19989
rect 244839 19961 244887 19989
rect 244577 11175 244887 19961
rect 244577 11147 244625 11175
rect 244653 11147 244687 11175
rect 244715 11147 244749 11175
rect 244777 11147 244811 11175
rect 244839 11147 244887 11175
rect 244577 11113 244887 11147
rect 244577 11085 244625 11113
rect 244653 11085 244687 11113
rect 244715 11085 244749 11113
rect 244777 11085 244811 11113
rect 244839 11085 244887 11113
rect 244577 11051 244887 11085
rect 244577 11023 244625 11051
rect 244653 11023 244687 11051
rect 244715 11023 244749 11051
rect 244777 11023 244811 11051
rect 244839 11023 244887 11051
rect 244577 10989 244887 11023
rect 244577 10961 244625 10989
rect 244653 10961 244687 10989
rect 244715 10961 244749 10989
rect 244777 10961 244811 10989
rect 244839 10961 244887 10989
rect 244577 2175 244887 10961
rect 244577 2147 244625 2175
rect 244653 2147 244687 2175
rect 244715 2147 244749 2175
rect 244777 2147 244811 2175
rect 244839 2147 244887 2175
rect 244577 2113 244887 2147
rect 244577 2085 244625 2113
rect 244653 2085 244687 2113
rect 244715 2085 244749 2113
rect 244777 2085 244811 2113
rect 244839 2085 244887 2113
rect 244577 2051 244887 2085
rect 244577 2023 244625 2051
rect 244653 2023 244687 2051
rect 244715 2023 244749 2051
rect 244777 2023 244811 2051
rect 244839 2023 244887 2051
rect 244577 1989 244887 2023
rect 244577 1961 244625 1989
rect 244653 1961 244687 1989
rect 244715 1961 244749 1989
rect 244777 1961 244811 1989
rect 244839 1961 244887 1989
rect 244577 -80 244887 1961
rect 244577 -108 244625 -80
rect 244653 -108 244687 -80
rect 244715 -108 244749 -80
rect 244777 -108 244811 -80
rect 244839 -108 244887 -80
rect 244577 -142 244887 -108
rect 244577 -170 244625 -142
rect 244653 -170 244687 -142
rect 244715 -170 244749 -142
rect 244777 -170 244811 -142
rect 244839 -170 244887 -142
rect 244577 -204 244887 -170
rect 244577 -232 244625 -204
rect 244653 -232 244687 -204
rect 244715 -232 244749 -204
rect 244777 -232 244811 -204
rect 244839 -232 244887 -204
rect 244577 -266 244887 -232
rect 244577 -294 244625 -266
rect 244653 -294 244687 -266
rect 244715 -294 244749 -266
rect 244777 -294 244811 -266
rect 244839 -294 244887 -266
rect 244577 -822 244887 -294
rect 246437 299086 246747 299134
rect 246437 299058 246485 299086
rect 246513 299058 246547 299086
rect 246575 299058 246609 299086
rect 246637 299058 246671 299086
rect 246699 299058 246747 299086
rect 246437 299024 246747 299058
rect 246437 298996 246485 299024
rect 246513 298996 246547 299024
rect 246575 298996 246609 299024
rect 246637 298996 246671 299024
rect 246699 298996 246747 299024
rect 246437 298962 246747 298996
rect 246437 298934 246485 298962
rect 246513 298934 246547 298962
rect 246575 298934 246609 298962
rect 246637 298934 246671 298962
rect 246699 298934 246747 298962
rect 246437 298900 246747 298934
rect 246437 298872 246485 298900
rect 246513 298872 246547 298900
rect 246575 298872 246609 298900
rect 246637 298872 246671 298900
rect 246699 298872 246747 298900
rect 246437 293175 246747 298872
rect 246437 293147 246485 293175
rect 246513 293147 246547 293175
rect 246575 293147 246609 293175
rect 246637 293147 246671 293175
rect 246699 293147 246747 293175
rect 246437 293113 246747 293147
rect 246437 293085 246485 293113
rect 246513 293085 246547 293113
rect 246575 293085 246609 293113
rect 246637 293085 246671 293113
rect 246699 293085 246747 293113
rect 246437 293051 246747 293085
rect 246437 293023 246485 293051
rect 246513 293023 246547 293051
rect 246575 293023 246609 293051
rect 246637 293023 246671 293051
rect 246699 293023 246747 293051
rect 246437 292989 246747 293023
rect 246437 292961 246485 292989
rect 246513 292961 246547 292989
rect 246575 292961 246609 292989
rect 246637 292961 246671 292989
rect 246699 292961 246747 292989
rect 246437 284175 246747 292961
rect 246437 284147 246485 284175
rect 246513 284147 246547 284175
rect 246575 284147 246609 284175
rect 246637 284147 246671 284175
rect 246699 284147 246747 284175
rect 246437 284113 246747 284147
rect 246437 284085 246485 284113
rect 246513 284085 246547 284113
rect 246575 284085 246609 284113
rect 246637 284085 246671 284113
rect 246699 284085 246747 284113
rect 246437 284051 246747 284085
rect 246437 284023 246485 284051
rect 246513 284023 246547 284051
rect 246575 284023 246609 284051
rect 246637 284023 246671 284051
rect 246699 284023 246747 284051
rect 246437 283989 246747 284023
rect 246437 283961 246485 283989
rect 246513 283961 246547 283989
rect 246575 283961 246609 283989
rect 246637 283961 246671 283989
rect 246699 283961 246747 283989
rect 246437 275175 246747 283961
rect 246437 275147 246485 275175
rect 246513 275147 246547 275175
rect 246575 275147 246609 275175
rect 246637 275147 246671 275175
rect 246699 275147 246747 275175
rect 246437 275113 246747 275147
rect 246437 275085 246485 275113
rect 246513 275085 246547 275113
rect 246575 275085 246609 275113
rect 246637 275085 246671 275113
rect 246699 275085 246747 275113
rect 246437 275051 246747 275085
rect 246437 275023 246485 275051
rect 246513 275023 246547 275051
rect 246575 275023 246609 275051
rect 246637 275023 246671 275051
rect 246699 275023 246747 275051
rect 246437 274989 246747 275023
rect 246437 274961 246485 274989
rect 246513 274961 246547 274989
rect 246575 274961 246609 274989
rect 246637 274961 246671 274989
rect 246699 274961 246747 274989
rect 246437 266175 246747 274961
rect 246437 266147 246485 266175
rect 246513 266147 246547 266175
rect 246575 266147 246609 266175
rect 246637 266147 246671 266175
rect 246699 266147 246747 266175
rect 246437 266113 246747 266147
rect 246437 266085 246485 266113
rect 246513 266085 246547 266113
rect 246575 266085 246609 266113
rect 246637 266085 246671 266113
rect 246699 266085 246747 266113
rect 246437 266051 246747 266085
rect 246437 266023 246485 266051
rect 246513 266023 246547 266051
rect 246575 266023 246609 266051
rect 246637 266023 246671 266051
rect 246699 266023 246747 266051
rect 246437 265989 246747 266023
rect 246437 265961 246485 265989
rect 246513 265961 246547 265989
rect 246575 265961 246609 265989
rect 246637 265961 246671 265989
rect 246699 265961 246747 265989
rect 246437 257175 246747 265961
rect 246437 257147 246485 257175
rect 246513 257147 246547 257175
rect 246575 257147 246609 257175
rect 246637 257147 246671 257175
rect 246699 257147 246747 257175
rect 246437 257113 246747 257147
rect 246437 257085 246485 257113
rect 246513 257085 246547 257113
rect 246575 257085 246609 257113
rect 246637 257085 246671 257113
rect 246699 257085 246747 257113
rect 246437 257051 246747 257085
rect 246437 257023 246485 257051
rect 246513 257023 246547 257051
rect 246575 257023 246609 257051
rect 246637 257023 246671 257051
rect 246699 257023 246747 257051
rect 246437 256989 246747 257023
rect 246437 256961 246485 256989
rect 246513 256961 246547 256989
rect 246575 256961 246609 256989
rect 246637 256961 246671 256989
rect 246699 256961 246747 256989
rect 246437 248175 246747 256961
rect 246437 248147 246485 248175
rect 246513 248147 246547 248175
rect 246575 248147 246609 248175
rect 246637 248147 246671 248175
rect 246699 248147 246747 248175
rect 246437 248113 246747 248147
rect 246437 248085 246485 248113
rect 246513 248085 246547 248113
rect 246575 248085 246609 248113
rect 246637 248085 246671 248113
rect 246699 248085 246747 248113
rect 246437 248051 246747 248085
rect 246437 248023 246485 248051
rect 246513 248023 246547 248051
rect 246575 248023 246609 248051
rect 246637 248023 246671 248051
rect 246699 248023 246747 248051
rect 246437 247989 246747 248023
rect 246437 247961 246485 247989
rect 246513 247961 246547 247989
rect 246575 247961 246609 247989
rect 246637 247961 246671 247989
rect 246699 247961 246747 247989
rect 246437 239175 246747 247961
rect 246437 239147 246485 239175
rect 246513 239147 246547 239175
rect 246575 239147 246609 239175
rect 246637 239147 246671 239175
rect 246699 239147 246747 239175
rect 246437 239113 246747 239147
rect 246437 239085 246485 239113
rect 246513 239085 246547 239113
rect 246575 239085 246609 239113
rect 246637 239085 246671 239113
rect 246699 239085 246747 239113
rect 246437 239051 246747 239085
rect 246437 239023 246485 239051
rect 246513 239023 246547 239051
rect 246575 239023 246609 239051
rect 246637 239023 246671 239051
rect 246699 239023 246747 239051
rect 246437 238989 246747 239023
rect 246437 238961 246485 238989
rect 246513 238961 246547 238989
rect 246575 238961 246609 238989
rect 246637 238961 246671 238989
rect 246699 238961 246747 238989
rect 246437 230175 246747 238961
rect 246437 230147 246485 230175
rect 246513 230147 246547 230175
rect 246575 230147 246609 230175
rect 246637 230147 246671 230175
rect 246699 230147 246747 230175
rect 246437 230113 246747 230147
rect 246437 230085 246485 230113
rect 246513 230085 246547 230113
rect 246575 230085 246609 230113
rect 246637 230085 246671 230113
rect 246699 230085 246747 230113
rect 246437 230051 246747 230085
rect 246437 230023 246485 230051
rect 246513 230023 246547 230051
rect 246575 230023 246609 230051
rect 246637 230023 246671 230051
rect 246699 230023 246747 230051
rect 246437 229989 246747 230023
rect 246437 229961 246485 229989
rect 246513 229961 246547 229989
rect 246575 229961 246609 229989
rect 246637 229961 246671 229989
rect 246699 229961 246747 229989
rect 246437 221175 246747 229961
rect 246437 221147 246485 221175
rect 246513 221147 246547 221175
rect 246575 221147 246609 221175
rect 246637 221147 246671 221175
rect 246699 221147 246747 221175
rect 246437 221113 246747 221147
rect 246437 221085 246485 221113
rect 246513 221085 246547 221113
rect 246575 221085 246609 221113
rect 246637 221085 246671 221113
rect 246699 221085 246747 221113
rect 246437 221051 246747 221085
rect 246437 221023 246485 221051
rect 246513 221023 246547 221051
rect 246575 221023 246609 221051
rect 246637 221023 246671 221051
rect 246699 221023 246747 221051
rect 246437 220989 246747 221023
rect 246437 220961 246485 220989
rect 246513 220961 246547 220989
rect 246575 220961 246609 220989
rect 246637 220961 246671 220989
rect 246699 220961 246747 220989
rect 246437 212175 246747 220961
rect 246437 212147 246485 212175
rect 246513 212147 246547 212175
rect 246575 212147 246609 212175
rect 246637 212147 246671 212175
rect 246699 212147 246747 212175
rect 246437 212113 246747 212147
rect 246437 212085 246485 212113
rect 246513 212085 246547 212113
rect 246575 212085 246609 212113
rect 246637 212085 246671 212113
rect 246699 212085 246747 212113
rect 246437 212051 246747 212085
rect 246437 212023 246485 212051
rect 246513 212023 246547 212051
rect 246575 212023 246609 212051
rect 246637 212023 246671 212051
rect 246699 212023 246747 212051
rect 246437 211989 246747 212023
rect 246437 211961 246485 211989
rect 246513 211961 246547 211989
rect 246575 211961 246609 211989
rect 246637 211961 246671 211989
rect 246699 211961 246747 211989
rect 246437 203175 246747 211961
rect 246437 203147 246485 203175
rect 246513 203147 246547 203175
rect 246575 203147 246609 203175
rect 246637 203147 246671 203175
rect 246699 203147 246747 203175
rect 246437 203113 246747 203147
rect 246437 203085 246485 203113
rect 246513 203085 246547 203113
rect 246575 203085 246609 203113
rect 246637 203085 246671 203113
rect 246699 203085 246747 203113
rect 246437 203051 246747 203085
rect 246437 203023 246485 203051
rect 246513 203023 246547 203051
rect 246575 203023 246609 203051
rect 246637 203023 246671 203051
rect 246699 203023 246747 203051
rect 246437 202989 246747 203023
rect 246437 202961 246485 202989
rect 246513 202961 246547 202989
rect 246575 202961 246609 202989
rect 246637 202961 246671 202989
rect 246699 202961 246747 202989
rect 246437 194175 246747 202961
rect 246437 194147 246485 194175
rect 246513 194147 246547 194175
rect 246575 194147 246609 194175
rect 246637 194147 246671 194175
rect 246699 194147 246747 194175
rect 246437 194113 246747 194147
rect 246437 194085 246485 194113
rect 246513 194085 246547 194113
rect 246575 194085 246609 194113
rect 246637 194085 246671 194113
rect 246699 194085 246747 194113
rect 246437 194051 246747 194085
rect 246437 194023 246485 194051
rect 246513 194023 246547 194051
rect 246575 194023 246609 194051
rect 246637 194023 246671 194051
rect 246699 194023 246747 194051
rect 246437 193989 246747 194023
rect 246437 193961 246485 193989
rect 246513 193961 246547 193989
rect 246575 193961 246609 193989
rect 246637 193961 246671 193989
rect 246699 193961 246747 193989
rect 246437 185175 246747 193961
rect 246437 185147 246485 185175
rect 246513 185147 246547 185175
rect 246575 185147 246609 185175
rect 246637 185147 246671 185175
rect 246699 185147 246747 185175
rect 246437 185113 246747 185147
rect 246437 185085 246485 185113
rect 246513 185085 246547 185113
rect 246575 185085 246609 185113
rect 246637 185085 246671 185113
rect 246699 185085 246747 185113
rect 246437 185051 246747 185085
rect 246437 185023 246485 185051
rect 246513 185023 246547 185051
rect 246575 185023 246609 185051
rect 246637 185023 246671 185051
rect 246699 185023 246747 185051
rect 246437 184989 246747 185023
rect 246437 184961 246485 184989
rect 246513 184961 246547 184989
rect 246575 184961 246609 184989
rect 246637 184961 246671 184989
rect 246699 184961 246747 184989
rect 246437 176175 246747 184961
rect 246437 176147 246485 176175
rect 246513 176147 246547 176175
rect 246575 176147 246609 176175
rect 246637 176147 246671 176175
rect 246699 176147 246747 176175
rect 246437 176113 246747 176147
rect 246437 176085 246485 176113
rect 246513 176085 246547 176113
rect 246575 176085 246609 176113
rect 246637 176085 246671 176113
rect 246699 176085 246747 176113
rect 246437 176051 246747 176085
rect 246437 176023 246485 176051
rect 246513 176023 246547 176051
rect 246575 176023 246609 176051
rect 246637 176023 246671 176051
rect 246699 176023 246747 176051
rect 246437 175989 246747 176023
rect 246437 175961 246485 175989
rect 246513 175961 246547 175989
rect 246575 175961 246609 175989
rect 246637 175961 246671 175989
rect 246699 175961 246747 175989
rect 246437 167175 246747 175961
rect 246437 167147 246485 167175
rect 246513 167147 246547 167175
rect 246575 167147 246609 167175
rect 246637 167147 246671 167175
rect 246699 167147 246747 167175
rect 246437 167113 246747 167147
rect 246437 167085 246485 167113
rect 246513 167085 246547 167113
rect 246575 167085 246609 167113
rect 246637 167085 246671 167113
rect 246699 167085 246747 167113
rect 246437 167051 246747 167085
rect 246437 167023 246485 167051
rect 246513 167023 246547 167051
rect 246575 167023 246609 167051
rect 246637 167023 246671 167051
rect 246699 167023 246747 167051
rect 246437 166989 246747 167023
rect 246437 166961 246485 166989
rect 246513 166961 246547 166989
rect 246575 166961 246609 166989
rect 246637 166961 246671 166989
rect 246699 166961 246747 166989
rect 246437 158175 246747 166961
rect 246437 158147 246485 158175
rect 246513 158147 246547 158175
rect 246575 158147 246609 158175
rect 246637 158147 246671 158175
rect 246699 158147 246747 158175
rect 246437 158113 246747 158147
rect 246437 158085 246485 158113
rect 246513 158085 246547 158113
rect 246575 158085 246609 158113
rect 246637 158085 246671 158113
rect 246699 158085 246747 158113
rect 246437 158051 246747 158085
rect 246437 158023 246485 158051
rect 246513 158023 246547 158051
rect 246575 158023 246609 158051
rect 246637 158023 246671 158051
rect 246699 158023 246747 158051
rect 246437 157989 246747 158023
rect 246437 157961 246485 157989
rect 246513 157961 246547 157989
rect 246575 157961 246609 157989
rect 246637 157961 246671 157989
rect 246699 157961 246747 157989
rect 246437 149175 246747 157961
rect 246437 149147 246485 149175
rect 246513 149147 246547 149175
rect 246575 149147 246609 149175
rect 246637 149147 246671 149175
rect 246699 149147 246747 149175
rect 246437 149113 246747 149147
rect 246437 149085 246485 149113
rect 246513 149085 246547 149113
rect 246575 149085 246609 149113
rect 246637 149085 246671 149113
rect 246699 149085 246747 149113
rect 246437 149051 246747 149085
rect 246437 149023 246485 149051
rect 246513 149023 246547 149051
rect 246575 149023 246609 149051
rect 246637 149023 246671 149051
rect 246699 149023 246747 149051
rect 246437 148989 246747 149023
rect 246437 148961 246485 148989
rect 246513 148961 246547 148989
rect 246575 148961 246609 148989
rect 246637 148961 246671 148989
rect 246699 148961 246747 148989
rect 246437 140175 246747 148961
rect 246437 140147 246485 140175
rect 246513 140147 246547 140175
rect 246575 140147 246609 140175
rect 246637 140147 246671 140175
rect 246699 140147 246747 140175
rect 246437 140113 246747 140147
rect 246437 140085 246485 140113
rect 246513 140085 246547 140113
rect 246575 140085 246609 140113
rect 246637 140085 246671 140113
rect 246699 140085 246747 140113
rect 246437 140051 246747 140085
rect 246437 140023 246485 140051
rect 246513 140023 246547 140051
rect 246575 140023 246609 140051
rect 246637 140023 246671 140051
rect 246699 140023 246747 140051
rect 246437 139989 246747 140023
rect 246437 139961 246485 139989
rect 246513 139961 246547 139989
rect 246575 139961 246609 139989
rect 246637 139961 246671 139989
rect 246699 139961 246747 139989
rect 246437 131175 246747 139961
rect 246437 131147 246485 131175
rect 246513 131147 246547 131175
rect 246575 131147 246609 131175
rect 246637 131147 246671 131175
rect 246699 131147 246747 131175
rect 246437 131113 246747 131147
rect 246437 131085 246485 131113
rect 246513 131085 246547 131113
rect 246575 131085 246609 131113
rect 246637 131085 246671 131113
rect 246699 131085 246747 131113
rect 246437 131051 246747 131085
rect 246437 131023 246485 131051
rect 246513 131023 246547 131051
rect 246575 131023 246609 131051
rect 246637 131023 246671 131051
rect 246699 131023 246747 131051
rect 246437 130989 246747 131023
rect 246437 130961 246485 130989
rect 246513 130961 246547 130989
rect 246575 130961 246609 130989
rect 246637 130961 246671 130989
rect 246699 130961 246747 130989
rect 246437 122175 246747 130961
rect 246437 122147 246485 122175
rect 246513 122147 246547 122175
rect 246575 122147 246609 122175
rect 246637 122147 246671 122175
rect 246699 122147 246747 122175
rect 246437 122113 246747 122147
rect 246437 122085 246485 122113
rect 246513 122085 246547 122113
rect 246575 122085 246609 122113
rect 246637 122085 246671 122113
rect 246699 122085 246747 122113
rect 246437 122051 246747 122085
rect 246437 122023 246485 122051
rect 246513 122023 246547 122051
rect 246575 122023 246609 122051
rect 246637 122023 246671 122051
rect 246699 122023 246747 122051
rect 246437 121989 246747 122023
rect 246437 121961 246485 121989
rect 246513 121961 246547 121989
rect 246575 121961 246609 121989
rect 246637 121961 246671 121989
rect 246699 121961 246747 121989
rect 246437 113175 246747 121961
rect 246437 113147 246485 113175
rect 246513 113147 246547 113175
rect 246575 113147 246609 113175
rect 246637 113147 246671 113175
rect 246699 113147 246747 113175
rect 246437 113113 246747 113147
rect 246437 113085 246485 113113
rect 246513 113085 246547 113113
rect 246575 113085 246609 113113
rect 246637 113085 246671 113113
rect 246699 113085 246747 113113
rect 246437 113051 246747 113085
rect 246437 113023 246485 113051
rect 246513 113023 246547 113051
rect 246575 113023 246609 113051
rect 246637 113023 246671 113051
rect 246699 113023 246747 113051
rect 246437 112989 246747 113023
rect 246437 112961 246485 112989
rect 246513 112961 246547 112989
rect 246575 112961 246609 112989
rect 246637 112961 246671 112989
rect 246699 112961 246747 112989
rect 246437 104175 246747 112961
rect 246437 104147 246485 104175
rect 246513 104147 246547 104175
rect 246575 104147 246609 104175
rect 246637 104147 246671 104175
rect 246699 104147 246747 104175
rect 246437 104113 246747 104147
rect 246437 104085 246485 104113
rect 246513 104085 246547 104113
rect 246575 104085 246609 104113
rect 246637 104085 246671 104113
rect 246699 104085 246747 104113
rect 246437 104051 246747 104085
rect 246437 104023 246485 104051
rect 246513 104023 246547 104051
rect 246575 104023 246609 104051
rect 246637 104023 246671 104051
rect 246699 104023 246747 104051
rect 246437 103989 246747 104023
rect 246437 103961 246485 103989
rect 246513 103961 246547 103989
rect 246575 103961 246609 103989
rect 246637 103961 246671 103989
rect 246699 103961 246747 103989
rect 246437 95175 246747 103961
rect 246437 95147 246485 95175
rect 246513 95147 246547 95175
rect 246575 95147 246609 95175
rect 246637 95147 246671 95175
rect 246699 95147 246747 95175
rect 246437 95113 246747 95147
rect 246437 95085 246485 95113
rect 246513 95085 246547 95113
rect 246575 95085 246609 95113
rect 246637 95085 246671 95113
rect 246699 95085 246747 95113
rect 246437 95051 246747 95085
rect 246437 95023 246485 95051
rect 246513 95023 246547 95051
rect 246575 95023 246609 95051
rect 246637 95023 246671 95051
rect 246699 95023 246747 95051
rect 246437 94989 246747 95023
rect 246437 94961 246485 94989
rect 246513 94961 246547 94989
rect 246575 94961 246609 94989
rect 246637 94961 246671 94989
rect 246699 94961 246747 94989
rect 246437 86175 246747 94961
rect 246437 86147 246485 86175
rect 246513 86147 246547 86175
rect 246575 86147 246609 86175
rect 246637 86147 246671 86175
rect 246699 86147 246747 86175
rect 246437 86113 246747 86147
rect 246437 86085 246485 86113
rect 246513 86085 246547 86113
rect 246575 86085 246609 86113
rect 246637 86085 246671 86113
rect 246699 86085 246747 86113
rect 246437 86051 246747 86085
rect 246437 86023 246485 86051
rect 246513 86023 246547 86051
rect 246575 86023 246609 86051
rect 246637 86023 246671 86051
rect 246699 86023 246747 86051
rect 246437 85989 246747 86023
rect 246437 85961 246485 85989
rect 246513 85961 246547 85989
rect 246575 85961 246609 85989
rect 246637 85961 246671 85989
rect 246699 85961 246747 85989
rect 246437 77175 246747 85961
rect 246437 77147 246485 77175
rect 246513 77147 246547 77175
rect 246575 77147 246609 77175
rect 246637 77147 246671 77175
rect 246699 77147 246747 77175
rect 246437 77113 246747 77147
rect 246437 77085 246485 77113
rect 246513 77085 246547 77113
rect 246575 77085 246609 77113
rect 246637 77085 246671 77113
rect 246699 77085 246747 77113
rect 246437 77051 246747 77085
rect 246437 77023 246485 77051
rect 246513 77023 246547 77051
rect 246575 77023 246609 77051
rect 246637 77023 246671 77051
rect 246699 77023 246747 77051
rect 246437 76989 246747 77023
rect 246437 76961 246485 76989
rect 246513 76961 246547 76989
rect 246575 76961 246609 76989
rect 246637 76961 246671 76989
rect 246699 76961 246747 76989
rect 246437 68175 246747 76961
rect 246437 68147 246485 68175
rect 246513 68147 246547 68175
rect 246575 68147 246609 68175
rect 246637 68147 246671 68175
rect 246699 68147 246747 68175
rect 246437 68113 246747 68147
rect 246437 68085 246485 68113
rect 246513 68085 246547 68113
rect 246575 68085 246609 68113
rect 246637 68085 246671 68113
rect 246699 68085 246747 68113
rect 246437 68051 246747 68085
rect 246437 68023 246485 68051
rect 246513 68023 246547 68051
rect 246575 68023 246609 68051
rect 246637 68023 246671 68051
rect 246699 68023 246747 68051
rect 246437 67989 246747 68023
rect 246437 67961 246485 67989
rect 246513 67961 246547 67989
rect 246575 67961 246609 67989
rect 246637 67961 246671 67989
rect 246699 67961 246747 67989
rect 246437 59175 246747 67961
rect 246437 59147 246485 59175
rect 246513 59147 246547 59175
rect 246575 59147 246609 59175
rect 246637 59147 246671 59175
rect 246699 59147 246747 59175
rect 246437 59113 246747 59147
rect 246437 59085 246485 59113
rect 246513 59085 246547 59113
rect 246575 59085 246609 59113
rect 246637 59085 246671 59113
rect 246699 59085 246747 59113
rect 246437 59051 246747 59085
rect 246437 59023 246485 59051
rect 246513 59023 246547 59051
rect 246575 59023 246609 59051
rect 246637 59023 246671 59051
rect 246699 59023 246747 59051
rect 246437 58989 246747 59023
rect 246437 58961 246485 58989
rect 246513 58961 246547 58989
rect 246575 58961 246609 58989
rect 246637 58961 246671 58989
rect 246699 58961 246747 58989
rect 246437 50175 246747 58961
rect 246437 50147 246485 50175
rect 246513 50147 246547 50175
rect 246575 50147 246609 50175
rect 246637 50147 246671 50175
rect 246699 50147 246747 50175
rect 246437 50113 246747 50147
rect 246437 50085 246485 50113
rect 246513 50085 246547 50113
rect 246575 50085 246609 50113
rect 246637 50085 246671 50113
rect 246699 50085 246747 50113
rect 246437 50051 246747 50085
rect 246437 50023 246485 50051
rect 246513 50023 246547 50051
rect 246575 50023 246609 50051
rect 246637 50023 246671 50051
rect 246699 50023 246747 50051
rect 246437 49989 246747 50023
rect 246437 49961 246485 49989
rect 246513 49961 246547 49989
rect 246575 49961 246609 49989
rect 246637 49961 246671 49989
rect 246699 49961 246747 49989
rect 246437 41175 246747 49961
rect 246437 41147 246485 41175
rect 246513 41147 246547 41175
rect 246575 41147 246609 41175
rect 246637 41147 246671 41175
rect 246699 41147 246747 41175
rect 246437 41113 246747 41147
rect 246437 41085 246485 41113
rect 246513 41085 246547 41113
rect 246575 41085 246609 41113
rect 246637 41085 246671 41113
rect 246699 41085 246747 41113
rect 246437 41051 246747 41085
rect 246437 41023 246485 41051
rect 246513 41023 246547 41051
rect 246575 41023 246609 41051
rect 246637 41023 246671 41051
rect 246699 41023 246747 41051
rect 246437 40989 246747 41023
rect 246437 40961 246485 40989
rect 246513 40961 246547 40989
rect 246575 40961 246609 40989
rect 246637 40961 246671 40989
rect 246699 40961 246747 40989
rect 246437 32175 246747 40961
rect 246437 32147 246485 32175
rect 246513 32147 246547 32175
rect 246575 32147 246609 32175
rect 246637 32147 246671 32175
rect 246699 32147 246747 32175
rect 246437 32113 246747 32147
rect 246437 32085 246485 32113
rect 246513 32085 246547 32113
rect 246575 32085 246609 32113
rect 246637 32085 246671 32113
rect 246699 32085 246747 32113
rect 246437 32051 246747 32085
rect 246437 32023 246485 32051
rect 246513 32023 246547 32051
rect 246575 32023 246609 32051
rect 246637 32023 246671 32051
rect 246699 32023 246747 32051
rect 246437 31989 246747 32023
rect 246437 31961 246485 31989
rect 246513 31961 246547 31989
rect 246575 31961 246609 31989
rect 246637 31961 246671 31989
rect 246699 31961 246747 31989
rect 246437 23175 246747 31961
rect 246437 23147 246485 23175
rect 246513 23147 246547 23175
rect 246575 23147 246609 23175
rect 246637 23147 246671 23175
rect 246699 23147 246747 23175
rect 246437 23113 246747 23147
rect 246437 23085 246485 23113
rect 246513 23085 246547 23113
rect 246575 23085 246609 23113
rect 246637 23085 246671 23113
rect 246699 23085 246747 23113
rect 246437 23051 246747 23085
rect 246437 23023 246485 23051
rect 246513 23023 246547 23051
rect 246575 23023 246609 23051
rect 246637 23023 246671 23051
rect 246699 23023 246747 23051
rect 246437 22989 246747 23023
rect 246437 22961 246485 22989
rect 246513 22961 246547 22989
rect 246575 22961 246609 22989
rect 246637 22961 246671 22989
rect 246699 22961 246747 22989
rect 246437 14175 246747 22961
rect 246437 14147 246485 14175
rect 246513 14147 246547 14175
rect 246575 14147 246609 14175
rect 246637 14147 246671 14175
rect 246699 14147 246747 14175
rect 246437 14113 246747 14147
rect 246437 14085 246485 14113
rect 246513 14085 246547 14113
rect 246575 14085 246609 14113
rect 246637 14085 246671 14113
rect 246699 14085 246747 14113
rect 246437 14051 246747 14085
rect 246437 14023 246485 14051
rect 246513 14023 246547 14051
rect 246575 14023 246609 14051
rect 246637 14023 246671 14051
rect 246699 14023 246747 14051
rect 246437 13989 246747 14023
rect 246437 13961 246485 13989
rect 246513 13961 246547 13989
rect 246575 13961 246609 13989
rect 246637 13961 246671 13989
rect 246699 13961 246747 13989
rect 246437 5175 246747 13961
rect 246437 5147 246485 5175
rect 246513 5147 246547 5175
rect 246575 5147 246609 5175
rect 246637 5147 246671 5175
rect 246699 5147 246747 5175
rect 246437 5113 246747 5147
rect 246437 5085 246485 5113
rect 246513 5085 246547 5113
rect 246575 5085 246609 5113
rect 246637 5085 246671 5113
rect 246699 5085 246747 5113
rect 246437 5051 246747 5085
rect 246437 5023 246485 5051
rect 246513 5023 246547 5051
rect 246575 5023 246609 5051
rect 246637 5023 246671 5051
rect 246699 5023 246747 5051
rect 246437 4989 246747 5023
rect 246437 4961 246485 4989
rect 246513 4961 246547 4989
rect 246575 4961 246609 4989
rect 246637 4961 246671 4989
rect 246699 4961 246747 4989
rect 246437 -560 246747 4961
rect 246437 -588 246485 -560
rect 246513 -588 246547 -560
rect 246575 -588 246609 -560
rect 246637 -588 246671 -560
rect 246699 -588 246747 -560
rect 246437 -622 246747 -588
rect 246437 -650 246485 -622
rect 246513 -650 246547 -622
rect 246575 -650 246609 -622
rect 246637 -650 246671 -622
rect 246699 -650 246747 -622
rect 246437 -684 246747 -650
rect 246437 -712 246485 -684
rect 246513 -712 246547 -684
rect 246575 -712 246609 -684
rect 246637 -712 246671 -684
rect 246699 -712 246747 -684
rect 246437 -746 246747 -712
rect 246437 -774 246485 -746
rect 246513 -774 246547 -746
rect 246575 -774 246609 -746
rect 246637 -774 246671 -746
rect 246699 -774 246747 -746
rect 246437 -822 246747 -774
rect 253577 298606 253887 299134
rect 253577 298578 253625 298606
rect 253653 298578 253687 298606
rect 253715 298578 253749 298606
rect 253777 298578 253811 298606
rect 253839 298578 253887 298606
rect 253577 298544 253887 298578
rect 253577 298516 253625 298544
rect 253653 298516 253687 298544
rect 253715 298516 253749 298544
rect 253777 298516 253811 298544
rect 253839 298516 253887 298544
rect 253577 298482 253887 298516
rect 253577 298454 253625 298482
rect 253653 298454 253687 298482
rect 253715 298454 253749 298482
rect 253777 298454 253811 298482
rect 253839 298454 253887 298482
rect 253577 298420 253887 298454
rect 253577 298392 253625 298420
rect 253653 298392 253687 298420
rect 253715 298392 253749 298420
rect 253777 298392 253811 298420
rect 253839 298392 253887 298420
rect 253577 290175 253887 298392
rect 253577 290147 253625 290175
rect 253653 290147 253687 290175
rect 253715 290147 253749 290175
rect 253777 290147 253811 290175
rect 253839 290147 253887 290175
rect 253577 290113 253887 290147
rect 253577 290085 253625 290113
rect 253653 290085 253687 290113
rect 253715 290085 253749 290113
rect 253777 290085 253811 290113
rect 253839 290085 253887 290113
rect 253577 290051 253887 290085
rect 253577 290023 253625 290051
rect 253653 290023 253687 290051
rect 253715 290023 253749 290051
rect 253777 290023 253811 290051
rect 253839 290023 253887 290051
rect 253577 289989 253887 290023
rect 253577 289961 253625 289989
rect 253653 289961 253687 289989
rect 253715 289961 253749 289989
rect 253777 289961 253811 289989
rect 253839 289961 253887 289989
rect 253577 281175 253887 289961
rect 253577 281147 253625 281175
rect 253653 281147 253687 281175
rect 253715 281147 253749 281175
rect 253777 281147 253811 281175
rect 253839 281147 253887 281175
rect 253577 281113 253887 281147
rect 253577 281085 253625 281113
rect 253653 281085 253687 281113
rect 253715 281085 253749 281113
rect 253777 281085 253811 281113
rect 253839 281085 253887 281113
rect 253577 281051 253887 281085
rect 253577 281023 253625 281051
rect 253653 281023 253687 281051
rect 253715 281023 253749 281051
rect 253777 281023 253811 281051
rect 253839 281023 253887 281051
rect 253577 280989 253887 281023
rect 253577 280961 253625 280989
rect 253653 280961 253687 280989
rect 253715 280961 253749 280989
rect 253777 280961 253811 280989
rect 253839 280961 253887 280989
rect 253577 272175 253887 280961
rect 253577 272147 253625 272175
rect 253653 272147 253687 272175
rect 253715 272147 253749 272175
rect 253777 272147 253811 272175
rect 253839 272147 253887 272175
rect 253577 272113 253887 272147
rect 253577 272085 253625 272113
rect 253653 272085 253687 272113
rect 253715 272085 253749 272113
rect 253777 272085 253811 272113
rect 253839 272085 253887 272113
rect 253577 272051 253887 272085
rect 253577 272023 253625 272051
rect 253653 272023 253687 272051
rect 253715 272023 253749 272051
rect 253777 272023 253811 272051
rect 253839 272023 253887 272051
rect 253577 271989 253887 272023
rect 253577 271961 253625 271989
rect 253653 271961 253687 271989
rect 253715 271961 253749 271989
rect 253777 271961 253811 271989
rect 253839 271961 253887 271989
rect 253577 263175 253887 271961
rect 253577 263147 253625 263175
rect 253653 263147 253687 263175
rect 253715 263147 253749 263175
rect 253777 263147 253811 263175
rect 253839 263147 253887 263175
rect 253577 263113 253887 263147
rect 253577 263085 253625 263113
rect 253653 263085 253687 263113
rect 253715 263085 253749 263113
rect 253777 263085 253811 263113
rect 253839 263085 253887 263113
rect 253577 263051 253887 263085
rect 253577 263023 253625 263051
rect 253653 263023 253687 263051
rect 253715 263023 253749 263051
rect 253777 263023 253811 263051
rect 253839 263023 253887 263051
rect 253577 262989 253887 263023
rect 253577 262961 253625 262989
rect 253653 262961 253687 262989
rect 253715 262961 253749 262989
rect 253777 262961 253811 262989
rect 253839 262961 253887 262989
rect 253577 254175 253887 262961
rect 253577 254147 253625 254175
rect 253653 254147 253687 254175
rect 253715 254147 253749 254175
rect 253777 254147 253811 254175
rect 253839 254147 253887 254175
rect 253577 254113 253887 254147
rect 253577 254085 253625 254113
rect 253653 254085 253687 254113
rect 253715 254085 253749 254113
rect 253777 254085 253811 254113
rect 253839 254085 253887 254113
rect 253577 254051 253887 254085
rect 253577 254023 253625 254051
rect 253653 254023 253687 254051
rect 253715 254023 253749 254051
rect 253777 254023 253811 254051
rect 253839 254023 253887 254051
rect 253577 253989 253887 254023
rect 253577 253961 253625 253989
rect 253653 253961 253687 253989
rect 253715 253961 253749 253989
rect 253777 253961 253811 253989
rect 253839 253961 253887 253989
rect 253577 245175 253887 253961
rect 253577 245147 253625 245175
rect 253653 245147 253687 245175
rect 253715 245147 253749 245175
rect 253777 245147 253811 245175
rect 253839 245147 253887 245175
rect 253577 245113 253887 245147
rect 253577 245085 253625 245113
rect 253653 245085 253687 245113
rect 253715 245085 253749 245113
rect 253777 245085 253811 245113
rect 253839 245085 253887 245113
rect 253577 245051 253887 245085
rect 253577 245023 253625 245051
rect 253653 245023 253687 245051
rect 253715 245023 253749 245051
rect 253777 245023 253811 245051
rect 253839 245023 253887 245051
rect 253577 244989 253887 245023
rect 253577 244961 253625 244989
rect 253653 244961 253687 244989
rect 253715 244961 253749 244989
rect 253777 244961 253811 244989
rect 253839 244961 253887 244989
rect 253577 236175 253887 244961
rect 253577 236147 253625 236175
rect 253653 236147 253687 236175
rect 253715 236147 253749 236175
rect 253777 236147 253811 236175
rect 253839 236147 253887 236175
rect 253577 236113 253887 236147
rect 253577 236085 253625 236113
rect 253653 236085 253687 236113
rect 253715 236085 253749 236113
rect 253777 236085 253811 236113
rect 253839 236085 253887 236113
rect 253577 236051 253887 236085
rect 253577 236023 253625 236051
rect 253653 236023 253687 236051
rect 253715 236023 253749 236051
rect 253777 236023 253811 236051
rect 253839 236023 253887 236051
rect 253577 235989 253887 236023
rect 253577 235961 253625 235989
rect 253653 235961 253687 235989
rect 253715 235961 253749 235989
rect 253777 235961 253811 235989
rect 253839 235961 253887 235989
rect 253577 227175 253887 235961
rect 253577 227147 253625 227175
rect 253653 227147 253687 227175
rect 253715 227147 253749 227175
rect 253777 227147 253811 227175
rect 253839 227147 253887 227175
rect 253577 227113 253887 227147
rect 253577 227085 253625 227113
rect 253653 227085 253687 227113
rect 253715 227085 253749 227113
rect 253777 227085 253811 227113
rect 253839 227085 253887 227113
rect 253577 227051 253887 227085
rect 253577 227023 253625 227051
rect 253653 227023 253687 227051
rect 253715 227023 253749 227051
rect 253777 227023 253811 227051
rect 253839 227023 253887 227051
rect 253577 226989 253887 227023
rect 253577 226961 253625 226989
rect 253653 226961 253687 226989
rect 253715 226961 253749 226989
rect 253777 226961 253811 226989
rect 253839 226961 253887 226989
rect 253577 218175 253887 226961
rect 253577 218147 253625 218175
rect 253653 218147 253687 218175
rect 253715 218147 253749 218175
rect 253777 218147 253811 218175
rect 253839 218147 253887 218175
rect 253577 218113 253887 218147
rect 253577 218085 253625 218113
rect 253653 218085 253687 218113
rect 253715 218085 253749 218113
rect 253777 218085 253811 218113
rect 253839 218085 253887 218113
rect 253577 218051 253887 218085
rect 253577 218023 253625 218051
rect 253653 218023 253687 218051
rect 253715 218023 253749 218051
rect 253777 218023 253811 218051
rect 253839 218023 253887 218051
rect 253577 217989 253887 218023
rect 253577 217961 253625 217989
rect 253653 217961 253687 217989
rect 253715 217961 253749 217989
rect 253777 217961 253811 217989
rect 253839 217961 253887 217989
rect 253577 209175 253887 217961
rect 253577 209147 253625 209175
rect 253653 209147 253687 209175
rect 253715 209147 253749 209175
rect 253777 209147 253811 209175
rect 253839 209147 253887 209175
rect 253577 209113 253887 209147
rect 253577 209085 253625 209113
rect 253653 209085 253687 209113
rect 253715 209085 253749 209113
rect 253777 209085 253811 209113
rect 253839 209085 253887 209113
rect 253577 209051 253887 209085
rect 253577 209023 253625 209051
rect 253653 209023 253687 209051
rect 253715 209023 253749 209051
rect 253777 209023 253811 209051
rect 253839 209023 253887 209051
rect 253577 208989 253887 209023
rect 253577 208961 253625 208989
rect 253653 208961 253687 208989
rect 253715 208961 253749 208989
rect 253777 208961 253811 208989
rect 253839 208961 253887 208989
rect 253577 200175 253887 208961
rect 253577 200147 253625 200175
rect 253653 200147 253687 200175
rect 253715 200147 253749 200175
rect 253777 200147 253811 200175
rect 253839 200147 253887 200175
rect 253577 200113 253887 200147
rect 253577 200085 253625 200113
rect 253653 200085 253687 200113
rect 253715 200085 253749 200113
rect 253777 200085 253811 200113
rect 253839 200085 253887 200113
rect 253577 200051 253887 200085
rect 253577 200023 253625 200051
rect 253653 200023 253687 200051
rect 253715 200023 253749 200051
rect 253777 200023 253811 200051
rect 253839 200023 253887 200051
rect 253577 199989 253887 200023
rect 253577 199961 253625 199989
rect 253653 199961 253687 199989
rect 253715 199961 253749 199989
rect 253777 199961 253811 199989
rect 253839 199961 253887 199989
rect 253577 191175 253887 199961
rect 253577 191147 253625 191175
rect 253653 191147 253687 191175
rect 253715 191147 253749 191175
rect 253777 191147 253811 191175
rect 253839 191147 253887 191175
rect 253577 191113 253887 191147
rect 253577 191085 253625 191113
rect 253653 191085 253687 191113
rect 253715 191085 253749 191113
rect 253777 191085 253811 191113
rect 253839 191085 253887 191113
rect 253577 191051 253887 191085
rect 253577 191023 253625 191051
rect 253653 191023 253687 191051
rect 253715 191023 253749 191051
rect 253777 191023 253811 191051
rect 253839 191023 253887 191051
rect 253577 190989 253887 191023
rect 253577 190961 253625 190989
rect 253653 190961 253687 190989
rect 253715 190961 253749 190989
rect 253777 190961 253811 190989
rect 253839 190961 253887 190989
rect 253577 182175 253887 190961
rect 253577 182147 253625 182175
rect 253653 182147 253687 182175
rect 253715 182147 253749 182175
rect 253777 182147 253811 182175
rect 253839 182147 253887 182175
rect 253577 182113 253887 182147
rect 253577 182085 253625 182113
rect 253653 182085 253687 182113
rect 253715 182085 253749 182113
rect 253777 182085 253811 182113
rect 253839 182085 253887 182113
rect 253577 182051 253887 182085
rect 253577 182023 253625 182051
rect 253653 182023 253687 182051
rect 253715 182023 253749 182051
rect 253777 182023 253811 182051
rect 253839 182023 253887 182051
rect 253577 181989 253887 182023
rect 253577 181961 253625 181989
rect 253653 181961 253687 181989
rect 253715 181961 253749 181989
rect 253777 181961 253811 181989
rect 253839 181961 253887 181989
rect 253577 173175 253887 181961
rect 253577 173147 253625 173175
rect 253653 173147 253687 173175
rect 253715 173147 253749 173175
rect 253777 173147 253811 173175
rect 253839 173147 253887 173175
rect 253577 173113 253887 173147
rect 253577 173085 253625 173113
rect 253653 173085 253687 173113
rect 253715 173085 253749 173113
rect 253777 173085 253811 173113
rect 253839 173085 253887 173113
rect 253577 173051 253887 173085
rect 253577 173023 253625 173051
rect 253653 173023 253687 173051
rect 253715 173023 253749 173051
rect 253777 173023 253811 173051
rect 253839 173023 253887 173051
rect 253577 172989 253887 173023
rect 253577 172961 253625 172989
rect 253653 172961 253687 172989
rect 253715 172961 253749 172989
rect 253777 172961 253811 172989
rect 253839 172961 253887 172989
rect 253577 164175 253887 172961
rect 253577 164147 253625 164175
rect 253653 164147 253687 164175
rect 253715 164147 253749 164175
rect 253777 164147 253811 164175
rect 253839 164147 253887 164175
rect 253577 164113 253887 164147
rect 253577 164085 253625 164113
rect 253653 164085 253687 164113
rect 253715 164085 253749 164113
rect 253777 164085 253811 164113
rect 253839 164085 253887 164113
rect 253577 164051 253887 164085
rect 253577 164023 253625 164051
rect 253653 164023 253687 164051
rect 253715 164023 253749 164051
rect 253777 164023 253811 164051
rect 253839 164023 253887 164051
rect 253577 163989 253887 164023
rect 253577 163961 253625 163989
rect 253653 163961 253687 163989
rect 253715 163961 253749 163989
rect 253777 163961 253811 163989
rect 253839 163961 253887 163989
rect 253577 155175 253887 163961
rect 253577 155147 253625 155175
rect 253653 155147 253687 155175
rect 253715 155147 253749 155175
rect 253777 155147 253811 155175
rect 253839 155147 253887 155175
rect 253577 155113 253887 155147
rect 253577 155085 253625 155113
rect 253653 155085 253687 155113
rect 253715 155085 253749 155113
rect 253777 155085 253811 155113
rect 253839 155085 253887 155113
rect 253577 155051 253887 155085
rect 253577 155023 253625 155051
rect 253653 155023 253687 155051
rect 253715 155023 253749 155051
rect 253777 155023 253811 155051
rect 253839 155023 253887 155051
rect 253577 154989 253887 155023
rect 253577 154961 253625 154989
rect 253653 154961 253687 154989
rect 253715 154961 253749 154989
rect 253777 154961 253811 154989
rect 253839 154961 253887 154989
rect 253577 146175 253887 154961
rect 253577 146147 253625 146175
rect 253653 146147 253687 146175
rect 253715 146147 253749 146175
rect 253777 146147 253811 146175
rect 253839 146147 253887 146175
rect 253577 146113 253887 146147
rect 253577 146085 253625 146113
rect 253653 146085 253687 146113
rect 253715 146085 253749 146113
rect 253777 146085 253811 146113
rect 253839 146085 253887 146113
rect 253577 146051 253887 146085
rect 253577 146023 253625 146051
rect 253653 146023 253687 146051
rect 253715 146023 253749 146051
rect 253777 146023 253811 146051
rect 253839 146023 253887 146051
rect 253577 145989 253887 146023
rect 253577 145961 253625 145989
rect 253653 145961 253687 145989
rect 253715 145961 253749 145989
rect 253777 145961 253811 145989
rect 253839 145961 253887 145989
rect 253577 137175 253887 145961
rect 253577 137147 253625 137175
rect 253653 137147 253687 137175
rect 253715 137147 253749 137175
rect 253777 137147 253811 137175
rect 253839 137147 253887 137175
rect 253577 137113 253887 137147
rect 253577 137085 253625 137113
rect 253653 137085 253687 137113
rect 253715 137085 253749 137113
rect 253777 137085 253811 137113
rect 253839 137085 253887 137113
rect 253577 137051 253887 137085
rect 253577 137023 253625 137051
rect 253653 137023 253687 137051
rect 253715 137023 253749 137051
rect 253777 137023 253811 137051
rect 253839 137023 253887 137051
rect 253577 136989 253887 137023
rect 253577 136961 253625 136989
rect 253653 136961 253687 136989
rect 253715 136961 253749 136989
rect 253777 136961 253811 136989
rect 253839 136961 253887 136989
rect 253577 128175 253887 136961
rect 253577 128147 253625 128175
rect 253653 128147 253687 128175
rect 253715 128147 253749 128175
rect 253777 128147 253811 128175
rect 253839 128147 253887 128175
rect 253577 128113 253887 128147
rect 253577 128085 253625 128113
rect 253653 128085 253687 128113
rect 253715 128085 253749 128113
rect 253777 128085 253811 128113
rect 253839 128085 253887 128113
rect 253577 128051 253887 128085
rect 253577 128023 253625 128051
rect 253653 128023 253687 128051
rect 253715 128023 253749 128051
rect 253777 128023 253811 128051
rect 253839 128023 253887 128051
rect 253577 127989 253887 128023
rect 253577 127961 253625 127989
rect 253653 127961 253687 127989
rect 253715 127961 253749 127989
rect 253777 127961 253811 127989
rect 253839 127961 253887 127989
rect 253577 119175 253887 127961
rect 253577 119147 253625 119175
rect 253653 119147 253687 119175
rect 253715 119147 253749 119175
rect 253777 119147 253811 119175
rect 253839 119147 253887 119175
rect 253577 119113 253887 119147
rect 253577 119085 253625 119113
rect 253653 119085 253687 119113
rect 253715 119085 253749 119113
rect 253777 119085 253811 119113
rect 253839 119085 253887 119113
rect 253577 119051 253887 119085
rect 253577 119023 253625 119051
rect 253653 119023 253687 119051
rect 253715 119023 253749 119051
rect 253777 119023 253811 119051
rect 253839 119023 253887 119051
rect 253577 118989 253887 119023
rect 253577 118961 253625 118989
rect 253653 118961 253687 118989
rect 253715 118961 253749 118989
rect 253777 118961 253811 118989
rect 253839 118961 253887 118989
rect 253577 110175 253887 118961
rect 253577 110147 253625 110175
rect 253653 110147 253687 110175
rect 253715 110147 253749 110175
rect 253777 110147 253811 110175
rect 253839 110147 253887 110175
rect 253577 110113 253887 110147
rect 253577 110085 253625 110113
rect 253653 110085 253687 110113
rect 253715 110085 253749 110113
rect 253777 110085 253811 110113
rect 253839 110085 253887 110113
rect 253577 110051 253887 110085
rect 253577 110023 253625 110051
rect 253653 110023 253687 110051
rect 253715 110023 253749 110051
rect 253777 110023 253811 110051
rect 253839 110023 253887 110051
rect 253577 109989 253887 110023
rect 253577 109961 253625 109989
rect 253653 109961 253687 109989
rect 253715 109961 253749 109989
rect 253777 109961 253811 109989
rect 253839 109961 253887 109989
rect 253577 101175 253887 109961
rect 253577 101147 253625 101175
rect 253653 101147 253687 101175
rect 253715 101147 253749 101175
rect 253777 101147 253811 101175
rect 253839 101147 253887 101175
rect 253577 101113 253887 101147
rect 253577 101085 253625 101113
rect 253653 101085 253687 101113
rect 253715 101085 253749 101113
rect 253777 101085 253811 101113
rect 253839 101085 253887 101113
rect 253577 101051 253887 101085
rect 253577 101023 253625 101051
rect 253653 101023 253687 101051
rect 253715 101023 253749 101051
rect 253777 101023 253811 101051
rect 253839 101023 253887 101051
rect 253577 100989 253887 101023
rect 253577 100961 253625 100989
rect 253653 100961 253687 100989
rect 253715 100961 253749 100989
rect 253777 100961 253811 100989
rect 253839 100961 253887 100989
rect 253577 92175 253887 100961
rect 253577 92147 253625 92175
rect 253653 92147 253687 92175
rect 253715 92147 253749 92175
rect 253777 92147 253811 92175
rect 253839 92147 253887 92175
rect 253577 92113 253887 92147
rect 253577 92085 253625 92113
rect 253653 92085 253687 92113
rect 253715 92085 253749 92113
rect 253777 92085 253811 92113
rect 253839 92085 253887 92113
rect 253577 92051 253887 92085
rect 253577 92023 253625 92051
rect 253653 92023 253687 92051
rect 253715 92023 253749 92051
rect 253777 92023 253811 92051
rect 253839 92023 253887 92051
rect 253577 91989 253887 92023
rect 253577 91961 253625 91989
rect 253653 91961 253687 91989
rect 253715 91961 253749 91989
rect 253777 91961 253811 91989
rect 253839 91961 253887 91989
rect 253577 83175 253887 91961
rect 253577 83147 253625 83175
rect 253653 83147 253687 83175
rect 253715 83147 253749 83175
rect 253777 83147 253811 83175
rect 253839 83147 253887 83175
rect 253577 83113 253887 83147
rect 253577 83085 253625 83113
rect 253653 83085 253687 83113
rect 253715 83085 253749 83113
rect 253777 83085 253811 83113
rect 253839 83085 253887 83113
rect 253577 83051 253887 83085
rect 253577 83023 253625 83051
rect 253653 83023 253687 83051
rect 253715 83023 253749 83051
rect 253777 83023 253811 83051
rect 253839 83023 253887 83051
rect 253577 82989 253887 83023
rect 253577 82961 253625 82989
rect 253653 82961 253687 82989
rect 253715 82961 253749 82989
rect 253777 82961 253811 82989
rect 253839 82961 253887 82989
rect 253577 74175 253887 82961
rect 253577 74147 253625 74175
rect 253653 74147 253687 74175
rect 253715 74147 253749 74175
rect 253777 74147 253811 74175
rect 253839 74147 253887 74175
rect 253577 74113 253887 74147
rect 253577 74085 253625 74113
rect 253653 74085 253687 74113
rect 253715 74085 253749 74113
rect 253777 74085 253811 74113
rect 253839 74085 253887 74113
rect 253577 74051 253887 74085
rect 253577 74023 253625 74051
rect 253653 74023 253687 74051
rect 253715 74023 253749 74051
rect 253777 74023 253811 74051
rect 253839 74023 253887 74051
rect 253577 73989 253887 74023
rect 253577 73961 253625 73989
rect 253653 73961 253687 73989
rect 253715 73961 253749 73989
rect 253777 73961 253811 73989
rect 253839 73961 253887 73989
rect 253577 65175 253887 73961
rect 253577 65147 253625 65175
rect 253653 65147 253687 65175
rect 253715 65147 253749 65175
rect 253777 65147 253811 65175
rect 253839 65147 253887 65175
rect 253577 65113 253887 65147
rect 253577 65085 253625 65113
rect 253653 65085 253687 65113
rect 253715 65085 253749 65113
rect 253777 65085 253811 65113
rect 253839 65085 253887 65113
rect 253577 65051 253887 65085
rect 253577 65023 253625 65051
rect 253653 65023 253687 65051
rect 253715 65023 253749 65051
rect 253777 65023 253811 65051
rect 253839 65023 253887 65051
rect 253577 64989 253887 65023
rect 253577 64961 253625 64989
rect 253653 64961 253687 64989
rect 253715 64961 253749 64989
rect 253777 64961 253811 64989
rect 253839 64961 253887 64989
rect 253577 56175 253887 64961
rect 253577 56147 253625 56175
rect 253653 56147 253687 56175
rect 253715 56147 253749 56175
rect 253777 56147 253811 56175
rect 253839 56147 253887 56175
rect 253577 56113 253887 56147
rect 253577 56085 253625 56113
rect 253653 56085 253687 56113
rect 253715 56085 253749 56113
rect 253777 56085 253811 56113
rect 253839 56085 253887 56113
rect 253577 56051 253887 56085
rect 253577 56023 253625 56051
rect 253653 56023 253687 56051
rect 253715 56023 253749 56051
rect 253777 56023 253811 56051
rect 253839 56023 253887 56051
rect 253577 55989 253887 56023
rect 253577 55961 253625 55989
rect 253653 55961 253687 55989
rect 253715 55961 253749 55989
rect 253777 55961 253811 55989
rect 253839 55961 253887 55989
rect 253577 47175 253887 55961
rect 253577 47147 253625 47175
rect 253653 47147 253687 47175
rect 253715 47147 253749 47175
rect 253777 47147 253811 47175
rect 253839 47147 253887 47175
rect 253577 47113 253887 47147
rect 253577 47085 253625 47113
rect 253653 47085 253687 47113
rect 253715 47085 253749 47113
rect 253777 47085 253811 47113
rect 253839 47085 253887 47113
rect 253577 47051 253887 47085
rect 253577 47023 253625 47051
rect 253653 47023 253687 47051
rect 253715 47023 253749 47051
rect 253777 47023 253811 47051
rect 253839 47023 253887 47051
rect 253577 46989 253887 47023
rect 253577 46961 253625 46989
rect 253653 46961 253687 46989
rect 253715 46961 253749 46989
rect 253777 46961 253811 46989
rect 253839 46961 253887 46989
rect 253577 38175 253887 46961
rect 253577 38147 253625 38175
rect 253653 38147 253687 38175
rect 253715 38147 253749 38175
rect 253777 38147 253811 38175
rect 253839 38147 253887 38175
rect 253577 38113 253887 38147
rect 253577 38085 253625 38113
rect 253653 38085 253687 38113
rect 253715 38085 253749 38113
rect 253777 38085 253811 38113
rect 253839 38085 253887 38113
rect 253577 38051 253887 38085
rect 253577 38023 253625 38051
rect 253653 38023 253687 38051
rect 253715 38023 253749 38051
rect 253777 38023 253811 38051
rect 253839 38023 253887 38051
rect 253577 37989 253887 38023
rect 253577 37961 253625 37989
rect 253653 37961 253687 37989
rect 253715 37961 253749 37989
rect 253777 37961 253811 37989
rect 253839 37961 253887 37989
rect 253577 29175 253887 37961
rect 253577 29147 253625 29175
rect 253653 29147 253687 29175
rect 253715 29147 253749 29175
rect 253777 29147 253811 29175
rect 253839 29147 253887 29175
rect 253577 29113 253887 29147
rect 253577 29085 253625 29113
rect 253653 29085 253687 29113
rect 253715 29085 253749 29113
rect 253777 29085 253811 29113
rect 253839 29085 253887 29113
rect 253577 29051 253887 29085
rect 253577 29023 253625 29051
rect 253653 29023 253687 29051
rect 253715 29023 253749 29051
rect 253777 29023 253811 29051
rect 253839 29023 253887 29051
rect 253577 28989 253887 29023
rect 253577 28961 253625 28989
rect 253653 28961 253687 28989
rect 253715 28961 253749 28989
rect 253777 28961 253811 28989
rect 253839 28961 253887 28989
rect 253577 20175 253887 28961
rect 253577 20147 253625 20175
rect 253653 20147 253687 20175
rect 253715 20147 253749 20175
rect 253777 20147 253811 20175
rect 253839 20147 253887 20175
rect 253577 20113 253887 20147
rect 253577 20085 253625 20113
rect 253653 20085 253687 20113
rect 253715 20085 253749 20113
rect 253777 20085 253811 20113
rect 253839 20085 253887 20113
rect 253577 20051 253887 20085
rect 253577 20023 253625 20051
rect 253653 20023 253687 20051
rect 253715 20023 253749 20051
rect 253777 20023 253811 20051
rect 253839 20023 253887 20051
rect 253577 19989 253887 20023
rect 253577 19961 253625 19989
rect 253653 19961 253687 19989
rect 253715 19961 253749 19989
rect 253777 19961 253811 19989
rect 253839 19961 253887 19989
rect 253577 11175 253887 19961
rect 253577 11147 253625 11175
rect 253653 11147 253687 11175
rect 253715 11147 253749 11175
rect 253777 11147 253811 11175
rect 253839 11147 253887 11175
rect 253577 11113 253887 11147
rect 253577 11085 253625 11113
rect 253653 11085 253687 11113
rect 253715 11085 253749 11113
rect 253777 11085 253811 11113
rect 253839 11085 253887 11113
rect 253577 11051 253887 11085
rect 253577 11023 253625 11051
rect 253653 11023 253687 11051
rect 253715 11023 253749 11051
rect 253777 11023 253811 11051
rect 253839 11023 253887 11051
rect 253577 10989 253887 11023
rect 253577 10961 253625 10989
rect 253653 10961 253687 10989
rect 253715 10961 253749 10989
rect 253777 10961 253811 10989
rect 253839 10961 253887 10989
rect 253577 2175 253887 10961
rect 253577 2147 253625 2175
rect 253653 2147 253687 2175
rect 253715 2147 253749 2175
rect 253777 2147 253811 2175
rect 253839 2147 253887 2175
rect 253577 2113 253887 2147
rect 253577 2085 253625 2113
rect 253653 2085 253687 2113
rect 253715 2085 253749 2113
rect 253777 2085 253811 2113
rect 253839 2085 253887 2113
rect 253577 2051 253887 2085
rect 253577 2023 253625 2051
rect 253653 2023 253687 2051
rect 253715 2023 253749 2051
rect 253777 2023 253811 2051
rect 253839 2023 253887 2051
rect 253577 1989 253887 2023
rect 253577 1961 253625 1989
rect 253653 1961 253687 1989
rect 253715 1961 253749 1989
rect 253777 1961 253811 1989
rect 253839 1961 253887 1989
rect 253577 -80 253887 1961
rect 253577 -108 253625 -80
rect 253653 -108 253687 -80
rect 253715 -108 253749 -80
rect 253777 -108 253811 -80
rect 253839 -108 253887 -80
rect 253577 -142 253887 -108
rect 253577 -170 253625 -142
rect 253653 -170 253687 -142
rect 253715 -170 253749 -142
rect 253777 -170 253811 -142
rect 253839 -170 253887 -142
rect 253577 -204 253887 -170
rect 253577 -232 253625 -204
rect 253653 -232 253687 -204
rect 253715 -232 253749 -204
rect 253777 -232 253811 -204
rect 253839 -232 253887 -204
rect 253577 -266 253887 -232
rect 253577 -294 253625 -266
rect 253653 -294 253687 -266
rect 253715 -294 253749 -266
rect 253777 -294 253811 -266
rect 253839 -294 253887 -266
rect 253577 -822 253887 -294
rect 255437 299086 255747 299134
rect 255437 299058 255485 299086
rect 255513 299058 255547 299086
rect 255575 299058 255609 299086
rect 255637 299058 255671 299086
rect 255699 299058 255747 299086
rect 255437 299024 255747 299058
rect 255437 298996 255485 299024
rect 255513 298996 255547 299024
rect 255575 298996 255609 299024
rect 255637 298996 255671 299024
rect 255699 298996 255747 299024
rect 255437 298962 255747 298996
rect 255437 298934 255485 298962
rect 255513 298934 255547 298962
rect 255575 298934 255609 298962
rect 255637 298934 255671 298962
rect 255699 298934 255747 298962
rect 255437 298900 255747 298934
rect 255437 298872 255485 298900
rect 255513 298872 255547 298900
rect 255575 298872 255609 298900
rect 255637 298872 255671 298900
rect 255699 298872 255747 298900
rect 255437 293175 255747 298872
rect 255437 293147 255485 293175
rect 255513 293147 255547 293175
rect 255575 293147 255609 293175
rect 255637 293147 255671 293175
rect 255699 293147 255747 293175
rect 255437 293113 255747 293147
rect 255437 293085 255485 293113
rect 255513 293085 255547 293113
rect 255575 293085 255609 293113
rect 255637 293085 255671 293113
rect 255699 293085 255747 293113
rect 255437 293051 255747 293085
rect 255437 293023 255485 293051
rect 255513 293023 255547 293051
rect 255575 293023 255609 293051
rect 255637 293023 255671 293051
rect 255699 293023 255747 293051
rect 255437 292989 255747 293023
rect 255437 292961 255485 292989
rect 255513 292961 255547 292989
rect 255575 292961 255609 292989
rect 255637 292961 255671 292989
rect 255699 292961 255747 292989
rect 255437 284175 255747 292961
rect 255437 284147 255485 284175
rect 255513 284147 255547 284175
rect 255575 284147 255609 284175
rect 255637 284147 255671 284175
rect 255699 284147 255747 284175
rect 255437 284113 255747 284147
rect 255437 284085 255485 284113
rect 255513 284085 255547 284113
rect 255575 284085 255609 284113
rect 255637 284085 255671 284113
rect 255699 284085 255747 284113
rect 255437 284051 255747 284085
rect 255437 284023 255485 284051
rect 255513 284023 255547 284051
rect 255575 284023 255609 284051
rect 255637 284023 255671 284051
rect 255699 284023 255747 284051
rect 255437 283989 255747 284023
rect 255437 283961 255485 283989
rect 255513 283961 255547 283989
rect 255575 283961 255609 283989
rect 255637 283961 255671 283989
rect 255699 283961 255747 283989
rect 255437 275175 255747 283961
rect 255437 275147 255485 275175
rect 255513 275147 255547 275175
rect 255575 275147 255609 275175
rect 255637 275147 255671 275175
rect 255699 275147 255747 275175
rect 255437 275113 255747 275147
rect 255437 275085 255485 275113
rect 255513 275085 255547 275113
rect 255575 275085 255609 275113
rect 255637 275085 255671 275113
rect 255699 275085 255747 275113
rect 255437 275051 255747 275085
rect 255437 275023 255485 275051
rect 255513 275023 255547 275051
rect 255575 275023 255609 275051
rect 255637 275023 255671 275051
rect 255699 275023 255747 275051
rect 255437 274989 255747 275023
rect 255437 274961 255485 274989
rect 255513 274961 255547 274989
rect 255575 274961 255609 274989
rect 255637 274961 255671 274989
rect 255699 274961 255747 274989
rect 255437 266175 255747 274961
rect 255437 266147 255485 266175
rect 255513 266147 255547 266175
rect 255575 266147 255609 266175
rect 255637 266147 255671 266175
rect 255699 266147 255747 266175
rect 255437 266113 255747 266147
rect 255437 266085 255485 266113
rect 255513 266085 255547 266113
rect 255575 266085 255609 266113
rect 255637 266085 255671 266113
rect 255699 266085 255747 266113
rect 255437 266051 255747 266085
rect 255437 266023 255485 266051
rect 255513 266023 255547 266051
rect 255575 266023 255609 266051
rect 255637 266023 255671 266051
rect 255699 266023 255747 266051
rect 255437 265989 255747 266023
rect 255437 265961 255485 265989
rect 255513 265961 255547 265989
rect 255575 265961 255609 265989
rect 255637 265961 255671 265989
rect 255699 265961 255747 265989
rect 255437 257175 255747 265961
rect 255437 257147 255485 257175
rect 255513 257147 255547 257175
rect 255575 257147 255609 257175
rect 255637 257147 255671 257175
rect 255699 257147 255747 257175
rect 255437 257113 255747 257147
rect 255437 257085 255485 257113
rect 255513 257085 255547 257113
rect 255575 257085 255609 257113
rect 255637 257085 255671 257113
rect 255699 257085 255747 257113
rect 255437 257051 255747 257085
rect 255437 257023 255485 257051
rect 255513 257023 255547 257051
rect 255575 257023 255609 257051
rect 255637 257023 255671 257051
rect 255699 257023 255747 257051
rect 255437 256989 255747 257023
rect 255437 256961 255485 256989
rect 255513 256961 255547 256989
rect 255575 256961 255609 256989
rect 255637 256961 255671 256989
rect 255699 256961 255747 256989
rect 255437 248175 255747 256961
rect 255437 248147 255485 248175
rect 255513 248147 255547 248175
rect 255575 248147 255609 248175
rect 255637 248147 255671 248175
rect 255699 248147 255747 248175
rect 255437 248113 255747 248147
rect 255437 248085 255485 248113
rect 255513 248085 255547 248113
rect 255575 248085 255609 248113
rect 255637 248085 255671 248113
rect 255699 248085 255747 248113
rect 255437 248051 255747 248085
rect 255437 248023 255485 248051
rect 255513 248023 255547 248051
rect 255575 248023 255609 248051
rect 255637 248023 255671 248051
rect 255699 248023 255747 248051
rect 255437 247989 255747 248023
rect 255437 247961 255485 247989
rect 255513 247961 255547 247989
rect 255575 247961 255609 247989
rect 255637 247961 255671 247989
rect 255699 247961 255747 247989
rect 255437 239175 255747 247961
rect 255437 239147 255485 239175
rect 255513 239147 255547 239175
rect 255575 239147 255609 239175
rect 255637 239147 255671 239175
rect 255699 239147 255747 239175
rect 255437 239113 255747 239147
rect 255437 239085 255485 239113
rect 255513 239085 255547 239113
rect 255575 239085 255609 239113
rect 255637 239085 255671 239113
rect 255699 239085 255747 239113
rect 255437 239051 255747 239085
rect 255437 239023 255485 239051
rect 255513 239023 255547 239051
rect 255575 239023 255609 239051
rect 255637 239023 255671 239051
rect 255699 239023 255747 239051
rect 255437 238989 255747 239023
rect 255437 238961 255485 238989
rect 255513 238961 255547 238989
rect 255575 238961 255609 238989
rect 255637 238961 255671 238989
rect 255699 238961 255747 238989
rect 255437 230175 255747 238961
rect 255437 230147 255485 230175
rect 255513 230147 255547 230175
rect 255575 230147 255609 230175
rect 255637 230147 255671 230175
rect 255699 230147 255747 230175
rect 255437 230113 255747 230147
rect 255437 230085 255485 230113
rect 255513 230085 255547 230113
rect 255575 230085 255609 230113
rect 255637 230085 255671 230113
rect 255699 230085 255747 230113
rect 255437 230051 255747 230085
rect 255437 230023 255485 230051
rect 255513 230023 255547 230051
rect 255575 230023 255609 230051
rect 255637 230023 255671 230051
rect 255699 230023 255747 230051
rect 255437 229989 255747 230023
rect 255437 229961 255485 229989
rect 255513 229961 255547 229989
rect 255575 229961 255609 229989
rect 255637 229961 255671 229989
rect 255699 229961 255747 229989
rect 255437 221175 255747 229961
rect 255437 221147 255485 221175
rect 255513 221147 255547 221175
rect 255575 221147 255609 221175
rect 255637 221147 255671 221175
rect 255699 221147 255747 221175
rect 255437 221113 255747 221147
rect 255437 221085 255485 221113
rect 255513 221085 255547 221113
rect 255575 221085 255609 221113
rect 255637 221085 255671 221113
rect 255699 221085 255747 221113
rect 255437 221051 255747 221085
rect 255437 221023 255485 221051
rect 255513 221023 255547 221051
rect 255575 221023 255609 221051
rect 255637 221023 255671 221051
rect 255699 221023 255747 221051
rect 255437 220989 255747 221023
rect 255437 220961 255485 220989
rect 255513 220961 255547 220989
rect 255575 220961 255609 220989
rect 255637 220961 255671 220989
rect 255699 220961 255747 220989
rect 255437 212175 255747 220961
rect 255437 212147 255485 212175
rect 255513 212147 255547 212175
rect 255575 212147 255609 212175
rect 255637 212147 255671 212175
rect 255699 212147 255747 212175
rect 255437 212113 255747 212147
rect 255437 212085 255485 212113
rect 255513 212085 255547 212113
rect 255575 212085 255609 212113
rect 255637 212085 255671 212113
rect 255699 212085 255747 212113
rect 255437 212051 255747 212085
rect 255437 212023 255485 212051
rect 255513 212023 255547 212051
rect 255575 212023 255609 212051
rect 255637 212023 255671 212051
rect 255699 212023 255747 212051
rect 255437 211989 255747 212023
rect 255437 211961 255485 211989
rect 255513 211961 255547 211989
rect 255575 211961 255609 211989
rect 255637 211961 255671 211989
rect 255699 211961 255747 211989
rect 255437 203175 255747 211961
rect 255437 203147 255485 203175
rect 255513 203147 255547 203175
rect 255575 203147 255609 203175
rect 255637 203147 255671 203175
rect 255699 203147 255747 203175
rect 255437 203113 255747 203147
rect 255437 203085 255485 203113
rect 255513 203085 255547 203113
rect 255575 203085 255609 203113
rect 255637 203085 255671 203113
rect 255699 203085 255747 203113
rect 255437 203051 255747 203085
rect 255437 203023 255485 203051
rect 255513 203023 255547 203051
rect 255575 203023 255609 203051
rect 255637 203023 255671 203051
rect 255699 203023 255747 203051
rect 255437 202989 255747 203023
rect 255437 202961 255485 202989
rect 255513 202961 255547 202989
rect 255575 202961 255609 202989
rect 255637 202961 255671 202989
rect 255699 202961 255747 202989
rect 255437 194175 255747 202961
rect 255437 194147 255485 194175
rect 255513 194147 255547 194175
rect 255575 194147 255609 194175
rect 255637 194147 255671 194175
rect 255699 194147 255747 194175
rect 255437 194113 255747 194147
rect 255437 194085 255485 194113
rect 255513 194085 255547 194113
rect 255575 194085 255609 194113
rect 255637 194085 255671 194113
rect 255699 194085 255747 194113
rect 255437 194051 255747 194085
rect 255437 194023 255485 194051
rect 255513 194023 255547 194051
rect 255575 194023 255609 194051
rect 255637 194023 255671 194051
rect 255699 194023 255747 194051
rect 255437 193989 255747 194023
rect 255437 193961 255485 193989
rect 255513 193961 255547 193989
rect 255575 193961 255609 193989
rect 255637 193961 255671 193989
rect 255699 193961 255747 193989
rect 255437 185175 255747 193961
rect 255437 185147 255485 185175
rect 255513 185147 255547 185175
rect 255575 185147 255609 185175
rect 255637 185147 255671 185175
rect 255699 185147 255747 185175
rect 255437 185113 255747 185147
rect 255437 185085 255485 185113
rect 255513 185085 255547 185113
rect 255575 185085 255609 185113
rect 255637 185085 255671 185113
rect 255699 185085 255747 185113
rect 255437 185051 255747 185085
rect 255437 185023 255485 185051
rect 255513 185023 255547 185051
rect 255575 185023 255609 185051
rect 255637 185023 255671 185051
rect 255699 185023 255747 185051
rect 255437 184989 255747 185023
rect 255437 184961 255485 184989
rect 255513 184961 255547 184989
rect 255575 184961 255609 184989
rect 255637 184961 255671 184989
rect 255699 184961 255747 184989
rect 255437 176175 255747 184961
rect 255437 176147 255485 176175
rect 255513 176147 255547 176175
rect 255575 176147 255609 176175
rect 255637 176147 255671 176175
rect 255699 176147 255747 176175
rect 255437 176113 255747 176147
rect 255437 176085 255485 176113
rect 255513 176085 255547 176113
rect 255575 176085 255609 176113
rect 255637 176085 255671 176113
rect 255699 176085 255747 176113
rect 255437 176051 255747 176085
rect 255437 176023 255485 176051
rect 255513 176023 255547 176051
rect 255575 176023 255609 176051
rect 255637 176023 255671 176051
rect 255699 176023 255747 176051
rect 255437 175989 255747 176023
rect 255437 175961 255485 175989
rect 255513 175961 255547 175989
rect 255575 175961 255609 175989
rect 255637 175961 255671 175989
rect 255699 175961 255747 175989
rect 255437 167175 255747 175961
rect 255437 167147 255485 167175
rect 255513 167147 255547 167175
rect 255575 167147 255609 167175
rect 255637 167147 255671 167175
rect 255699 167147 255747 167175
rect 255437 167113 255747 167147
rect 255437 167085 255485 167113
rect 255513 167085 255547 167113
rect 255575 167085 255609 167113
rect 255637 167085 255671 167113
rect 255699 167085 255747 167113
rect 255437 167051 255747 167085
rect 255437 167023 255485 167051
rect 255513 167023 255547 167051
rect 255575 167023 255609 167051
rect 255637 167023 255671 167051
rect 255699 167023 255747 167051
rect 255437 166989 255747 167023
rect 255437 166961 255485 166989
rect 255513 166961 255547 166989
rect 255575 166961 255609 166989
rect 255637 166961 255671 166989
rect 255699 166961 255747 166989
rect 255437 158175 255747 166961
rect 255437 158147 255485 158175
rect 255513 158147 255547 158175
rect 255575 158147 255609 158175
rect 255637 158147 255671 158175
rect 255699 158147 255747 158175
rect 255437 158113 255747 158147
rect 255437 158085 255485 158113
rect 255513 158085 255547 158113
rect 255575 158085 255609 158113
rect 255637 158085 255671 158113
rect 255699 158085 255747 158113
rect 255437 158051 255747 158085
rect 255437 158023 255485 158051
rect 255513 158023 255547 158051
rect 255575 158023 255609 158051
rect 255637 158023 255671 158051
rect 255699 158023 255747 158051
rect 255437 157989 255747 158023
rect 255437 157961 255485 157989
rect 255513 157961 255547 157989
rect 255575 157961 255609 157989
rect 255637 157961 255671 157989
rect 255699 157961 255747 157989
rect 255437 149175 255747 157961
rect 255437 149147 255485 149175
rect 255513 149147 255547 149175
rect 255575 149147 255609 149175
rect 255637 149147 255671 149175
rect 255699 149147 255747 149175
rect 255437 149113 255747 149147
rect 255437 149085 255485 149113
rect 255513 149085 255547 149113
rect 255575 149085 255609 149113
rect 255637 149085 255671 149113
rect 255699 149085 255747 149113
rect 255437 149051 255747 149085
rect 255437 149023 255485 149051
rect 255513 149023 255547 149051
rect 255575 149023 255609 149051
rect 255637 149023 255671 149051
rect 255699 149023 255747 149051
rect 255437 148989 255747 149023
rect 255437 148961 255485 148989
rect 255513 148961 255547 148989
rect 255575 148961 255609 148989
rect 255637 148961 255671 148989
rect 255699 148961 255747 148989
rect 255437 140175 255747 148961
rect 255437 140147 255485 140175
rect 255513 140147 255547 140175
rect 255575 140147 255609 140175
rect 255637 140147 255671 140175
rect 255699 140147 255747 140175
rect 255437 140113 255747 140147
rect 255437 140085 255485 140113
rect 255513 140085 255547 140113
rect 255575 140085 255609 140113
rect 255637 140085 255671 140113
rect 255699 140085 255747 140113
rect 255437 140051 255747 140085
rect 255437 140023 255485 140051
rect 255513 140023 255547 140051
rect 255575 140023 255609 140051
rect 255637 140023 255671 140051
rect 255699 140023 255747 140051
rect 255437 139989 255747 140023
rect 255437 139961 255485 139989
rect 255513 139961 255547 139989
rect 255575 139961 255609 139989
rect 255637 139961 255671 139989
rect 255699 139961 255747 139989
rect 255437 131175 255747 139961
rect 255437 131147 255485 131175
rect 255513 131147 255547 131175
rect 255575 131147 255609 131175
rect 255637 131147 255671 131175
rect 255699 131147 255747 131175
rect 255437 131113 255747 131147
rect 255437 131085 255485 131113
rect 255513 131085 255547 131113
rect 255575 131085 255609 131113
rect 255637 131085 255671 131113
rect 255699 131085 255747 131113
rect 255437 131051 255747 131085
rect 255437 131023 255485 131051
rect 255513 131023 255547 131051
rect 255575 131023 255609 131051
rect 255637 131023 255671 131051
rect 255699 131023 255747 131051
rect 255437 130989 255747 131023
rect 255437 130961 255485 130989
rect 255513 130961 255547 130989
rect 255575 130961 255609 130989
rect 255637 130961 255671 130989
rect 255699 130961 255747 130989
rect 255437 122175 255747 130961
rect 255437 122147 255485 122175
rect 255513 122147 255547 122175
rect 255575 122147 255609 122175
rect 255637 122147 255671 122175
rect 255699 122147 255747 122175
rect 255437 122113 255747 122147
rect 255437 122085 255485 122113
rect 255513 122085 255547 122113
rect 255575 122085 255609 122113
rect 255637 122085 255671 122113
rect 255699 122085 255747 122113
rect 255437 122051 255747 122085
rect 255437 122023 255485 122051
rect 255513 122023 255547 122051
rect 255575 122023 255609 122051
rect 255637 122023 255671 122051
rect 255699 122023 255747 122051
rect 255437 121989 255747 122023
rect 255437 121961 255485 121989
rect 255513 121961 255547 121989
rect 255575 121961 255609 121989
rect 255637 121961 255671 121989
rect 255699 121961 255747 121989
rect 255437 113175 255747 121961
rect 255437 113147 255485 113175
rect 255513 113147 255547 113175
rect 255575 113147 255609 113175
rect 255637 113147 255671 113175
rect 255699 113147 255747 113175
rect 255437 113113 255747 113147
rect 255437 113085 255485 113113
rect 255513 113085 255547 113113
rect 255575 113085 255609 113113
rect 255637 113085 255671 113113
rect 255699 113085 255747 113113
rect 255437 113051 255747 113085
rect 255437 113023 255485 113051
rect 255513 113023 255547 113051
rect 255575 113023 255609 113051
rect 255637 113023 255671 113051
rect 255699 113023 255747 113051
rect 255437 112989 255747 113023
rect 255437 112961 255485 112989
rect 255513 112961 255547 112989
rect 255575 112961 255609 112989
rect 255637 112961 255671 112989
rect 255699 112961 255747 112989
rect 255437 104175 255747 112961
rect 255437 104147 255485 104175
rect 255513 104147 255547 104175
rect 255575 104147 255609 104175
rect 255637 104147 255671 104175
rect 255699 104147 255747 104175
rect 255437 104113 255747 104147
rect 255437 104085 255485 104113
rect 255513 104085 255547 104113
rect 255575 104085 255609 104113
rect 255637 104085 255671 104113
rect 255699 104085 255747 104113
rect 255437 104051 255747 104085
rect 255437 104023 255485 104051
rect 255513 104023 255547 104051
rect 255575 104023 255609 104051
rect 255637 104023 255671 104051
rect 255699 104023 255747 104051
rect 255437 103989 255747 104023
rect 255437 103961 255485 103989
rect 255513 103961 255547 103989
rect 255575 103961 255609 103989
rect 255637 103961 255671 103989
rect 255699 103961 255747 103989
rect 255437 95175 255747 103961
rect 255437 95147 255485 95175
rect 255513 95147 255547 95175
rect 255575 95147 255609 95175
rect 255637 95147 255671 95175
rect 255699 95147 255747 95175
rect 255437 95113 255747 95147
rect 255437 95085 255485 95113
rect 255513 95085 255547 95113
rect 255575 95085 255609 95113
rect 255637 95085 255671 95113
rect 255699 95085 255747 95113
rect 255437 95051 255747 95085
rect 255437 95023 255485 95051
rect 255513 95023 255547 95051
rect 255575 95023 255609 95051
rect 255637 95023 255671 95051
rect 255699 95023 255747 95051
rect 255437 94989 255747 95023
rect 255437 94961 255485 94989
rect 255513 94961 255547 94989
rect 255575 94961 255609 94989
rect 255637 94961 255671 94989
rect 255699 94961 255747 94989
rect 255437 86175 255747 94961
rect 255437 86147 255485 86175
rect 255513 86147 255547 86175
rect 255575 86147 255609 86175
rect 255637 86147 255671 86175
rect 255699 86147 255747 86175
rect 255437 86113 255747 86147
rect 255437 86085 255485 86113
rect 255513 86085 255547 86113
rect 255575 86085 255609 86113
rect 255637 86085 255671 86113
rect 255699 86085 255747 86113
rect 255437 86051 255747 86085
rect 255437 86023 255485 86051
rect 255513 86023 255547 86051
rect 255575 86023 255609 86051
rect 255637 86023 255671 86051
rect 255699 86023 255747 86051
rect 255437 85989 255747 86023
rect 255437 85961 255485 85989
rect 255513 85961 255547 85989
rect 255575 85961 255609 85989
rect 255637 85961 255671 85989
rect 255699 85961 255747 85989
rect 255437 77175 255747 85961
rect 255437 77147 255485 77175
rect 255513 77147 255547 77175
rect 255575 77147 255609 77175
rect 255637 77147 255671 77175
rect 255699 77147 255747 77175
rect 255437 77113 255747 77147
rect 255437 77085 255485 77113
rect 255513 77085 255547 77113
rect 255575 77085 255609 77113
rect 255637 77085 255671 77113
rect 255699 77085 255747 77113
rect 255437 77051 255747 77085
rect 255437 77023 255485 77051
rect 255513 77023 255547 77051
rect 255575 77023 255609 77051
rect 255637 77023 255671 77051
rect 255699 77023 255747 77051
rect 255437 76989 255747 77023
rect 255437 76961 255485 76989
rect 255513 76961 255547 76989
rect 255575 76961 255609 76989
rect 255637 76961 255671 76989
rect 255699 76961 255747 76989
rect 255437 68175 255747 76961
rect 255437 68147 255485 68175
rect 255513 68147 255547 68175
rect 255575 68147 255609 68175
rect 255637 68147 255671 68175
rect 255699 68147 255747 68175
rect 255437 68113 255747 68147
rect 255437 68085 255485 68113
rect 255513 68085 255547 68113
rect 255575 68085 255609 68113
rect 255637 68085 255671 68113
rect 255699 68085 255747 68113
rect 255437 68051 255747 68085
rect 255437 68023 255485 68051
rect 255513 68023 255547 68051
rect 255575 68023 255609 68051
rect 255637 68023 255671 68051
rect 255699 68023 255747 68051
rect 255437 67989 255747 68023
rect 255437 67961 255485 67989
rect 255513 67961 255547 67989
rect 255575 67961 255609 67989
rect 255637 67961 255671 67989
rect 255699 67961 255747 67989
rect 255437 59175 255747 67961
rect 255437 59147 255485 59175
rect 255513 59147 255547 59175
rect 255575 59147 255609 59175
rect 255637 59147 255671 59175
rect 255699 59147 255747 59175
rect 255437 59113 255747 59147
rect 255437 59085 255485 59113
rect 255513 59085 255547 59113
rect 255575 59085 255609 59113
rect 255637 59085 255671 59113
rect 255699 59085 255747 59113
rect 255437 59051 255747 59085
rect 255437 59023 255485 59051
rect 255513 59023 255547 59051
rect 255575 59023 255609 59051
rect 255637 59023 255671 59051
rect 255699 59023 255747 59051
rect 255437 58989 255747 59023
rect 255437 58961 255485 58989
rect 255513 58961 255547 58989
rect 255575 58961 255609 58989
rect 255637 58961 255671 58989
rect 255699 58961 255747 58989
rect 255437 50175 255747 58961
rect 255437 50147 255485 50175
rect 255513 50147 255547 50175
rect 255575 50147 255609 50175
rect 255637 50147 255671 50175
rect 255699 50147 255747 50175
rect 255437 50113 255747 50147
rect 255437 50085 255485 50113
rect 255513 50085 255547 50113
rect 255575 50085 255609 50113
rect 255637 50085 255671 50113
rect 255699 50085 255747 50113
rect 255437 50051 255747 50085
rect 255437 50023 255485 50051
rect 255513 50023 255547 50051
rect 255575 50023 255609 50051
rect 255637 50023 255671 50051
rect 255699 50023 255747 50051
rect 255437 49989 255747 50023
rect 255437 49961 255485 49989
rect 255513 49961 255547 49989
rect 255575 49961 255609 49989
rect 255637 49961 255671 49989
rect 255699 49961 255747 49989
rect 255437 41175 255747 49961
rect 255437 41147 255485 41175
rect 255513 41147 255547 41175
rect 255575 41147 255609 41175
rect 255637 41147 255671 41175
rect 255699 41147 255747 41175
rect 255437 41113 255747 41147
rect 255437 41085 255485 41113
rect 255513 41085 255547 41113
rect 255575 41085 255609 41113
rect 255637 41085 255671 41113
rect 255699 41085 255747 41113
rect 255437 41051 255747 41085
rect 255437 41023 255485 41051
rect 255513 41023 255547 41051
rect 255575 41023 255609 41051
rect 255637 41023 255671 41051
rect 255699 41023 255747 41051
rect 255437 40989 255747 41023
rect 255437 40961 255485 40989
rect 255513 40961 255547 40989
rect 255575 40961 255609 40989
rect 255637 40961 255671 40989
rect 255699 40961 255747 40989
rect 255437 32175 255747 40961
rect 255437 32147 255485 32175
rect 255513 32147 255547 32175
rect 255575 32147 255609 32175
rect 255637 32147 255671 32175
rect 255699 32147 255747 32175
rect 255437 32113 255747 32147
rect 255437 32085 255485 32113
rect 255513 32085 255547 32113
rect 255575 32085 255609 32113
rect 255637 32085 255671 32113
rect 255699 32085 255747 32113
rect 255437 32051 255747 32085
rect 255437 32023 255485 32051
rect 255513 32023 255547 32051
rect 255575 32023 255609 32051
rect 255637 32023 255671 32051
rect 255699 32023 255747 32051
rect 255437 31989 255747 32023
rect 255437 31961 255485 31989
rect 255513 31961 255547 31989
rect 255575 31961 255609 31989
rect 255637 31961 255671 31989
rect 255699 31961 255747 31989
rect 255437 23175 255747 31961
rect 255437 23147 255485 23175
rect 255513 23147 255547 23175
rect 255575 23147 255609 23175
rect 255637 23147 255671 23175
rect 255699 23147 255747 23175
rect 255437 23113 255747 23147
rect 255437 23085 255485 23113
rect 255513 23085 255547 23113
rect 255575 23085 255609 23113
rect 255637 23085 255671 23113
rect 255699 23085 255747 23113
rect 255437 23051 255747 23085
rect 255437 23023 255485 23051
rect 255513 23023 255547 23051
rect 255575 23023 255609 23051
rect 255637 23023 255671 23051
rect 255699 23023 255747 23051
rect 255437 22989 255747 23023
rect 255437 22961 255485 22989
rect 255513 22961 255547 22989
rect 255575 22961 255609 22989
rect 255637 22961 255671 22989
rect 255699 22961 255747 22989
rect 255437 14175 255747 22961
rect 255437 14147 255485 14175
rect 255513 14147 255547 14175
rect 255575 14147 255609 14175
rect 255637 14147 255671 14175
rect 255699 14147 255747 14175
rect 255437 14113 255747 14147
rect 255437 14085 255485 14113
rect 255513 14085 255547 14113
rect 255575 14085 255609 14113
rect 255637 14085 255671 14113
rect 255699 14085 255747 14113
rect 255437 14051 255747 14085
rect 255437 14023 255485 14051
rect 255513 14023 255547 14051
rect 255575 14023 255609 14051
rect 255637 14023 255671 14051
rect 255699 14023 255747 14051
rect 255437 13989 255747 14023
rect 255437 13961 255485 13989
rect 255513 13961 255547 13989
rect 255575 13961 255609 13989
rect 255637 13961 255671 13989
rect 255699 13961 255747 13989
rect 255437 5175 255747 13961
rect 255437 5147 255485 5175
rect 255513 5147 255547 5175
rect 255575 5147 255609 5175
rect 255637 5147 255671 5175
rect 255699 5147 255747 5175
rect 255437 5113 255747 5147
rect 255437 5085 255485 5113
rect 255513 5085 255547 5113
rect 255575 5085 255609 5113
rect 255637 5085 255671 5113
rect 255699 5085 255747 5113
rect 255437 5051 255747 5085
rect 255437 5023 255485 5051
rect 255513 5023 255547 5051
rect 255575 5023 255609 5051
rect 255637 5023 255671 5051
rect 255699 5023 255747 5051
rect 255437 4989 255747 5023
rect 255437 4961 255485 4989
rect 255513 4961 255547 4989
rect 255575 4961 255609 4989
rect 255637 4961 255671 4989
rect 255699 4961 255747 4989
rect 255437 -560 255747 4961
rect 255437 -588 255485 -560
rect 255513 -588 255547 -560
rect 255575 -588 255609 -560
rect 255637 -588 255671 -560
rect 255699 -588 255747 -560
rect 255437 -622 255747 -588
rect 255437 -650 255485 -622
rect 255513 -650 255547 -622
rect 255575 -650 255609 -622
rect 255637 -650 255671 -622
rect 255699 -650 255747 -622
rect 255437 -684 255747 -650
rect 255437 -712 255485 -684
rect 255513 -712 255547 -684
rect 255575 -712 255609 -684
rect 255637 -712 255671 -684
rect 255699 -712 255747 -684
rect 255437 -746 255747 -712
rect 255437 -774 255485 -746
rect 255513 -774 255547 -746
rect 255575 -774 255609 -746
rect 255637 -774 255671 -746
rect 255699 -774 255747 -746
rect 255437 -822 255747 -774
rect 262577 298606 262887 299134
rect 262577 298578 262625 298606
rect 262653 298578 262687 298606
rect 262715 298578 262749 298606
rect 262777 298578 262811 298606
rect 262839 298578 262887 298606
rect 262577 298544 262887 298578
rect 262577 298516 262625 298544
rect 262653 298516 262687 298544
rect 262715 298516 262749 298544
rect 262777 298516 262811 298544
rect 262839 298516 262887 298544
rect 262577 298482 262887 298516
rect 262577 298454 262625 298482
rect 262653 298454 262687 298482
rect 262715 298454 262749 298482
rect 262777 298454 262811 298482
rect 262839 298454 262887 298482
rect 262577 298420 262887 298454
rect 262577 298392 262625 298420
rect 262653 298392 262687 298420
rect 262715 298392 262749 298420
rect 262777 298392 262811 298420
rect 262839 298392 262887 298420
rect 262577 290175 262887 298392
rect 262577 290147 262625 290175
rect 262653 290147 262687 290175
rect 262715 290147 262749 290175
rect 262777 290147 262811 290175
rect 262839 290147 262887 290175
rect 262577 290113 262887 290147
rect 262577 290085 262625 290113
rect 262653 290085 262687 290113
rect 262715 290085 262749 290113
rect 262777 290085 262811 290113
rect 262839 290085 262887 290113
rect 262577 290051 262887 290085
rect 262577 290023 262625 290051
rect 262653 290023 262687 290051
rect 262715 290023 262749 290051
rect 262777 290023 262811 290051
rect 262839 290023 262887 290051
rect 262577 289989 262887 290023
rect 262577 289961 262625 289989
rect 262653 289961 262687 289989
rect 262715 289961 262749 289989
rect 262777 289961 262811 289989
rect 262839 289961 262887 289989
rect 262577 281175 262887 289961
rect 262577 281147 262625 281175
rect 262653 281147 262687 281175
rect 262715 281147 262749 281175
rect 262777 281147 262811 281175
rect 262839 281147 262887 281175
rect 262577 281113 262887 281147
rect 262577 281085 262625 281113
rect 262653 281085 262687 281113
rect 262715 281085 262749 281113
rect 262777 281085 262811 281113
rect 262839 281085 262887 281113
rect 262577 281051 262887 281085
rect 262577 281023 262625 281051
rect 262653 281023 262687 281051
rect 262715 281023 262749 281051
rect 262777 281023 262811 281051
rect 262839 281023 262887 281051
rect 262577 280989 262887 281023
rect 262577 280961 262625 280989
rect 262653 280961 262687 280989
rect 262715 280961 262749 280989
rect 262777 280961 262811 280989
rect 262839 280961 262887 280989
rect 262577 272175 262887 280961
rect 262577 272147 262625 272175
rect 262653 272147 262687 272175
rect 262715 272147 262749 272175
rect 262777 272147 262811 272175
rect 262839 272147 262887 272175
rect 262577 272113 262887 272147
rect 262577 272085 262625 272113
rect 262653 272085 262687 272113
rect 262715 272085 262749 272113
rect 262777 272085 262811 272113
rect 262839 272085 262887 272113
rect 262577 272051 262887 272085
rect 262577 272023 262625 272051
rect 262653 272023 262687 272051
rect 262715 272023 262749 272051
rect 262777 272023 262811 272051
rect 262839 272023 262887 272051
rect 262577 271989 262887 272023
rect 262577 271961 262625 271989
rect 262653 271961 262687 271989
rect 262715 271961 262749 271989
rect 262777 271961 262811 271989
rect 262839 271961 262887 271989
rect 262577 263175 262887 271961
rect 262577 263147 262625 263175
rect 262653 263147 262687 263175
rect 262715 263147 262749 263175
rect 262777 263147 262811 263175
rect 262839 263147 262887 263175
rect 262577 263113 262887 263147
rect 262577 263085 262625 263113
rect 262653 263085 262687 263113
rect 262715 263085 262749 263113
rect 262777 263085 262811 263113
rect 262839 263085 262887 263113
rect 262577 263051 262887 263085
rect 262577 263023 262625 263051
rect 262653 263023 262687 263051
rect 262715 263023 262749 263051
rect 262777 263023 262811 263051
rect 262839 263023 262887 263051
rect 262577 262989 262887 263023
rect 262577 262961 262625 262989
rect 262653 262961 262687 262989
rect 262715 262961 262749 262989
rect 262777 262961 262811 262989
rect 262839 262961 262887 262989
rect 262577 254175 262887 262961
rect 262577 254147 262625 254175
rect 262653 254147 262687 254175
rect 262715 254147 262749 254175
rect 262777 254147 262811 254175
rect 262839 254147 262887 254175
rect 262577 254113 262887 254147
rect 262577 254085 262625 254113
rect 262653 254085 262687 254113
rect 262715 254085 262749 254113
rect 262777 254085 262811 254113
rect 262839 254085 262887 254113
rect 262577 254051 262887 254085
rect 262577 254023 262625 254051
rect 262653 254023 262687 254051
rect 262715 254023 262749 254051
rect 262777 254023 262811 254051
rect 262839 254023 262887 254051
rect 262577 253989 262887 254023
rect 262577 253961 262625 253989
rect 262653 253961 262687 253989
rect 262715 253961 262749 253989
rect 262777 253961 262811 253989
rect 262839 253961 262887 253989
rect 262577 245175 262887 253961
rect 262577 245147 262625 245175
rect 262653 245147 262687 245175
rect 262715 245147 262749 245175
rect 262777 245147 262811 245175
rect 262839 245147 262887 245175
rect 262577 245113 262887 245147
rect 262577 245085 262625 245113
rect 262653 245085 262687 245113
rect 262715 245085 262749 245113
rect 262777 245085 262811 245113
rect 262839 245085 262887 245113
rect 262577 245051 262887 245085
rect 262577 245023 262625 245051
rect 262653 245023 262687 245051
rect 262715 245023 262749 245051
rect 262777 245023 262811 245051
rect 262839 245023 262887 245051
rect 262577 244989 262887 245023
rect 262577 244961 262625 244989
rect 262653 244961 262687 244989
rect 262715 244961 262749 244989
rect 262777 244961 262811 244989
rect 262839 244961 262887 244989
rect 262577 236175 262887 244961
rect 262577 236147 262625 236175
rect 262653 236147 262687 236175
rect 262715 236147 262749 236175
rect 262777 236147 262811 236175
rect 262839 236147 262887 236175
rect 262577 236113 262887 236147
rect 262577 236085 262625 236113
rect 262653 236085 262687 236113
rect 262715 236085 262749 236113
rect 262777 236085 262811 236113
rect 262839 236085 262887 236113
rect 262577 236051 262887 236085
rect 262577 236023 262625 236051
rect 262653 236023 262687 236051
rect 262715 236023 262749 236051
rect 262777 236023 262811 236051
rect 262839 236023 262887 236051
rect 262577 235989 262887 236023
rect 262577 235961 262625 235989
rect 262653 235961 262687 235989
rect 262715 235961 262749 235989
rect 262777 235961 262811 235989
rect 262839 235961 262887 235989
rect 262577 227175 262887 235961
rect 262577 227147 262625 227175
rect 262653 227147 262687 227175
rect 262715 227147 262749 227175
rect 262777 227147 262811 227175
rect 262839 227147 262887 227175
rect 262577 227113 262887 227147
rect 262577 227085 262625 227113
rect 262653 227085 262687 227113
rect 262715 227085 262749 227113
rect 262777 227085 262811 227113
rect 262839 227085 262887 227113
rect 262577 227051 262887 227085
rect 262577 227023 262625 227051
rect 262653 227023 262687 227051
rect 262715 227023 262749 227051
rect 262777 227023 262811 227051
rect 262839 227023 262887 227051
rect 262577 226989 262887 227023
rect 262577 226961 262625 226989
rect 262653 226961 262687 226989
rect 262715 226961 262749 226989
rect 262777 226961 262811 226989
rect 262839 226961 262887 226989
rect 262577 218175 262887 226961
rect 262577 218147 262625 218175
rect 262653 218147 262687 218175
rect 262715 218147 262749 218175
rect 262777 218147 262811 218175
rect 262839 218147 262887 218175
rect 262577 218113 262887 218147
rect 262577 218085 262625 218113
rect 262653 218085 262687 218113
rect 262715 218085 262749 218113
rect 262777 218085 262811 218113
rect 262839 218085 262887 218113
rect 262577 218051 262887 218085
rect 262577 218023 262625 218051
rect 262653 218023 262687 218051
rect 262715 218023 262749 218051
rect 262777 218023 262811 218051
rect 262839 218023 262887 218051
rect 262577 217989 262887 218023
rect 262577 217961 262625 217989
rect 262653 217961 262687 217989
rect 262715 217961 262749 217989
rect 262777 217961 262811 217989
rect 262839 217961 262887 217989
rect 262577 209175 262887 217961
rect 262577 209147 262625 209175
rect 262653 209147 262687 209175
rect 262715 209147 262749 209175
rect 262777 209147 262811 209175
rect 262839 209147 262887 209175
rect 262577 209113 262887 209147
rect 262577 209085 262625 209113
rect 262653 209085 262687 209113
rect 262715 209085 262749 209113
rect 262777 209085 262811 209113
rect 262839 209085 262887 209113
rect 262577 209051 262887 209085
rect 262577 209023 262625 209051
rect 262653 209023 262687 209051
rect 262715 209023 262749 209051
rect 262777 209023 262811 209051
rect 262839 209023 262887 209051
rect 262577 208989 262887 209023
rect 262577 208961 262625 208989
rect 262653 208961 262687 208989
rect 262715 208961 262749 208989
rect 262777 208961 262811 208989
rect 262839 208961 262887 208989
rect 262577 200175 262887 208961
rect 262577 200147 262625 200175
rect 262653 200147 262687 200175
rect 262715 200147 262749 200175
rect 262777 200147 262811 200175
rect 262839 200147 262887 200175
rect 262577 200113 262887 200147
rect 262577 200085 262625 200113
rect 262653 200085 262687 200113
rect 262715 200085 262749 200113
rect 262777 200085 262811 200113
rect 262839 200085 262887 200113
rect 262577 200051 262887 200085
rect 262577 200023 262625 200051
rect 262653 200023 262687 200051
rect 262715 200023 262749 200051
rect 262777 200023 262811 200051
rect 262839 200023 262887 200051
rect 262577 199989 262887 200023
rect 262577 199961 262625 199989
rect 262653 199961 262687 199989
rect 262715 199961 262749 199989
rect 262777 199961 262811 199989
rect 262839 199961 262887 199989
rect 262577 191175 262887 199961
rect 262577 191147 262625 191175
rect 262653 191147 262687 191175
rect 262715 191147 262749 191175
rect 262777 191147 262811 191175
rect 262839 191147 262887 191175
rect 262577 191113 262887 191147
rect 262577 191085 262625 191113
rect 262653 191085 262687 191113
rect 262715 191085 262749 191113
rect 262777 191085 262811 191113
rect 262839 191085 262887 191113
rect 262577 191051 262887 191085
rect 262577 191023 262625 191051
rect 262653 191023 262687 191051
rect 262715 191023 262749 191051
rect 262777 191023 262811 191051
rect 262839 191023 262887 191051
rect 262577 190989 262887 191023
rect 262577 190961 262625 190989
rect 262653 190961 262687 190989
rect 262715 190961 262749 190989
rect 262777 190961 262811 190989
rect 262839 190961 262887 190989
rect 262577 182175 262887 190961
rect 262577 182147 262625 182175
rect 262653 182147 262687 182175
rect 262715 182147 262749 182175
rect 262777 182147 262811 182175
rect 262839 182147 262887 182175
rect 262577 182113 262887 182147
rect 262577 182085 262625 182113
rect 262653 182085 262687 182113
rect 262715 182085 262749 182113
rect 262777 182085 262811 182113
rect 262839 182085 262887 182113
rect 262577 182051 262887 182085
rect 262577 182023 262625 182051
rect 262653 182023 262687 182051
rect 262715 182023 262749 182051
rect 262777 182023 262811 182051
rect 262839 182023 262887 182051
rect 262577 181989 262887 182023
rect 262577 181961 262625 181989
rect 262653 181961 262687 181989
rect 262715 181961 262749 181989
rect 262777 181961 262811 181989
rect 262839 181961 262887 181989
rect 262577 173175 262887 181961
rect 262577 173147 262625 173175
rect 262653 173147 262687 173175
rect 262715 173147 262749 173175
rect 262777 173147 262811 173175
rect 262839 173147 262887 173175
rect 262577 173113 262887 173147
rect 262577 173085 262625 173113
rect 262653 173085 262687 173113
rect 262715 173085 262749 173113
rect 262777 173085 262811 173113
rect 262839 173085 262887 173113
rect 262577 173051 262887 173085
rect 262577 173023 262625 173051
rect 262653 173023 262687 173051
rect 262715 173023 262749 173051
rect 262777 173023 262811 173051
rect 262839 173023 262887 173051
rect 262577 172989 262887 173023
rect 262577 172961 262625 172989
rect 262653 172961 262687 172989
rect 262715 172961 262749 172989
rect 262777 172961 262811 172989
rect 262839 172961 262887 172989
rect 262577 164175 262887 172961
rect 262577 164147 262625 164175
rect 262653 164147 262687 164175
rect 262715 164147 262749 164175
rect 262777 164147 262811 164175
rect 262839 164147 262887 164175
rect 262577 164113 262887 164147
rect 262577 164085 262625 164113
rect 262653 164085 262687 164113
rect 262715 164085 262749 164113
rect 262777 164085 262811 164113
rect 262839 164085 262887 164113
rect 262577 164051 262887 164085
rect 262577 164023 262625 164051
rect 262653 164023 262687 164051
rect 262715 164023 262749 164051
rect 262777 164023 262811 164051
rect 262839 164023 262887 164051
rect 262577 163989 262887 164023
rect 262577 163961 262625 163989
rect 262653 163961 262687 163989
rect 262715 163961 262749 163989
rect 262777 163961 262811 163989
rect 262839 163961 262887 163989
rect 262577 155175 262887 163961
rect 262577 155147 262625 155175
rect 262653 155147 262687 155175
rect 262715 155147 262749 155175
rect 262777 155147 262811 155175
rect 262839 155147 262887 155175
rect 262577 155113 262887 155147
rect 262577 155085 262625 155113
rect 262653 155085 262687 155113
rect 262715 155085 262749 155113
rect 262777 155085 262811 155113
rect 262839 155085 262887 155113
rect 262577 155051 262887 155085
rect 262577 155023 262625 155051
rect 262653 155023 262687 155051
rect 262715 155023 262749 155051
rect 262777 155023 262811 155051
rect 262839 155023 262887 155051
rect 262577 154989 262887 155023
rect 262577 154961 262625 154989
rect 262653 154961 262687 154989
rect 262715 154961 262749 154989
rect 262777 154961 262811 154989
rect 262839 154961 262887 154989
rect 262577 146175 262887 154961
rect 262577 146147 262625 146175
rect 262653 146147 262687 146175
rect 262715 146147 262749 146175
rect 262777 146147 262811 146175
rect 262839 146147 262887 146175
rect 262577 146113 262887 146147
rect 262577 146085 262625 146113
rect 262653 146085 262687 146113
rect 262715 146085 262749 146113
rect 262777 146085 262811 146113
rect 262839 146085 262887 146113
rect 262577 146051 262887 146085
rect 262577 146023 262625 146051
rect 262653 146023 262687 146051
rect 262715 146023 262749 146051
rect 262777 146023 262811 146051
rect 262839 146023 262887 146051
rect 262577 145989 262887 146023
rect 262577 145961 262625 145989
rect 262653 145961 262687 145989
rect 262715 145961 262749 145989
rect 262777 145961 262811 145989
rect 262839 145961 262887 145989
rect 262577 137175 262887 145961
rect 262577 137147 262625 137175
rect 262653 137147 262687 137175
rect 262715 137147 262749 137175
rect 262777 137147 262811 137175
rect 262839 137147 262887 137175
rect 262577 137113 262887 137147
rect 262577 137085 262625 137113
rect 262653 137085 262687 137113
rect 262715 137085 262749 137113
rect 262777 137085 262811 137113
rect 262839 137085 262887 137113
rect 262577 137051 262887 137085
rect 262577 137023 262625 137051
rect 262653 137023 262687 137051
rect 262715 137023 262749 137051
rect 262777 137023 262811 137051
rect 262839 137023 262887 137051
rect 262577 136989 262887 137023
rect 262577 136961 262625 136989
rect 262653 136961 262687 136989
rect 262715 136961 262749 136989
rect 262777 136961 262811 136989
rect 262839 136961 262887 136989
rect 262577 128175 262887 136961
rect 262577 128147 262625 128175
rect 262653 128147 262687 128175
rect 262715 128147 262749 128175
rect 262777 128147 262811 128175
rect 262839 128147 262887 128175
rect 262577 128113 262887 128147
rect 262577 128085 262625 128113
rect 262653 128085 262687 128113
rect 262715 128085 262749 128113
rect 262777 128085 262811 128113
rect 262839 128085 262887 128113
rect 262577 128051 262887 128085
rect 262577 128023 262625 128051
rect 262653 128023 262687 128051
rect 262715 128023 262749 128051
rect 262777 128023 262811 128051
rect 262839 128023 262887 128051
rect 262577 127989 262887 128023
rect 262577 127961 262625 127989
rect 262653 127961 262687 127989
rect 262715 127961 262749 127989
rect 262777 127961 262811 127989
rect 262839 127961 262887 127989
rect 262577 119175 262887 127961
rect 262577 119147 262625 119175
rect 262653 119147 262687 119175
rect 262715 119147 262749 119175
rect 262777 119147 262811 119175
rect 262839 119147 262887 119175
rect 262577 119113 262887 119147
rect 262577 119085 262625 119113
rect 262653 119085 262687 119113
rect 262715 119085 262749 119113
rect 262777 119085 262811 119113
rect 262839 119085 262887 119113
rect 262577 119051 262887 119085
rect 262577 119023 262625 119051
rect 262653 119023 262687 119051
rect 262715 119023 262749 119051
rect 262777 119023 262811 119051
rect 262839 119023 262887 119051
rect 262577 118989 262887 119023
rect 262577 118961 262625 118989
rect 262653 118961 262687 118989
rect 262715 118961 262749 118989
rect 262777 118961 262811 118989
rect 262839 118961 262887 118989
rect 262577 110175 262887 118961
rect 262577 110147 262625 110175
rect 262653 110147 262687 110175
rect 262715 110147 262749 110175
rect 262777 110147 262811 110175
rect 262839 110147 262887 110175
rect 262577 110113 262887 110147
rect 262577 110085 262625 110113
rect 262653 110085 262687 110113
rect 262715 110085 262749 110113
rect 262777 110085 262811 110113
rect 262839 110085 262887 110113
rect 262577 110051 262887 110085
rect 262577 110023 262625 110051
rect 262653 110023 262687 110051
rect 262715 110023 262749 110051
rect 262777 110023 262811 110051
rect 262839 110023 262887 110051
rect 262577 109989 262887 110023
rect 262577 109961 262625 109989
rect 262653 109961 262687 109989
rect 262715 109961 262749 109989
rect 262777 109961 262811 109989
rect 262839 109961 262887 109989
rect 262577 101175 262887 109961
rect 262577 101147 262625 101175
rect 262653 101147 262687 101175
rect 262715 101147 262749 101175
rect 262777 101147 262811 101175
rect 262839 101147 262887 101175
rect 262577 101113 262887 101147
rect 262577 101085 262625 101113
rect 262653 101085 262687 101113
rect 262715 101085 262749 101113
rect 262777 101085 262811 101113
rect 262839 101085 262887 101113
rect 262577 101051 262887 101085
rect 262577 101023 262625 101051
rect 262653 101023 262687 101051
rect 262715 101023 262749 101051
rect 262777 101023 262811 101051
rect 262839 101023 262887 101051
rect 262577 100989 262887 101023
rect 262577 100961 262625 100989
rect 262653 100961 262687 100989
rect 262715 100961 262749 100989
rect 262777 100961 262811 100989
rect 262839 100961 262887 100989
rect 262577 92175 262887 100961
rect 262577 92147 262625 92175
rect 262653 92147 262687 92175
rect 262715 92147 262749 92175
rect 262777 92147 262811 92175
rect 262839 92147 262887 92175
rect 262577 92113 262887 92147
rect 262577 92085 262625 92113
rect 262653 92085 262687 92113
rect 262715 92085 262749 92113
rect 262777 92085 262811 92113
rect 262839 92085 262887 92113
rect 262577 92051 262887 92085
rect 262577 92023 262625 92051
rect 262653 92023 262687 92051
rect 262715 92023 262749 92051
rect 262777 92023 262811 92051
rect 262839 92023 262887 92051
rect 262577 91989 262887 92023
rect 262577 91961 262625 91989
rect 262653 91961 262687 91989
rect 262715 91961 262749 91989
rect 262777 91961 262811 91989
rect 262839 91961 262887 91989
rect 262577 83175 262887 91961
rect 262577 83147 262625 83175
rect 262653 83147 262687 83175
rect 262715 83147 262749 83175
rect 262777 83147 262811 83175
rect 262839 83147 262887 83175
rect 262577 83113 262887 83147
rect 262577 83085 262625 83113
rect 262653 83085 262687 83113
rect 262715 83085 262749 83113
rect 262777 83085 262811 83113
rect 262839 83085 262887 83113
rect 262577 83051 262887 83085
rect 262577 83023 262625 83051
rect 262653 83023 262687 83051
rect 262715 83023 262749 83051
rect 262777 83023 262811 83051
rect 262839 83023 262887 83051
rect 262577 82989 262887 83023
rect 262577 82961 262625 82989
rect 262653 82961 262687 82989
rect 262715 82961 262749 82989
rect 262777 82961 262811 82989
rect 262839 82961 262887 82989
rect 262577 74175 262887 82961
rect 262577 74147 262625 74175
rect 262653 74147 262687 74175
rect 262715 74147 262749 74175
rect 262777 74147 262811 74175
rect 262839 74147 262887 74175
rect 262577 74113 262887 74147
rect 262577 74085 262625 74113
rect 262653 74085 262687 74113
rect 262715 74085 262749 74113
rect 262777 74085 262811 74113
rect 262839 74085 262887 74113
rect 262577 74051 262887 74085
rect 262577 74023 262625 74051
rect 262653 74023 262687 74051
rect 262715 74023 262749 74051
rect 262777 74023 262811 74051
rect 262839 74023 262887 74051
rect 262577 73989 262887 74023
rect 262577 73961 262625 73989
rect 262653 73961 262687 73989
rect 262715 73961 262749 73989
rect 262777 73961 262811 73989
rect 262839 73961 262887 73989
rect 262577 65175 262887 73961
rect 262577 65147 262625 65175
rect 262653 65147 262687 65175
rect 262715 65147 262749 65175
rect 262777 65147 262811 65175
rect 262839 65147 262887 65175
rect 262577 65113 262887 65147
rect 262577 65085 262625 65113
rect 262653 65085 262687 65113
rect 262715 65085 262749 65113
rect 262777 65085 262811 65113
rect 262839 65085 262887 65113
rect 262577 65051 262887 65085
rect 262577 65023 262625 65051
rect 262653 65023 262687 65051
rect 262715 65023 262749 65051
rect 262777 65023 262811 65051
rect 262839 65023 262887 65051
rect 262577 64989 262887 65023
rect 262577 64961 262625 64989
rect 262653 64961 262687 64989
rect 262715 64961 262749 64989
rect 262777 64961 262811 64989
rect 262839 64961 262887 64989
rect 262577 56175 262887 64961
rect 262577 56147 262625 56175
rect 262653 56147 262687 56175
rect 262715 56147 262749 56175
rect 262777 56147 262811 56175
rect 262839 56147 262887 56175
rect 262577 56113 262887 56147
rect 262577 56085 262625 56113
rect 262653 56085 262687 56113
rect 262715 56085 262749 56113
rect 262777 56085 262811 56113
rect 262839 56085 262887 56113
rect 262577 56051 262887 56085
rect 262577 56023 262625 56051
rect 262653 56023 262687 56051
rect 262715 56023 262749 56051
rect 262777 56023 262811 56051
rect 262839 56023 262887 56051
rect 262577 55989 262887 56023
rect 262577 55961 262625 55989
rect 262653 55961 262687 55989
rect 262715 55961 262749 55989
rect 262777 55961 262811 55989
rect 262839 55961 262887 55989
rect 262577 47175 262887 55961
rect 262577 47147 262625 47175
rect 262653 47147 262687 47175
rect 262715 47147 262749 47175
rect 262777 47147 262811 47175
rect 262839 47147 262887 47175
rect 262577 47113 262887 47147
rect 262577 47085 262625 47113
rect 262653 47085 262687 47113
rect 262715 47085 262749 47113
rect 262777 47085 262811 47113
rect 262839 47085 262887 47113
rect 262577 47051 262887 47085
rect 262577 47023 262625 47051
rect 262653 47023 262687 47051
rect 262715 47023 262749 47051
rect 262777 47023 262811 47051
rect 262839 47023 262887 47051
rect 262577 46989 262887 47023
rect 262577 46961 262625 46989
rect 262653 46961 262687 46989
rect 262715 46961 262749 46989
rect 262777 46961 262811 46989
rect 262839 46961 262887 46989
rect 262577 38175 262887 46961
rect 262577 38147 262625 38175
rect 262653 38147 262687 38175
rect 262715 38147 262749 38175
rect 262777 38147 262811 38175
rect 262839 38147 262887 38175
rect 262577 38113 262887 38147
rect 262577 38085 262625 38113
rect 262653 38085 262687 38113
rect 262715 38085 262749 38113
rect 262777 38085 262811 38113
rect 262839 38085 262887 38113
rect 262577 38051 262887 38085
rect 262577 38023 262625 38051
rect 262653 38023 262687 38051
rect 262715 38023 262749 38051
rect 262777 38023 262811 38051
rect 262839 38023 262887 38051
rect 262577 37989 262887 38023
rect 262577 37961 262625 37989
rect 262653 37961 262687 37989
rect 262715 37961 262749 37989
rect 262777 37961 262811 37989
rect 262839 37961 262887 37989
rect 262577 29175 262887 37961
rect 262577 29147 262625 29175
rect 262653 29147 262687 29175
rect 262715 29147 262749 29175
rect 262777 29147 262811 29175
rect 262839 29147 262887 29175
rect 262577 29113 262887 29147
rect 262577 29085 262625 29113
rect 262653 29085 262687 29113
rect 262715 29085 262749 29113
rect 262777 29085 262811 29113
rect 262839 29085 262887 29113
rect 262577 29051 262887 29085
rect 262577 29023 262625 29051
rect 262653 29023 262687 29051
rect 262715 29023 262749 29051
rect 262777 29023 262811 29051
rect 262839 29023 262887 29051
rect 262577 28989 262887 29023
rect 262577 28961 262625 28989
rect 262653 28961 262687 28989
rect 262715 28961 262749 28989
rect 262777 28961 262811 28989
rect 262839 28961 262887 28989
rect 262577 20175 262887 28961
rect 262577 20147 262625 20175
rect 262653 20147 262687 20175
rect 262715 20147 262749 20175
rect 262777 20147 262811 20175
rect 262839 20147 262887 20175
rect 262577 20113 262887 20147
rect 262577 20085 262625 20113
rect 262653 20085 262687 20113
rect 262715 20085 262749 20113
rect 262777 20085 262811 20113
rect 262839 20085 262887 20113
rect 262577 20051 262887 20085
rect 262577 20023 262625 20051
rect 262653 20023 262687 20051
rect 262715 20023 262749 20051
rect 262777 20023 262811 20051
rect 262839 20023 262887 20051
rect 262577 19989 262887 20023
rect 262577 19961 262625 19989
rect 262653 19961 262687 19989
rect 262715 19961 262749 19989
rect 262777 19961 262811 19989
rect 262839 19961 262887 19989
rect 262577 11175 262887 19961
rect 262577 11147 262625 11175
rect 262653 11147 262687 11175
rect 262715 11147 262749 11175
rect 262777 11147 262811 11175
rect 262839 11147 262887 11175
rect 262577 11113 262887 11147
rect 262577 11085 262625 11113
rect 262653 11085 262687 11113
rect 262715 11085 262749 11113
rect 262777 11085 262811 11113
rect 262839 11085 262887 11113
rect 262577 11051 262887 11085
rect 262577 11023 262625 11051
rect 262653 11023 262687 11051
rect 262715 11023 262749 11051
rect 262777 11023 262811 11051
rect 262839 11023 262887 11051
rect 262577 10989 262887 11023
rect 262577 10961 262625 10989
rect 262653 10961 262687 10989
rect 262715 10961 262749 10989
rect 262777 10961 262811 10989
rect 262839 10961 262887 10989
rect 262577 2175 262887 10961
rect 262577 2147 262625 2175
rect 262653 2147 262687 2175
rect 262715 2147 262749 2175
rect 262777 2147 262811 2175
rect 262839 2147 262887 2175
rect 262577 2113 262887 2147
rect 262577 2085 262625 2113
rect 262653 2085 262687 2113
rect 262715 2085 262749 2113
rect 262777 2085 262811 2113
rect 262839 2085 262887 2113
rect 262577 2051 262887 2085
rect 262577 2023 262625 2051
rect 262653 2023 262687 2051
rect 262715 2023 262749 2051
rect 262777 2023 262811 2051
rect 262839 2023 262887 2051
rect 262577 1989 262887 2023
rect 262577 1961 262625 1989
rect 262653 1961 262687 1989
rect 262715 1961 262749 1989
rect 262777 1961 262811 1989
rect 262839 1961 262887 1989
rect 262577 -80 262887 1961
rect 262577 -108 262625 -80
rect 262653 -108 262687 -80
rect 262715 -108 262749 -80
rect 262777 -108 262811 -80
rect 262839 -108 262887 -80
rect 262577 -142 262887 -108
rect 262577 -170 262625 -142
rect 262653 -170 262687 -142
rect 262715 -170 262749 -142
rect 262777 -170 262811 -142
rect 262839 -170 262887 -142
rect 262577 -204 262887 -170
rect 262577 -232 262625 -204
rect 262653 -232 262687 -204
rect 262715 -232 262749 -204
rect 262777 -232 262811 -204
rect 262839 -232 262887 -204
rect 262577 -266 262887 -232
rect 262577 -294 262625 -266
rect 262653 -294 262687 -266
rect 262715 -294 262749 -266
rect 262777 -294 262811 -266
rect 262839 -294 262887 -266
rect 262577 -822 262887 -294
rect 264437 299086 264747 299134
rect 264437 299058 264485 299086
rect 264513 299058 264547 299086
rect 264575 299058 264609 299086
rect 264637 299058 264671 299086
rect 264699 299058 264747 299086
rect 264437 299024 264747 299058
rect 264437 298996 264485 299024
rect 264513 298996 264547 299024
rect 264575 298996 264609 299024
rect 264637 298996 264671 299024
rect 264699 298996 264747 299024
rect 264437 298962 264747 298996
rect 264437 298934 264485 298962
rect 264513 298934 264547 298962
rect 264575 298934 264609 298962
rect 264637 298934 264671 298962
rect 264699 298934 264747 298962
rect 264437 298900 264747 298934
rect 264437 298872 264485 298900
rect 264513 298872 264547 298900
rect 264575 298872 264609 298900
rect 264637 298872 264671 298900
rect 264699 298872 264747 298900
rect 264437 293175 264747 298872
rect 264437 293147 264485 293175
rect 264513 293147 264547 293175
rect 264575 293147 264609 293175
rect 264637 293147 264671 293175
rect 264699 293147 264747 293175
rect 264437 293113 264747 293147
rect 264437 293085 264485 293113
rect 264513 293085 264547 293113
rect 264575 293085 264609 293113
rect 264637 293085 264671 293113
rect 264699 293085 264747 293113
rect 264437 293051 264747 293085
rect 264437 293023 264485 293051
rect 264513 293023 264547 293051
rect 264575 293023 264609 293051
rect 264637 293023 264671 293051
rect 264699 293023 264747 293051
rect 264437 292989 264747 293023
rect 264437 292961 264485 292989
rect 264513 292961 264547 292989
rect 264575 292961 264609 292989
rect 264637 292961 264671 292989
rect 264699 292961 264747 292989
rect 264437 284175 264747 292961
rect 264437 284147 264485 284175
rect 264513 284147 264547 284175
rect 264575 284147 264609 284175
rect 264637 284147 264671 284175
rect 264699 284147 264747 284175
rect 264437 284113 264747 284147
rect 264437 284085 264485 284113
rect 264513 284085 264547 284113
rect 264575 284085 264609 284113
rect 264637 284085 264671 284113
rect 264699 284085 264747 284113
rect 264437 284051 264747 284085
rect 264437 284023 264485 284051
rect 264513 284023 264547 284051
rect 264575 284023 264609 284051
rect 264637 284023 264671 284051
rect 264699 284023 264747 284051
rect 264437 283989 264747 284023
rect 264437 283961 264485 283989
rect 264513 283961 264547 283989
rect 264575 283961 264609 283989
rect 264637 283961 264671 283989
rect 264699 283961 264747 283989
rect 264437 275175 264747 283961
rect 264437 275147 264485 275175
rect 264513 275147 264547 275175
rect 264575 275147 264609 275175
rect 264637 275147 264671 275175
rect 264699 275147 264747 275175
rect 264437 275113 264747 275147
rect 264437 275085 264485 275113
rect 264513 275085 264547 275113
rect 264575 275085 264609 275113
rect 264637 275085 264671 275113
rect 264699 275085 264747 275113
rect 264437 275051 264747 275085
rect 264437 275023 264485 275051
rect 264513 275023 264547 275051
rect 264575 275023 264609 275051
rect 264637 275023 264671 275051
rect 264699 275023 264747 275051
rect 264437 274989 264747 275023
rect 264437 274961 264485 274989
rect 264513 274961 264547 274989
rect 264575 274961 264609 274989
rect 264637 274961 264671 274989
rect 264699 274961 264747 274989
rect 264437 266175 264747 274961
rect 264437 266147 264485 266175
rect 264513 266147 264547 266175
rect 264575 266147 264609 266175
rect 264637 266147 264671 266175
rect 264699 266147 264747 266175
rect 264437 266113 264747 266147
rect 264437 266085 264485 266113
rect 264513 266085 264547 266113
rect 264575 266085 264609 266113
rect 264637 266085 264671 266113
rect 264699 266085 264747 266113
rect 264437 266051 264747 266085
rect 264437 266023 264485 266051
rect 264513 266023 264547 266051
rect 264575 266023 264609 266051
rect 264637 266023 264671 266051
rect 264699 266023 264747 266051
rect 264437 265989 264747 266023
rect 264437 265961 264485 265989
rect 264513 265961 264547 265989
rect 264575 265961 264609 265989
rect 264637 265961 264671 265989
rect 264699 265961 264747 265989
rect 264437 257175 264747 265961
rect 264437 257147 264485 257175
rect 264513 257147 264547 257175
rect 264575 257147 264609 257175
rect 264637 257147 264671 257175
rect 264699 257147 264747 257175
rect 264437 257113 264747 257147
rect 264437 257085 264485 257113
rect 264513 257085 264547 257113
rect 264575 257085 264609 257113
rect 264637 257085 264671 257113
rect 264699 257085 264747 257113
rect 264437 257051 264747 257085
rect 264437 257023 264485 257051
rect 264513 257023 264547 257051
rect 264575 257023 264609 257051
rect 264637 257023 264671 257051
rect 264699 257023 264747 257051
rect 264437 256989 264747 257023
rect 264437 256961 264485 256989
rect 264513 256961 264547 256989
rect 264575 256961 264609 256989
rect 264637 256961 264671 256989
rect 264699 256961 264747 256989
rect 264437 248175 264747 256961
rect 264437 248147 264485 248175
rect 264513 248147 264547 248175
rect 264575 248147 264609 248175
rect 264637 248147 264671 248175
rect 264699 248147 264747 248175
rect 264437 248113 264747 248147
rect 264437 248085 264485 248113
rect 264513 248085 264547 248113
rect 264575 248085 264609 248113
rect 264637 248085 264671 248113
rect 264699 248085 264747 248113
rect 264437 248051 264747 248085
rect 264437 248023 264485 248051
rect 264513 248023 264547 248051
rect 264575 248023 264609 248051
rect 264637 248023 264671 248051
rect 264699 248023 264747 248051
rect 264437 247989 264747 248023
rect 264437 247961 264485 247989
rect 264513 247961 264547 247989
rect 264575 247961 264609 247989
rect 264637 247961 264671 247989
rect 264699 247961 264747 247989
rect 264437 239175 264747 247961
rect 264437 239147 264485 239175
rect 264513 239147 264547 239175
rect 264575 239147 264609 239175
rect 264637 239147 264671 239175
rect 264699 239147 264747 239175
rect 264437 239113 264747 239147
rect 264437 239085 264485 239113
rect 264513 239085 264547 239113
rect 264575 239085 264609 239113
rect 264637 239085 264671 239113
rect 264699 239085 264747 239113
rect 264437 239051 264747 239085
rect 264437 239023 264485 239051
rect 264513 239023 264547 239051
rect 264575 239023 264609 239051
rect 264637 239023 264671 239051
rect 264699 239023 264747 239051
rect 264437 238989 264747 239023
rect 264437 238961 264485 238989
rect 264513 238961 264547 238989
rect 264575 238961 264609 238989
rect 264637 238961 264671 238989
rect 264699 238961 264747 238989
rect 264437 230175 264747 238961
rect 264437 230147 264485 230175
rect 264513 230147 264547 230175
rect 264575 230147 264609 230175
rect 264637 230147 264671 230175
rect 264699 230147 264747 230175
rect 264437 230113 264747 230147
rect 264437 230085 264485 230113
rect 264513 230085 264547 230113
rect 264575 230085 264609 230113
rect 264637 230085 264671 230113
rect 264699 230085 264747 230113
rect 264437 230051 264747 230085
rect 264437 230023 264485 230051
rect 264513 230023 264547 230051
rect 264575 230023 264609 230051
rect 264637 230023 264671 230051
rect 264699 230023 264747 230051
rect 264437 229989 264747 230023
rect 264437 229961 264485 229989
rect 264513 229961 264547 229989
rect 264575 229961 264609 229989
rect 264637 229961 264671 229989
rect 264699 229961 264747 229989
rect 264437 221175 264747 229961
rect 264437 221147 264485 221175
rect 264513 221147 264547 221175
rect 264575 221147 264609 221175
rect 264637 221147 264671 221175
rect 264699 221147 264747 221175
rect 264437 221113 264747 221147
rect 264437 221085 264485 221113
rect 264513 221085 264547 221113
rect 264575 221085 264609 221113
rect 264637 221085 264671 221113
rect 264699 221085 264747 221113
rect 264437 221051 264747 221085
rect 264437 221023 264485 221051
rect 264513 221023 264547 221051
rect 264575 221023 264609 221051
rect 264637 221023 264671 221051
rect 264699 221023 264747 221051
rect 264437 220989 264747 221023
rect 264437 220961 264485 220989
rect 264513 220961 264547 220989
rect 264575 220961 264609 220989
rect 264637 220961 264671 220989
rect 264699 220961 264747 220989
rect 264437 212175 264747 220961
rect 264437 212147 264485 212175
rect 264513 212147 264547 212175
rect 264575 212147 264609 212175
rect 264637 212147 264671 212175
rect 264699 212147 264747 212175
rect 264437 212113 264747 212147
rect 264437 212085 264485 212113
rect 264513 212085 264547 212113
rect 264575 212085 264609 212113
rect 264637 212085 264671 212113
rect 264699 212085 264747 212113
rect 264437 212051 264747 212085
rect 264437 212023 264485 212051
rect 264513 212023 264547 212051
rect 264575 212023 264609 212051
rect 264637 212023 264671 212051
rect 264699 212023 264747 212051
rect 264437 211989 264747 212023
rect 264437 211961 264485 211989
rect 264513 211961 264547 211989
rect 264575 211961 264609 211989
rect 264637 211961 264671 211989
rect 264699 211961 264747 211989
rect 264437 203175 264747 211961
rect 264437 203147 264485 203175
rect 264513 203147 264547 203175
rect 264575 203147 264609 203175
rect 264637 203147 264671 203175
rect 264699 203147 264747 203175
rect 264437 203113 264747 203147
rect 264437 203085 264485 203113
rect 264513 203085 264547 203113
rect 264575 203085 264609 203113
rect 264637 203085 264671 203113
rect 264699 203085 264747 203113
rect 264437 203051 264747 203085
rect 264437 203023 264485 203051
rect 264513 203023 264547 203051
rect 264575 203023 264609 203051
rect 264637 203023 264671 203051
rect 264699 203023 264747 203051
rect 264437 202989 264747 203023
rect 264437 202961 264485 202989
rect 264513 202961 264547 202989
rect 264575 202961 264609 202989
rect 264637 202961 264671 202989
rect 264699 202961 264747 202989
rect 264437 194175 264747 202961
rect 264437 194147 264485 194175
rect 264513 194147 264547 194175
rect 264575 194147 264609 194175
rect 264637 194147 264671 194175
rect 264699 194147 264747 194175
rect 264437 194113 264747 194147
rect 264437 194085 264485 194113
rect 264513 194085 264547 194113
rect 264575 194085 264609 194113
rect 264637 194085 264671 194113
rect 264699 194085 264747 194113
rect 264437 194051 264747 194085
rect 264437 194023 264485 194051
rect 264513 194023 264547 194051
rect 264575 194023 264609 194051
rect 264637 194023 264671 194051
rect 264699 194023 264747 194051
rect 264437 193989 264747 194023
rect 264437 193961 264485 193989
rect 264513 193961 264547 193989
rect 264575 193961 264609 193989
rect 264637 193961 264671 193989
rect 264699 193961 264747 193989
rect 264437 185175 264747 193961
rect 264437 185147 264485 185175
rect 264513 185147 264547 185175
rect 264575 185147 264609 185175
rect 264637 185147 264671 185175
rect 264699 185147 264747 185175
rect 264437 185113 264747 185147
rect 264437 185085 264485 185113
rect 264513 185085 264547 185113
rect 264575 185085 264609 185113
rect 264637 185085 264671 185113
rect 264699 185085 264747 185113
rect 264437 185051 264747 185085
rect 264437 185023 264485 185051
rect 264513 185023 264547 185051
rect 264575 185023 264609 185051
rect 264637 185023 264671 185051
rect 264699 185023 264747 185051
rect 264437 184989 264747 185023
rect 264437 184961 264485 184989
rect 264513 184961 264547 184989
rect 264575 184961 264609 184989
rect 264637 184961 264671 184989
rect 264699 184961 264747 184989
rect 264437 176175 264747 184961
rect 264437 176147 264485 176175
rect 264513 176147 264547 176175
rect 264575 176147 264609 176175
rect 264637 176147 264671 176175
rect 264699 176147 264747 176175
rect 264437 176113 264747 176147
rect 264437 176085 264485 176113
rect 264513 176085 264547 176113
rect 264575 176085 264609 176113
rect 264637 176085 264671 176113
rect 264699 176085 264747 176113
rect 264437 176051 264747 176085
rect 264437 176023 264485 176051
rect 264513 176023 264547 176051
rect 264575 176023 264609 176051
rect 264637 176023 264671 176051
rect 264699 176023 264747 176051
rect 264437 175989 264747 176023
rect 264437 175961 264485 175989
rect 264513 175961 264547 175989
rect 264575 175961 264609 175989
rect 264637 175961 264671 175989
rect 264699 175961 264747 175989
rect 264437 167175 264747 175961
rect 264437 167147 264485 167175
rect 264513 167147 264547 167175
rect 264575 167147 264609 167175
rect 264637 167147 264671 167175
rect 264699 167147 264747 167175
rect 264437 167113 264747 167147
rect 264437 167085 264485 167113
rect 264513 167085 264547 167113
rect 264575 167085 264609 167113
rect 264637 167085 264671 167113
rect 264699 167085 264747 167113
rect 264437 167051 264747 167085
rect 264437 167023 264485 167051
rect 264513 167023 264547 167051
rect 264575 167023 264609 167051
rect 264637 167023 264671 167051
rect 264699 167023 264747 167051
rect 264437 166989 264747 167023
rect 264437 166961 264485 166989
rect 264513 166961 264547 166989
rect 264575 166961 264609 166989
rect 264637 166961 264671 166989
rect 264699 166961 264747 166989
rect 264437 158175 264747 166961
rect 264437 158147 264485 158175
rect 264513 158147 264547 158175
rect 264575 158147 264609 158175
rect 264637 158147 264671 158175
rect 264699 158147 264747 158175
rect 264437 158113 264747 158147
rect 264437 158085 264485 158113
rect 264513 158085 264547 158113
rect 264575 158085 264609 158113
rect 264637 158085 264671 158113
rect 264699 158085 264747 158113
rect 264437 158051 264747 158085
rect 264437 158023 264485 158051
rect 264513 158023 264547 158051
rect 264575 158023 264609 158051
rect 264637 158023 264671 158051
rect 264699 158023 264747 158051
rect 264437 157989 264747 158023
rect 264437 157961 264485 157989
rect 264513 157961 264547 157989
rect 264575 157961 264609 157989
rect 264637 157961 264671 157989
rect 264699 157961 264747 157989
rect 264437 149175 264747 157961
rect 264437 149147 264485 149175
rect 264513 149147 264547 149175
rect 264575 149147 264609 149175
rect 264637 149147 264671 149175
rect 264699 149147 264747 149175
rect 264437 149113 264747 149147
rect 264437 149085 264485 149113
rect 264513 149085 264547 149113
rect 264575 149085 264609 149113
rect 264637 149085 264671 149113
rect 264699 149085 264747 149113
rect 264437 149051 264747 149085
rect 264437 149023 264485 149051
rect 264513 149023 264547 149051
rect 264575 149023 264609 149051
rect 264637 149023 264671 149051
rect 264699 149023 264747 149051
rect 264437 148989 264747 149023
rect 264437 148961 264485 148989
rect 264513 148961 264547 148989
rect 264575 148961 264609 148989
rect 264637 148961 264671 148989
rect 264699 148961 264747 148989
rect 264437 140175 264747 148961
rect 264437 140147 264485 140175
rect 264513 140147 264547 140175
rect 264575 140147 264609 140175
rect 264637 140147 264671 140175
rect 264699 140147 264747 140175
rect 264437 140113 264747 140147
rect 264437 140085 264485 140113
rect 264513 140085 264547 140113
rect 264575 140085 264609 140113
rect 264637 140085 264671 140113
rect 264699 140085 264747 140113
rect 264437 140051 264747 140085
rect 264437 140023 264485 140051
rect 264513 140023 264547 140051
rect 264575 140023 264609 140051
rect 264637 140023 264671 140051
rect 264699 140023 264747 140051
rect 264437 139989 264747 140023
rect 264437 139961 264485 139989
rect 264513 139961 264547 139989
rect 264575 139961 264609 139989
rect 264637 139961 264671 139989
rect 264699 139961 264747 139989
rect 264437 131175 264747 139961
rect 264437 131147 264485 131175
rect 264513 131147 264547 131175
rect 264575 131147 264609 131175
rect 264637 131147 264671 131175
rect 264699 131147 264747 131175
rect 264437 131113 264747 131147
rect 264437 131085 264485 131113
rect 264513 131085 264547 131113
rect 264575 131085 264609 131113
rect 264637 131085 264671 131113
rect 264699 131085 264747 131113
rect 264437 131051 264747 131085
rect 264437 131023 264485 131051
rect 264513 131023 264547 131051
rect 264575 131023 264609 131051
rect 264637 131023 264671 131051
rect 264699 131023 264747 131051
rect 264437 130989 264747 131023
rect 264437 130961 264485 130989
rect 264513 130961 264547 130989
rect 264575 130961 264609 130989
rect 264637 130961 264671 130989
rect 264699 130961 264747 130989
rect 264437 122175 264747 130961
rect 264437 122147 264485 122175
rect 264513 122147 264547 122175
rect 264575 122147 264609 122175
rect 264637 122147 264671 122175
rect 264699 122147 264747 122175
rect 264437 122113 264747 122147
rect 264437 122085 264485 122113
rect 264513 122085 264547 122113
rect 264575 122085 264609 122113
rect 264637 122085 264671 122113
rect 264699 122085 264747 122113
rect 264437 122051 264747 122085
rect 264437 122023 264485 122051
rect 264513 122023 264547 122051
rect 264575 122023 264609 122051
rect 264637 122023 264671 122051
rect 264699 122023 264747 122051
rect 264437 121989 264747 122023
rect 264437 121961 264485 121989
rect 264513 121961 264547 121989
rect 264575 121961 264609 121989
rect 264637 121961 264671 121989
rect 264699 121961 264747 121989
rect 264437 113175 264747 121961
rect 264437 113147 264485 113175
rect 264513 113147 264547 113175
rect 264575 113147 264609 113175
rect 264637 113147 264671 113175
rect 264699 113147 264747 113175
rect 264437 113113 264747 113147
rect 264437 113085 264485 113113
rect 264513 113085 264547 113113
rect 264575 113085 264609 113113
rect 264637 113085 264671 113113
rect 264699 113085 264747 113113
rect 264437 113051 264747 113085
rect 264437 113023 264485 113051
rect 264513 113023 264547 113051
rect 264575 113023 264609 113051
rect 264637 113023 264671 113051
rect 264699 113023 264747 113051
rect 264437 112989 264747 113023
rect 264437 112961 264485 112989
rect 264513 112961 264547 112989
rect 264575 112961 264609 112989
rect 264637 112961 264671 112989
rect 264699 112961 264747 112989
rect 264437 104175 264747 112961
rect 264437 104147 264485 104175
rect 264513 104147 264547 104175
rect 264575 104147 264609 104175
rect 264637 104147 264671 104175
rect 264699 104147 264747 104175
rect 264437 104113 264747 104147
rect 264437 104085 264485 104113
rect 264513 104085 264547 104113
rect 264575 104085 264609 104113
rect 264637 104085 264671 104113
rect 264699 104085 264747 104113
rect 264437 104051 264747 104085
rect 264437 104023 264485 104051
rect 264513 104023 264547 104051
rect 264575 104023 264609 104051
rect 264637 104023 264671 104051
rect 264699 104023 264747 104051
rect 264437 103989 264747 104023
rect 264437 103961 264485 103989
rect 264513 103961 264547 103989
rect 264575 103961 264609 103989
rect 264637 103961 264671 103989
rect 264699 103961 264747 103989
rect 264437 95175 264747 103961
rect 264437 95147 264485 95175
rect 264513 95147 264547 95175
rect 264575 95147 264609 95175
rect 264637 95147 264671 95175
rect 264699 95147 264747 95175
rect 264437 95113 264747 95147
rect 264437 95085 264485 95113
rect 264513 95085 264547 95113
rect 264575 95085 264609 95113
rect 264637 95085 264671 95113
rect 264699 95085 264747 95113
rect 264437 95051 264747 95085
rect 264437 95023 264485 95051
rect 264513 95023 264547 95051
rect 264575 95023 264609 95051
rect 264637 95023 264671 95051
rect 264699 95023 264747 95051
rect 264437 94989 264747 95023
rect 264437 94961 264485 94989
rect 264513 94961 264547 94989
rect 264575 94961 264609 94989
rect 264637 94961 264671 94989
rect 264699 94961 264747 94989
rect 264437 86175 264747 94961
rect 264437 86147 264485 86175
rect 264513 86147 264547 86175
rect 264575 86147 264609 86175
rect 264637 86147 264671 86175
rect 264699 86147 264747 86175
rect 264437 86113 264747 86147
rect 264437 86085 264485 86113
rect 264513 86085 264547 86113
rect 264575 86085 264609 86113
rect 264637 86085 264671 86113
rect 264699 86085 264747 86113
rect 264437 86051 264747 86085
rect 264437 86023 264485 86051
rect 264513 86023 264547 86051
rect 264575 86023 264609 86051
rect 264637 86023 264671 86051
rect 264699 86023 264747 86051
rect 264437 85989 264747 86023
rect 264437 85961 264485 85989
rect 264513 85961 264547 85989
rect 264575 85961 264609 85989
rect 264637 85961 264671 85989
rect 264699 85961 264747 85989
rect 264437 77175 264747 85961
rect 264437 77147 264485 77175
rect 264513 77147 264547 77175
rect 264575 77147 264609 77175
rect 264637 77147 264671 77175
rect 264699 77147 264747 77175
rect 264437 77113 264747 77147
rect 264437 77085 264485 77113
rect 264513 77085 264547 77113
rect 264575 77085 264609 77113
rect 264637 77085 264671 77113
rect 264699 77085 264747 77113
rect 264437 77051 264747 77085
rect 264437 77023 264485 77051
rect 264513 77023 264547 77051
rect 264575 77023 264609 77051
rect 264637 77023 264671 77051
rect 264699 77023 264747 77051
rect 264437 76989 264747 77023
rect 264437 76961 264485 76989
rect 264513 76961 264547 76989
rect 264575 76961 264609 76989
rect 264637 76961 264671 76989
rect 264699 76961 264747 76989
rect 264437 68175 264747 76961
rect 264437 68147 264485 68175
rect 264513 68147 264547 68175
rect 264575 68147 264609 68175
rect 264637 68147 264671 68175
rect 264699 68147 264747 68175
rect 264437 68113 264747 68147
rect 264437 68085 264485 68113
rect 264513 68085 264547 68113
rect 264575 68085 264609 68113
rect 264637 68085 264671 68113
rect 264699 68085 264747 68113
rect 264437 68051 264747 68085
rect 264437 68023 264485 68051
rect 264513 68023 264547 68051
rect 264575 68023 264609 68051
rect 264637 68023 264671 68051
rect 264699 68023 264747 68051
rect 264437 67989 264747 68023
rect 264437 67961 264485 67989
rect 264513 67961 264547 67989
rect 264575 67961 264609 67989
rect 264637 67961 264671 67989
rect 264699 67961 264747 67989
rect 264437 59175 264747 67961
rect 264437 59147 264485 59175
rect 264513 59147 264547 59175
rect 264575 59147 264609 59175
rect 264637 59147 264671 59175
rect 264699 59147 264747 59175
rect 264437 59113 264747 59147
rect 264437 59085 264485 59113
rect 264513 59085 264547 59113
rect 264575 59085 264609 59113
rect 264637 59085 264671 59113
rect 264699 59085 264747 59113
rect 264437 59051 264747 59085
rect 264437 59023 264485 59051
rect 264513 59023 264547 59051
rect 264575 59023 264609 59051
rect 264637 59023 264671 59051
rect 264699 59023 264747 59051
rect 264437 58989 264747 59023
rect 264437 58961 264485 58989
rect 264513 58961 264547 58989
rect 264575 58961 264609 58989
rect 264637 58961 264671 58989
rect 264699 58961 264747 58989
rect 264437 50175 264747 58961
rect 264437 50147 264485 50175
rect 264513 50147 264547 50175
rect 264575 50147 264609 50175
rect 264637 50147 264671 50175
rect 264699 50147 264747 50175
rect 264437 50113 264747 50147
rect 264437 50085 264485 50113
rect 264513 50085 264547 50113
rect 264575 50085 264609 50113
rect 264637 50085 264671 50113
rect 264699 50085 264747 50113
rect 264437 50051 264747 50085
rect 264437 50023 264485 50051
rect 264513 50023 264547 50051
rect 264575 50023 264609 50051
rect 264637 50023 264671 50051
rect 264699 50023 264747 50051
rect 264437 49989 264747 50023
rect 264437 49961 264485 49989
rect 264513 49961 264547 49989
rect 264575 49961 264609 49989
rect 264637 49961 264671 49989
rect 264699 49961 264747 49989
rect 264437 41175 264747 49961
rect 264437 41147 264485 41175
rect 264513 41147 264547 41175
rect 264575 41147 264609 41175
rect 264637 41147 264671 41175
rect 264699 41147 264747 41175
rect 264437 41113 264747 41147
rect 264437 41085 264485 41113
rect 264513 41085 264547 41113
rect 264575 41085 264609 41113
rect 264637 41085 264671 41113
rect 264699 41085 264747 41113
rect 264437 41051 264747 41085
rect 264437 41023 264485 41051
rect 264513 41023 264547 41051
rect 264575 41023 264609 41051
rect 264637 41023 264671 41051
rect 264699 41023 264747 41051
rect 264437 40989 264747 41023
rect 264437 40961 264485 40989
rect 264513 40961 264547 40989
rect 264575 40961 264609 40989
rect 264637 40961 264671 40989
rect 264699 40961 264747 40989
rect 264437 32175 264747 40961
rect 264437 32147 264485 32175
rect 264513 32147 264547 32175
rect 264575 32147 264609 32175
rect 264637 32147 264671 32175
rect 264699 32147 264747 32175
rect 264437 32113 264747 32147
rect 264437 32085 264485 32113
rect 264513 32085 264547 32113
rect 264575 32085 264609 32113
rect 264637 32085 264671 32113
rect 264699 32085 264747 32113
rect 264437 32051 264747 32085
rect 264437 32023 264485 32051
rect 264513 32023 264547 32051
rect 264575 32023 264609 32051
rect 264637 32023 264671 32051
rect 264699 32023 264747 32051
rect 264437 31989 264747 32023
rect 264437 31961 264485 31989
rect 264513 31961 264547 31989
rect 264575 31961 264609 31989
rect 264637 31961 264671 31989
rect 264699 31961 264747 31989
rect 264437 23175 264747 31961
rect 264437 23147 264485 23175
rect 264513 23147 264547 23175
rect 264575 23147 264609 23175
rect 264637 23147 264671 23175
rect 264699 23147 264747 23175
rect 264437 23113 264747 23147
rect 264437 23085 264485 23113
rect 264513 23085 264547 23113
rect 264575 23085 264609 23113
rect 264637 23085 264671 23113
rect 264699 23085 264747 23113
rect 264437 23051 264747 23085
rect 264437 23023 264485 23051
rect 264513 23023 264547 23051
rect 264575 23023 264609 23051
rect 264637 23023 264671 23051
rect 264699 23023 264747 23051
rect 264437 22989 264747 23023
rect 264437 22961 264485 22989
rect 264513 22961 264547 22989
rect 264575 22961 264609 22989
rect 264637 22961 264671 22989
rect 264699 22961 264747 22989
rect 264437 14175 264747 22961
rect 264437 14147 264485 14175
rect 264513 14147 264547 14175
rect 264575 14147 264609 14175
rect 264637 14147 264671 14175
rect 264699 14147 264747 14175
rect 264437 14113 264747 14147
rect 264437 14085 264485 14113
rect 264513 14085 264547 14113
rect 264575 14085 264609 14113
rect 264637 14085 264671 14113
rect 264699 14085 264747 14113
rect 264437 14051 264747 14085
rect 264437 14023 264485 14051
rect 264513 14023 264547 14051
rect 264575 14023 264609 14051
rect 264637 14023 264671 14051
rect 264699 14023 264747 14051
rect 264437 13989 264747 14023
rect 264437 13961 264485 13989
rect 264513 13961 264547 13989
rect 264575 13961 264609 13989
rect 264637 13961 264671 13989
rect 264699 13961 264747 13989
rect 264437 5175 264747 13961
rect 264437 5147 264485 5175
rect 264513 5147 264547 5175
rect 264575 5147 264609 5175
rect 264637 5147 264671 5175
rect 264699 5147 264747 5175
rect 264437 5113 264747 5147
rect 264437 5085 264485 5113
rect 264513 5085 264547 5113
rect 264575 5085 264609 5113
rect 264637 5085 264671 5113
rect 264699 5085 264747 5113
rect 264437 5051 264747 5085
rect 264437 5023 264485 5051
rect 264513 5023 264547 5051
rect 264575 5023 264609 5051
rect 264637 5023 264671 5051
rect 264699 5023 264747 5051
rect 264437 4989 264747 5023
rect 264437 4961 264485 4989
rect 264513 4961 264547 4989
rect 264575 4961 264609 4989
rect 264637 4961 264671 4989
rect 264699 4961 264747 4989
rect 264437 -560 264747 4961
rect 264437 -588 264485 -560
rect 264513 -588 264547 -560
rect 264575 -588 264609 -560
rect 264637 -588 264671 -560
rect 264699 -588 264747 -560
rect 264437 -622 264747 -588
rect 264437 -650 264485 -622
rect 264513 -650 264547 -622
rect 264575 -650 264609 -622
rect 264637 -650 264671 -622
rect 264699 -650 264747 -622
rect 264437 -684 264747 -650
rect 264437 -712 264485 -684
rect 264513 -712 264547 -684
rect 264575 -712 264609 -684
rect 264637 -712 264671 -684
rect 264699 -712 264747 -684
rect 264437 -746 264747 -712
rect 264437 -774 264485 -746
rect 264513 -774 264547 -746
rect 264575 -774 264609 -746
rect 264637 -774 264671 -746
rect 264699 -774 264747 -746
rect 264437 -822 264747 -774
rect 271577 298606 271887 299134
rect 271577 298578 271625 298606
rect 271653 298578 271687 298606
rect 271715 298578 271749 298606
rect 271777 298578 271811 298606
rect 271839 298578 271887 298606
rect 271577 298544 271887 298578
rect 271577 298516 271625 298544
rect 271653 298516 271687 298544
rect 271715 298516 271749 298544
rect 271777 298516 271811 298544
rect 271839 298516 271887 298544
rect 271577 298482 271887 298516
rect 271577 298454 271625 298482
rect 271653 298454 271687 298482
rect 271715 298454 271749 298482
rect 271777 298454 271811 298482
rect 271839 298454 271887 298482
rect 271577 298420 271887 298454
rect 271577 298392 271625 298420
rect 271653 298392 271687 298420
rect 271715 298392 271749 298420
rect 271777 298392 271811 298420
rect 271839 298392 271887 298420
rect 271577 290175 271887 298392
rect 271577 290147 271625 290175
rect 271653 290147 271687 290175
rect 271715 290147 271749 290175
rect 271777 290147 271811 290175
rect 271839 290147 271887 290175
rect 271577 290113 271887 290147
rect 271577 290085 271625 290113
rect 271653 290085 271687 290113
rect 271715 290085 271749 290113
rect 271777 290085 271811 290113
rect 271839 290085 271887 290113
rect 271577 290051 271887 290085
rect 271577 290023 271625 290051
rect 271653 290023 271687 290051
rect 271715 290023 271749 290051
rect 271777 290023 271811 290051
rect 271839 290023 271887 290051
rect 271577 289989 271887 290023
rect 271577 289961 271625 289989
rect 271653 289961 271687 289989
rect 271715 289961 271749 289989
rect 271777 289961 271811 289989
rect 271839 289961 271887 289989
rect 271577 281175 271887 289961
rect 271577 281147 271625 281175
rect 271653 281147 271687 281175
rect 271715 281147 271749 281175
rect 271777 281147 271811 281175
rect 271839 281147 271887 281175
rect 271577 281113 271887 281147
rect 271577 281085 271625 281113
rect 271653 281085 271687 281113
rect 271715 281085 271749 281113
rect 271777 281085 271811 281113
rect 271839 281085 271887 281113
rect 271577 281051 271887 281085
rect 271577 281023 271625 281051
rect 271653 281023 271687 281051
rect 271715 281023 271749 281051
rect 271777 281023 271811 281051
rect 271839 281023 271887 281051
rect 271577 280989 271887 281023
rect 271577 280961 271625 280989
rect 271653 280961 271687 280989
rect 271715 280961 271749 280989
rect 271777 280961 271811 280989
rect 271839 280961 271887 280989
rect 271577 272175 271887 280961
rect 271577 272147 271625 272175
rect 271653 272147 271687 272175
rect 271715 272147 271749 272175
rect 271777 272147 271811 272175
rect 271839 272147 271887 272175
rect 271577 272113 271887 272147
rect 271577 272085 271625 272113
rect 271653 272085 271687 272113
rect 271715 272085 271749 272113
rect 271777 272085 271811 272113
rect 271839 272085 271887 272113
rect 271577 272051 271887 272085
rect 271577 272023 271625 272051
rect 271653 272023 271687 272051
rect 271715 272023 271749 272051
rect 271777 272023 271811 272051
rect 271839 272023 271887 272051
rect 271577 271989 271887 272023
rect 271577 271961 271625 271989
rect 271653 271961 271687 271989
rect 271715 271961 271749 271989
rect 271777 271961 271811 271989
rect 271839 271961 271887 271989
rect 271577 263175 271887 271961
rect 271577 263147 271625 263175
rect 271653 263147 271687 263175
rect 271715 263147 271749 263175
rect 271777 263147 271811 263175
rect 271839 263147 271887 263175
rect 271577 263113 271887 263147
rect 271577 263085 271625 263113
rect 271653 263085 271687 263113
rect 271715 263085 271749 263113
rect 271777 263085 271811 263113
rect 271839 263085 271887 263113
rect 271577 263051 271887 263085
rect 271577 263023 271625 263051
rect 271653 263023 271687 263051
rect 271715 263023 271749 263051
rect 271777 263023 271811 263051
rect 271839 263023 271887 263051
rect 271577 262989 271887 263023
rect 271577 262961 271625 262989
rect 271653 262961 271687 262989
rect 271715 262961 271749 262989
rect 271777 262961 271811 262989
rect 271839 262961 271887 262989
rect 271577 254175 271887 262961
rect 271577 254147 271625 254175
rect 271653 254147 271687 254175
rect 271715 254147 271749 254175
rect 271777 254147 271811 254175
rect 271839 254147 271887 254175
rect 271577 254113 271887 254147
rect 271577 254085 271625 254113
rect 271653 254085 271687 254113
rect 271715 254085 271749 254113
rect 271777 254085 271811 254113
rect 271839 254085 271887 254113
rect 271577 254051 271887 254085
rect 271577 254023 271625 254051
rect 271653 254023 271687 254051
rect 271715 254023 271749 254051
rect 271777 254023 271811 254051
rect 271839 254023 271887 254051
rect 271577 253989 271887 254023
rect 271577 253961 271625 253989
rect 271653 253961 271687 253989
rect 271715 253961 271749 253989
rect 271777 253961 271811 253989
rect 271839 253961 271887 253989
rect 271577 245175 271887 253961
rect 271577 245147 271625 245175
rect 271653 245147 271687 245175
rect 271715 245147 271749 245175
rect 271777 245147 271811 245175
rect 271839 245147 271887 245175
rect 271577 245113 271887 245147
rect 271577 245085 271625 245113
rect 271653 245085 271687 245113
rect 271715 245085 271749 245113
rect 271777 245085 271811 245113
rect 271839 245085 271887 245113
rect 271577 245051 271887 245085
rect 271577 245023 271625 245051
rect 271653 245023 271687 245051
rect 271715 245023 271749 245051
rect 271777 245023 271811 245051
rect 271839 245023 271887 245051
rect 271577 244989 271887 245023
rect 271577 244961 271625 244989
rect 271653 244961 271687 244989
rect 271715 244961 271749 244989
rect 271777 244961 271811 244989
rect 271839 244961 271887 244989
rect 271577 236175 271887 244961
rect 271577 236147 271625 236175
rect 271653 236147 271687 236175
rect 271715 236147 271749 236175
rect 271777 236147 271811 236175
rect 271839 236147 271887 236175
rect 271577 236113 271887 236147
rect 271577 236085 271625 236113
rect 271653 236085 271687 236113
rect 271715 236085 271749 236113
rect 271777 236085 271811 236113
rect 271839 236085 271887 236113
rect 271577 236051 271887 236085
rect 271577 236023 271625 236051
rect 271653 236023 271687 236051
rect 271715 236023 271749 236051
rect 271777 236023 271811 236051
rect 271839 236023 271887 236051
rect 271577 235989 271887 236023
rect 271577 235961 271625 235989
rect 271653 235961 271687 235989
rect 271715 235961 271749 235989
rect 271777 235961 271811 235989
rect 271839 235961 271887 235989
rect 271577 227175 271887 235961
rect 271577 227147 271625 227175
rect 271653 227147 271687 227175
rect 271715 227147 271749 227175
rect 271777 227147 271811 227175
rect 271839 227147 271887 227175
rect 271577 227113 271887 227147
rect 271577 227085 271625 227113
rect 271653 227085 271687 227113
rect 271715 227085 271749 227113
rect 271777 227085 271811 227113
rect 271839 227085 271887 227113
rect 271577 227051 271887 227085
rect 271577 227023 271625 227051
rect 271653 227023 271687 227051
rect 271715 227023 271749 227051
rect 271777 227023 271811 227051
rect 271839 227023 271887 227051
rect 271577 226989 271887 227023
rect 271577 226961 271625 226989
rect 271653 226961 271687 226989
rect 271715 226961 271749 226989
rect 271777 226961 271811 226989
rect 271839 226961 271887 226989
rect 271577 218175 271887 226961
rect 271577 218147 271625 218175
rect 271653 218147 271687 218175
rect 271715 218147 271749 218175
rect 271777 218147 271811 218175
rect 271839 218147 271887 218175
rect 271577 218113 271887 218147
rect 271577 218085 271625 218113
rect 271653 218085 271687 218113
rect 271715 218085 271749 218113
rect 271777 218085 271811 218113
rect 271839 218085 271887 218113
rect 271577 218051 271887 218085
rect 271577 218023 271625 218051
rect 271653 218023 271687 218051
rect 271715 218023 271749 218051
rect 271777 218023 271811 218051
rect 271839 218023 271887 218051
rect 271577 217989 271887 218023
rect 271577 217961 271625 217989
rect 271653 217961 271687 217989
rect 271715 217961 271749 217989
rect 271777 217961 271811 217989
rect 271839 217961 271887 217989
rect 271577 209175 271887 217961
rect 271577 209147 271625 209175
rect 271653 209147 271687 209175
rect 271715 209147 271749 209175
rect 271777 209147 271811 209175
rect 271839 209147 271887 209175
rect 271577 209113 271887 209147
rect 271577 209085 271625 209113
rect 271653 209085 271687 209113
rect 271715 209085 271749 209113
rect 271777 209085 271811 209113
rect 271839 209085 271887 209113
rect 271577 209051 271887 209085
rect 271577 209023 271625 209051
rect 271653 209023 271687 209051
rect 271715 209023 271749 209051
rect 271777 209023 271811 209051
rect 271839 209023 271887 209051
rect 271577 208989 271887 209023
rect 271577 208961 271625 208989
rect 271653 208961 271687 208989
rect 271715 208961 271749 208989
rect 271777 208961 271811 208989
rect 271839 208961 271887 208989
rect 271577 200175 271887 208961
rect 271577 200147 271625 200175
rect 271653 200147 271687 200175
rect 271715 200147 271749 200175
rect 271777 200147 271811 200175
rect 271839 200147 271887 200175
rect 271577 200113 271887 200147
rect 271577 200085 271625 200113
rect 271653 200085 271687 200113
rect 271715 200085 271749 200113
rect 271777 200085 271811 200113
rect 271839 200085 271887 200113
rect 271577 200051 271887 200085
rect 271577 200023 271625 200051
rect 271653 200023 271687 200051
rect 271715 200023 271749 200051
rect 271777 200023 271811 200051
rect 271839 200023 271887 200051
rect 271577 199989 271887 200023
rect 271577 199961 271625 199989
rect 271653 199961 271687 199989
rect 271715 199961 271749 199989
rect 271777 199961 271811 199989
rect 271839 199961 271887 199989
rect 271577 191175 271887 199961
rect 271577 191147 271625 191175
rect 271653 191147 271687 191175
rect 271715 191147 271749 191175
rect 271777 191147 271811 191175
rect 271839 191147 271887 191175
rect 271577 191113 271887 191147
rect 271577 191085 271625 191113
rect 271653 191085 271687 191113
rect 271715 191085 271749 191113
rect 271777 191085 271811 191113
rect 271839 191085 271887 191113
rect 271577 191051 271887 191085
rect 271577 191023 271625 191051
rect 271653 191023 271687 191051
rect 271715 191023 271749 191051
rect 271777 191023 271811 191051
rect 271839 191023 271887 191051
rect 271577 190989 271887 191023
rect 271577 190961 271625 190989
rect 271653 190961 271687 190989
rect 271715 190961 271749 190989
rect 271777 190961 271811 190989
rect 271839 190961 271887 190989
rect 271577 182175 271887 190961
rect 271577 182147 271625 182175
rect 271653 182147 271687 182175
rect 271715 182147 271749 182175
rect 271777 182147 271811 182175
rect 271839 182147 271887 182175
rect 271577 182113 271887 182147
rect 271577 182085 271625 182113
rect 271653 182085 271687 182113
rect 271715 182085 271749 182113
rect 271777 182085 271811 182113
rect 271839 182085 271887 182113
rect 271577 182051 271887 182085
rect 271577 182023 271625 182051
rect 271653 182023 271687 182051
rect 271715 182023 271749 182051
rect 271777 182023 271811 182051
rect 271839 182023 271887 182051
rect 271577 181989 271887 182023
rect 271577 181961 271625 181989
rect 271653 181961 271687 181989
rect 271715 181961 271749 181989
rect 271777 181961 271811 181989
rect 271839 181961 271887 181989
rect 271577 173175 271887 181961
rect 271577 173147 271625 173175
rect 271653 173147 271687 173175
rect 271715 173147 271749 173175
rect 271777 173147 271811 173175
rect 271839 173147 271887 173175
rect 271577 173113 271887 173147
rect 271577 173085 271625 173113
rect 271653 173085 271687 173113
rect 271715 173085 271749 173113
rect 271777 173085 271811 173113
rect 271839 173085 271887 173113
rect 271577 173051 271887 173085
rect 271577 173023 271625 173051
rect 271653 173023 271687 173051
rect 271715 173023 271749 173051
rect 271777 173023 271811 173051
rect 271839 173023 271887 173051
rect 271577 172989 271887 173023
rect 271577 172961 271625 172989
rect 271653 172961 271687 172989
rect 271715 172961 271749 172989
rect 271777 172961 271811 172989
rect 271839 172961 271887 172989
rect 271577 164175 271887 172961
rect 271577 164147 271625 164175
rect 271653 164147 271687 164175
rect 271715 164147 271749 164175
rect 271777 164147 271811 164175
rect 271839 164147 271887 164175
rect 271577 164113 271887 164147
rect 271577 164085 271625 164113
rect 271653 164085 271687 164113
rect 271715 164085 271749 164113
rect 271777 164085 271811 164113
rect 271839 164085 271887 164113
rect 271577 164051 271887 164085
rect 271577 164023 271625 164051
rect 271653 164023 271687 164051
rect 271715 164023 271749 164051
rect 271777 164023 271811 164051
rect 271839 164023 271887 164051
rect 271577 163989 271887 164023
rect 271577 163961 271625 163989
rect 271653 163961 271687 163989
rect 271715 163961 271749 163989
rect 271777 163961 271811 163989
rect 271839 163961 271887 163989
rect 271577 155175 271887 163961
rect 271577 155147 271625 155175
rect 271653 155147 271687 155175
rect 271715 155147 271749 155175
rect 271777 155147 271811 155175
rect 271839 155147 271887 155175
rect 271577 155113 271887 155147
rect 271577 155085 271625 155113
rect 271653 155085 271687 155113
rect 271715 155085 271749 155113
rect 271777 155085 271811 155113
rect 271839 155085 271887 155113
rect 271577 155051 271887 155085
rect 271577 155023 271625 155051
rect 271653 155023 271687 155051
rect 271715 155023 271749 155051
rect 271777 155023 271811 155051
rect 271839 155023 271887 155051
rect 271577 154989 271887 155023
rect 271577 154961 271625 154989
rect 271653 154961 271687 154989
rect 271715 154961 271749 154989
rect 271777 154961 271811 154989
rect 271839 154961 271887 154989
rect 271577 146175 271887 154961
rect 271577 146147 271625 146175
rect 271653 146147 271687 146175
rect 271715 146147 271749 146175
rect 271777 146147 271811 146175
rect 271839 146147 271887 146175
rect 271577 146113 271887 146147
rect 271577 146085 271625 146113
rect 271653 146085 271687 146113
rect 271715 146085 271749 146113
rect 271777 146085 271811 146113
rect 271839 146085 271887 146113
rect 271577 146051 271887 146085
rect 271577 146023 271625 146051
rect 271653 146023 271687 146051
rect 271715 146023 271749 146051
rect 271777 146023 271811 146051
rect 271839 146023 271887 146051
rect 271577 145989 271887 146023
rect 271577 145961 271625 145989
rect 271653 145961 271687 145989
rect 271715 145961 271749 145989
rect 271777 145961 271811 145989
rect 271839 145961 271887 145989
rect 271577 137175 271887 145961
rect 271577 137147 271625 137175
rect 271653 137147 271687 137175
rect 271715 137147 271749 137175
rect 271777 137147 271811 137175
rect 271839 137147 271887 137175
rect 271577 137113 271887 137147
rect 271577 137085 271625 137113
rect 271653 137085 271687 137113
rect 271715 137085 271749 137113
rect 271777 137085 271811 137113
rect 271839 137085 271887 137113
rect 271577 137051 271887 137085
rect 271577 137023 271625 137051
rect 271653 137023 271687 137051
rect 271715 137023 271749 137051
rect 271777 137023 271811 137051
rect 271839 137023 271887 137051
rect 271577 136989 271887 137023
rect 271577 136961 271625 136989
rect 271653 136961 271687 136989
rect 271715 136961 271749 136989
rect 271777 136961 271811 136989
rect 271839 136961 271887 136989
rect 271577 128175 271887 136961
rect 271577 128147 271625 128175
rect 271653 128147 271687 128175
rect 271715 128147 271749 128175
rect 271777 128147 271811 128175
rect 271839 128147 271887 128175
rect 271577 128113 271887 128147
rect 271577 128085 271625 128113
rect 271653 128085 271687 128113
rect 271715 128085 271749 128113
rect 271777 128085 271811 128113
rect 271839 128085 271887 128113
rect 271577 128051 271887 128085
rect 271577 128023 271625 128051
rect 271653 128023 271687 128051
rect 271715 128023 271749 128051
rect 271777 128023 271811 128051
rect 271839 128023 271887 128051
rect 271577 127989 271887 128023
rect 271577 127961 271625 127989
rect 271653 127961 271687 127989
rect 271715 127961 271749 127989
rect 271777 127961 271811 127989
rect 271839 127961 271887 127989
rect 271577 119175 271887 127961
rect 271577 119147 271625 119175
rect 271653 119147 271687 119175
rect 271715 119147 271749 119175
rect 271777 119147 271811 119175
rect 271839 119147 271887 119175
rect 271577 119113 271887 119147
rect 271577 119085 271625 119113
rect 271653 119085 271687 119113
rect 271715 119085 271749 119113
rect 271777 119085 271811 119113
rect 271839 119085 271887 119113
rect 271577 119051 271887 119085
rect 271577 119023 271625 119051
rect 271653 119023 271687 119051
rect 271715 119023 271749 119051
rect 271777 119023 271811 119051
rect 271839 119023 271887 119051
rect 271577 118989 271887 119023
rect 271577 118961 271625 118989
rect 271653 118961 271687 118989
rect 271715 118961 271749 118989
rect 271777 118961 271811 118989
rect 271839 118961 271887 118989
rect 271577 110175 271887 118961
rect 271577 110147 271625 110175
rect 271653 110147 271687 110175
rect 271715 110147 271749 110175
rect 271777 110147 271811 110175
rect 271839 110147 271887 110175
rect 271577 110113 271887 110147
rect 271577 110085 271625 110113
rect 271653 110085 271687 110113
rect 271715 110085 271749 110113
rect 271777 110085 271811 110113
rect 271839 110085 271887 110113
rect 271577 110051 271887 110085
rect 271577 110023 271625 110051
rect 271653 110023 271687 110051
rect 271715 110023 271749 110051
rect 271777 110023 271811 110051
rect 271839 110023 271887 110051
rect 271577 109989 271887 110023
rect 271577 109961 271625 109989
rect 271653 109961 271687 109989
rect 271715 109961 271749 109989
rect 271777 109961 271811 109989
rect 271839 109961 271887 109989
rect 271577 101175 271887 109961
rect 271577 101147 271625 101175
rect 271653 101147 271687 101175
rect 271715 101147 271749 101175
rect 271777 101147 271811 101175
rect 271839 101147 271887 101175
rect 271577 101113 271887 101147
rect 271577 101085 271625 101113
rect 271653 101085 271687 101113
rect 271715 101085 271749 101113
rect 271777 101085 271811 101113
rect 271839 101085 271887 101113
rect 271577 101051 271887 101085
rect 271577 101023 271625 101051
rect 271653 101023 271687 101051
rect 271715 101023 271749 101051
rect 271777 101023 271811 101051
rect 271839 101023 271887 101051
rect 271577 100989 271887 101023
rect 271577 100961 271625 100989
rect 271653 100961 271687 100989
rect 271715 100961 271749 100989
rect 271777 100961 271811 100989
rect 271839 100961 271887 100989
rect 271577 92175 271887 100961
rect 271577 92147 271625 92175
rect 271653 92147 271687 92175
rect 271715 92147 271749 92175
rect 271777 92147 271811 92175
rect 271839 92147 271887 92175
rect 271577 92113 271887 92147
rect 271577 92085 271625 92113
rect 271653 92085 271687 92113
rect 271715 92085 271749 92113
rect 271777 92085 271811 92113
rect 271839 92085 271887 92113
rect 271577 92051 271887 92085
rect 271577 92023 271625 92051
rect 271653 92023 271687 92051
rect 271715 92023 271749 92051
rect 271777 92023 271811 92051
rect 271839 92023 271887 92051
rect 271577 91989 271887 92023
rect 271577 91961 271625 91989
rect 271653 91961 271687 91989
rect 271715 91961 271749 91989
rect 271777 91961 271811 91989
rect 271839 91961 271887 91989
rect 271577 83175 271887 91961
rect 271577 83147 271625 83175
rect 271653 83147 271687 83175
rect 271715 83147 271749 83175
rect 271777 83147 271811 83175
rect 271839 83147 271887 83175
rect 271577 83113 271887 83147
rect 271577 83085 271625 83113
rect 271653 83085 271687 83113
rect 271715 83085 271749 83113
rect 271777 83085 271811 83113
rect 271839 83085 271887 83113
rect 271577 83051 271887 83085
rect 271577 83023 271625 83051
rect 271653 83023 271687 83051
rect 271715 83023 271749 83051
rect 271777 83023 271811 83051
rect 271839 83023 271887 83051
rect 271577 82989 271887 83023
rect 271577 82961 271625 82989
rect 271653 82961 271687 82989
rect 271715 82961 271749 82989
rect 271777 82961 271811 82989
rect 271839 82961 271887 82989
rect 271577 74175 271887 82961
rect 271577 74147 271625 74175
rect 271653 74147 271687 74175
rect 271715 74147 271749 74175
rect 271777 74147 271811 74175
rect 271839 74147 271887 74175
rect 271577 74113 271887 74147
rect 271577 74085 271625 74113
rect 271653 74085 271687 74113
rect 271715 74085 271749 74113
rect 271777 74085 271811 74113
rect 271839 74085 271887 74113
rect 271577 74051 271887 74085
rect 271577 74023 271625 74051
rect 271653 74023 271687 74051
rect 271715 74023 271749 74051
rect 271777 74023 271811 74051
rect 271839 74023 271887 74051
rect 271577 73989 271887 74023
rect 271577 73961 271625 73989
rect 271653 73961 271687 73989
rect 271715 73961 271749 73989
rect 271777 73961 271811 73989
rect 271839 73961 271887 73989
rect 271577 65175 271887 73961
rect 271577 65147 271625 65175
rect 271653 65147 271687 65175
rect 271715 65147 271749 65175
rect 271777 65147 271811 65175
rect 271839 65147 271887 65175
rect 271577 65113 271887 65147
rect 271577 65085 271625 65113
rect 271653 65085 271687 65113
rect 271715 65085 271749 65113
rect 271777 65085 271811 65113
rect 271839 65085 271887 65113
rect 271577 65051 271887 65085
rect 271577 65023 271625 65051
rect 271653 65023 271687 65051
rect 271715 65023 271749 65051
rect 271777 65023 271811 65051
rect 271839 65023 271887 65051
rect 271577 64989 271887 65023
rect 271577 64961 271625 64989
rect 271653 64961 271687 64989
rect 271715 64961 271749 64989
rect 271777 64961 271811 64989
rect 271839 64961 271887 64989
rect 271577 56175 271887 64961
rect 271577 56147 271625 56175
rect 271653 56147 271687 56175
rect 271715 56147 271749 56175
rect 271777 56147 271811 56175
rect 271839 56147 271887 56175
rect 271577 56113 271887 56147
rect 271577 56085 271625 56113
rect 271653 56085 271687 56113
rect 271715 56085 271749 56113
rect 271777 56085 271811 56113
rect 271839 56085 271887 56113
rect 271577 56051 271887 56085
rect 271577 56023 271625 56051
rect 271653 56023 271687 56051
rect 271715 56023 271749 56051
rect 271777 56023 271811 56051
rect 271839 56023 271887 56051
rect 271577 55989 271887 56023
rect 271577 55961 271625 55989
rect 271653 55961 271687 55989
rect 271715 55961 271749 55989
rect 271777 55961 271811 55989
rect 271839 55961 271887 55989
rect 271577 47175 271887 55961
rect 271577 47147 271625 47175
rect 271653 47147 271687 47175
rect 271715 47147 271749 47175
rect 271777 47147 271811 47175
rect 271839 47147 271887 47175
rect 271577 47113 271887 47147
rect 271577 47085 271625 47113
rect 271653 47085 271687 47113
rect 271715 47085 271749 47113
rect 271777 47085 271811 47113
rect 271839 47085 271887 47113
rect 271577 47051 271887 47085
rect 271577 47023 271625 47051
rect 271653 47023 271687 47051
rect 271715 47023 271749 47051
rect 271777 47023 271811 47051
rect 271839 47023 271887 47051
rect 271577 46989 271887 47023
rect 271577 46961 271625 46989
rect 271653 46961 271687 46989
rect 271715 46961 271749 46989
rect 271777 46961 271811 46989
rect 271839 46961 271887 46989
rect 271577 38175 271887 46961
rect 271577 38147 271625 38175
rect 271653 38147 271687 38175
rect 271715 38147 271749 38175
rect 271777 38147 271811 38175
rect 271839 38147 271887 38175
rect 271577 38113 271887 38147
rect 271577 38085 271625 38113
rect 271653 38085 271687 38113
rect 271715 38085 271749 38113
rect 271777 38085 271811 38113
rect 271839 38085 271887 38113
rect 271577 38051 271887 38085
rect 271577 38023 271625 38051
rect 271653 38023 271687 38051
rect 271715 38023 271749 38051
rect 271777 38023 271811 38051
rect 271839 38023 271887 38051
rect 271577 37989 271887 38023
rect 271577 37961 271625 37989
rect 271653 37961 271687 37989
rect 271715 37961 271749 37989
rect 271777 37961 271811 37989
rect 271839 37961 271887 37989
rect 271577 29175 271887 37961
rect 271577 29147 271625 29175
rect 271653 29147 271687 29175
rect 271715 29147 271749 29175
rect 271777 29147 271811 29175
rect 271839 29147 271887 29175
rect 271577 29113 271887 29147
rect 271577 29085 271625 29113
rect 271653 29085 271687 29113
rect 271715 29085 271749 29113
rect 271777 29085 271811 29113
rect 271839 29085 271887 29113
rect 271577 29051 271887 29085
rect 271577 29023 271625 29051
rect 271653 29023 271687 29051
rect 271715 29023 271749 29051
rect 271777 29023 271811 29051
rect 271839 29023 271887 29051
rect 271577 28989 271887 29023
rect 271577 28961 271625 28989
rect 271653 28961 271687 28989
rect 271715 28961 271749 28989
rect 271777 28961 271811 28989
rect 271839 28961 271887 28989
rect 271577 20175 271887 28961
rect 271577 20147 271625 20175
rect 271653 20147 271687 20175
rect 271715 20147 271749 20175
rect 271777 20147 271811 20175
rect 271839 20147 271887 20175
rect 271577 20113 271887 20147
rect 271577 20085 271625 20113
rect 271653 20085 271687 20113
rect 271715 20085 271749 20113
rect 271777 20085 271811 20113
rect 271839 20085 271887 20113
rect 271577 20051 271887 20085
rect 271577 20023 271625 20051
rect 271653 20023 271687 20051
rect 271715 20023 271749 20051
rect 271777 20023 271811 20051
rect 271839 20023 271887 20051
rect 271577 19989 271887 20023
rect 271577 19961 271625 19989
rect 271653 19961 271687 19989
rect 271715 19961 271749 19989
rect 271777 19961 271811 19989
rect 271839 19961 271887 19989
rect 271577 11175 271887 19961
rect 271577 11147 271625 11175
rect 271653 11147 271687 11175
rect 271715 11147 271749 11175
rect 271777 11147 271811 11175
rect 271839 11147 271887 11175
rect 271577 11113 271887 11147
rect 271577 11085 271625 11113
rect 271653 11085 271687 11113
rect 271715 11085 271749 11113
rect 271777 11085 271811 11113
rect 271839 11085 271887 11113
rect 271577 11051 271887 11085
rect 271577 11023 271625 11051
rect 271653 11023 271687 11051
rect 271715 11023 271749 11051
rect 271777 11023 271811 11051
rect 271839 11023 271887 11051
rect 271577 10989 271887 11023
rect 271577 10961 271625 10989
rect 271653 10961 271687 10989
rect 271715 10961 271749 10989
rect 271777 10961 271811 10989
rect 271839 10961 271887 10989
rect 271577 2175 271887 10961
rect 271577 2147 271625 2175
rect 271653 2147 271687 2175
rect 271715 2147 271749 2175
rect 271777 2147 271811 2175
rect 271839 2147 271887 2175
rect 271577 2113 271887 2147
rect 271577 2085 271625 2113
rect 271653 2085 271687 2113
rect 271715 2085 271749 2113
rect 271777 2085 271811 2113
rect 271839 2085 271887 2113
rect 271577 2051 271887 2085
rect 271577 2023 271625 2051
rect 271653 2023 271687 2051
rect 271715 2023 271749 2051
rect 271777 2023 271811 2051
rect 271839 2023 271887 2051
rect 271577 1989 271887 2023
rect 271577 1961 271625 1989
rect 271653 1961 271687 1989
rect 271715 1961 271749 1989
rect 271777 1961 271811 1989
rect 271839 1961 271887 1989
rect 271577 -80 271887 1961
rect 271577 -108 271625 -80
rect 271653 -108 271687 -80
rect 271715 -108 271749 -80
rect 271777 -108 271811 -80
rect 271839 -108 271887 -80
rect 271577 -142 271887 -108
rect 271577 -170 271625 -142
rect 271653 -170 271687 -142
rect 271715 -170 271749 -142
rect 271777 -170 271811 -142
rect 271839 -170 271887 -142
rect 271577 -204 271887 -170
rect 271577 -232 271625 -204
rect 271653 -232 271687 -204
rect 271715 -232 271749 -204
rect 271777 -232 271811 -204
rect 271839 -232 271887 -204
rect 271577 -266 271887 -232
rect 271577 -294 271625 -266
rect 271653 -294 271687 -266
rect 271715 -294 271749 -266
rect 271777 -294 271811 -266
rect 271839 -294 271887 -266
rect 271577 -822 271887 -294
rect 273437 299086 273747 299134
rect 273437 299058 273485 299086
rect 273513 299058 273547 299086
rect 273575 299058 273609 299086
rect 273637 299058 273671 299086
rect 273699 299058 273747 299086
rect 273437 299024 273747 299058
rect 273437 298996 273485 299024
rect 273513 298996 273547 299024
rect 273575 298996 273609 299024
rect 273637 298996 273671 299024
rect 273699 298996 273747 299024
rect 273437 298962 273747 298996
rect 273437 298934 273485 298962
rect 273513 298934 273547 298962
rect 273575 298934 273609 298962
rect 273637 298934 273671 298962
rect 273699 298934 273747 298962
rect 273437 298900 273747 298934
rect 273437 298872 273485 298900
rect 273513 298872 273547 298900
rect 273575 298872 273609 298900
rect 273637 298872 273671 298900
rect 273699 298872 273747 298900
rect 273437 293175 273747 298872
rect 273437 293147 273485 293175
rect 273513 293147 273547 293175
rect 273575 293147 273609 293175
rect 273637 293147 273671 293175
rect 273699 293147 273747 293175
rect 273437 293113 273747 293147
rect 273437 293085 273485 293113
rect 273513 293085 273547 293113
rect 273575 293085 273609 293113
rect 273637 293085 273671 293113
rect 273699 293085 273747 293113
rect 273437 293051 273747 293085
rect 273437 293023 273485 293051
rect 273513 293023 273547 293051
rect 273575 293023 273609 293051
rect 273637 293023 273671 293051
rect 273699 293023 273747 293051
rect 273437 292989 273747 293023
rect 273437 292961 273485 292989
rect 273513 292961 273547 292989
rect 273575 292961 273609 292989
rect 273637 292961 273671 292989
rect 273699 292961 273747 292989
rect 273437 284175 273747 292961
rect 273437 284147 273485 284175
rect 273513 284147 273547 284175
rect 273575 284147 273609 284175
rect 273637 284147 273671 284175
rect 273699 284147 273747 284175
rect 273437 284113 273747 284147
rect 273437 284085 273485 284113
rect 273513 284085 273547 284113
rect 273575 284085 273609 284113
rect 273637 284085 273671 284113
rect 273699 284085 273747 284113
rect 273437 284051 273747 284085
rect 273437 284023 273485 284051
rect 273513 284023 273547 284051
rect 273575 284023 273609 284051
rect 273637 284023 273671 284051
rect 273699 284023 273747 284051
rect 273437 283989 273747 284023
rect 273437 283961 273485 283989
rect 273513 283961 273547 283989
rect 273575 283961 273609 283989
rect 273637 283961 273671 283989
rect 273699 283961 273747 283989
rect 273437 275175 273747 283961
rect 273437 275147 273485 275175
rect 273513 275147 273547 275175
rect 273575 275147 273609 275175
rect 273637 275147 273671 275175
rect 273699 275147 273747 275175
rect 273437 275113 273747 275147
rect 273437 275085 273485 275113
rect 273513 275085 273547 275113
rect 273575 275085 273609 275113
rect 273637 275085 273671 275113
rect 273699 275085 273747 275113
rect 273437 275051 273747 275085
rect 273437 275023 273485 275051
rect 273513 275023 273547 275051
rect 273575 275023 273609 275051
rect 273637 275023 273671 275051
rect 273699 275023 273747 275051
rect 273437 274989 273747 275023
rect 273437 274961 273485 274989
rect 273513 274961 273547 274989
rect 273575 274961 273609 274989
rect 273637 274961 273671 274989
rect 273699 274961 273747 274989
rect 273437 266175 273747 274961
rect 273437 266147 273485 266175
rect 273513 266147 273547 266175
rect 273575 266147 273609 266175
rect 273637 266147 273671 266175
rect 273699 266147 273747 266175
rect 273437 266113 273747 266147
rect 273437 266085 273485 266113
rect 273513 266085 273547 266113
rect 273575 266085 273609 266113
rect 273637 266085 273671 266113
rect 273699 266085 273747 266113
rect 273437 266051 273747 266085
rect 273437 266023 273485 266051
rect 273513 266023 273547 266051
rect 273575 266023 273609 266051
rect 273637 266023 273671 266051
rect 273699 266023 273747 266051
rect 273437 265989 273747 266023
rect 273437 265961 273485 265989
rect 273513 265961 273547 265989
rect 273575 265961 273609 265989
rect 273637 265961 273671 265989
rect 273699 265961 273747 265989
rect 273437 257175 273747 265961
rect 273437 257147 273485 257175
rect 273513 257147 273547 257175
rect 273575 257147 273609 257175
rect 273637 257147 273671 257175
rect 273699 257147 273747 257175
rect 273437 257113 273747 257147
rect 273437 257085 273485 257113
rect 273513 257085 273547 257113
rect 273575 257085 273609 257113
rect 273637 257085 273671 257113
rect 273699 257085 273747 257113
rect 273437 257051 273747 257085
rect 273437 257023 273485 257051
rect 273513 257023 273547 257051
rect 273575 257023 273609 257051
rect 273637 257023 273671 257051
rect 273699 257023 273747 257051
rect 273437 256989 273747 257023
rect 273437 256961 273485 256989
rect 273513 256961 273547 256989
rect 273575 256961 273609 256989
rect 273637 256961 273671 256989
rect 273699 256961 273747 256989
rect 273437 248175 273747 256961
rect 273437 248147 273485 248175
rect 273513 248147 273547 248175
rect 273575 248147 273609 248175
rect 273637 248147 273671 248175
rect 273699 248147 273747 248175
rect 273437 248113 273747 248147
rect 273437 248085 273485 248113
rect 273513 248085 273547 248113
rect 273575 248085 273609 248113
rect 273637 248085 273671 248113
rect 273699 248085 273747 248113
rect 273437 248051 273747 248085
rect 273437 248023 273485 248051
rect 273513 248023 273547 248051
rect 273575 248023 273609 248051
rect 273637 248023 273671 248051
rect 273699 248023 273747 248051
rect 273437 247989 273747 248023
rect 273437 247961 273485 247989
rect 273513 247961 273547 247989
rect 273575 247961 273609 247989
rect 273637 247961 273671 247989
rect 273699 247961 273747 247989
rect 273437 239175 273747 247961
rect 273437 239147 273485 239175
rect 273513 239147 273547 239175
rect 273575 239147 273609 239175
rect 273637 239147 273671 239175
rect 273699 239147 273747 239175
rect 273437 239113 273747 239147
rect 273437 239085 273485 239113
rect 273513 239085 273547 239113
rect 273575 239085 273609 239113
rect 273637 239085 273671 239113
rect 273699 239085 273747 239113
rect 273437 239051 273747 239085
rect 273437 239023 273485 239051
rect 273513 239023 273547 239051
rect 273575 239023 273609 239051
rect 273637 239023 273671 239051
rect 273699 239023 273747 239051
rect 273437 238989 273747 239023
rect 273437 238961 273485 238989
rect 273513 238961 273547 238989
rect 273575 238961 273609 238989
rect 273637 238961 273671 238989
rect 273699 238961 273747 238989
rect 273437 230175 273747 238961
rect 273437 230147 273485 230175
rect 273513 230147 273547 230175
rect 273575 230147 273609 230175
rect 273637 230147 273671 230175
rect 273699 230147 273747 230175
rect 273437 230113 273747 230147
rect 273437 230085 273485 230113
rect 273513 230085 273547 230113
rect 273575 230085 273609 230113
rect 273637 230085 273671 230113
rect 273699 230085 273747 230113
rect 273437 230051 273747 230085
rect 273437 230023 273485 230051
rect 273513 230023 273547 230051
rect 273575 230023 273609 230051
rect 273637 230023 273671 230051
rect 273699 230023 273747 230051
rect 273437 229989 273747 230023
rect 273437 229961 273485 229989
rect 273513 229961 273547 229989
rect 273575 229961 273609 229989
rect 273637 229961 273671 229989
rect 273699 229961 273747 229989
rect 273437 221175 273747 229961
rect 273437 221147 273485 221175
rect 273513 221147 273547 221175
rect 273575 221147 273609 221175
rect 273637 221147 273671 221175
rect 273699 221147 273747 221175
rect 273437 221113 273747 221147
rect 273437 221085 273485 221113
rect 273513 221085 273547 221113
rect 273575 221085 273609 221113
rect 273637 221085 273671 221113
rect 273699 221085 273747 221113
rect 273437 221051 273747 221085
rect 273437 221023 273485 221051
rect 273513 221023 273547 221051
rect 273575 221023 273609 221051
rect 273637 221023 273671 221051
rect 273699 221023 273747 221051
rect 273437 220989 273747 221023
rect 273437 220961 273485 220989
rect 273513 220961 273547 220989
rect 273575 220961 273609 220989
rect 273637 220961 273671 220989
rect 273699 220961 273747 220989
rect 273437 212175 273747 220961
rect 273437 212147 273485 212175
rect 273513 212147 273547 212175
rect 273575 212147 273609 212175
rect 273637 212147 273671 212175
rect 273699 212147 273747 212175
rect 273437 212113 273747 212147
rect 273437 212085 273485 212113
rect 273513 212085 273547 212113
rect 273575 212085 273609 212113
rect 273637 212085 273671 212113
rect 273699 212085 273747 212113
rect 273437 212051 273747 212085
rect 273437 212023 273485 212051
rect 273513 212023 273547 212051
rect 273575 212023 273609 212051
rect 273637 212023 273671 212051
rect 273699 212023 273747 212051
rect 273437 211989 273747 212023
rect 273437 211961 273485 211989
rect 273513 211961 273547 211989
rect 273575 211961 273609 211989
rect 273637 211961 273671 211989
rect 273699 211961 273747 211989
rect 273437 203175 273747 211961
rect 273437 203147 273485 203175
rect 273513 203147 273547 203175
rect 273575 203147 273609 203175
rect 273637 203147 273671 203175
rect 273699 203147 273747 203175
rect 273437 203113 273747 203147
rect 273437 203085 273485 203113
rect 273513 203085 273547 203113
rect 273575 203085 273609 203113
rect 273637 203085 273671 203113
rect 273699 203085 273747 203113
rect 273437 203051 273747 203085
rect 273437 203023 273485 203051
rect 273513 203023 273547 203051
rect 273575 203023 273609 203051
rect 273637 203023 273671 203051
rect 273699 203023 273747 203051
rect 273437 202989 273747 203023
rect 273437 202961 273485 202989
rect 273513 202961 273547 202989
rect 273575 202961 273609 202989
rect 273637 202961 273671 202989
rect 273699 202961 273747 202989
rect 273437 194175 273747 202961
rect 273437 194147 273485 194175
rect 273513 194147 273547 194175
rect 273575 194147 273609 194175
rect 273637 194147 273671 194175
rect 273699 194147 273747 194175
rect 273437 194113 273747 194147
rect 273437 194085 273485 194113
rect 273513 194085 273547 194113
rect 273575 194085 273609 194113
rect 273637 194085 273671 194113
rect 273699 194085 273747 194113
rect 273437 194051 273747 194085
rect 273437 194023 273485 194051
rect 273513 194023 273547 194051
rect 273575 194023 273609 194051
rect 273637 194023 273671 194051
rect 273699 194023 273747 194051
rect 273437 193989 273747 194023
rect 273437 193961 273485 193989
rect 273513 193961 273547 193989
rect 273575 193961 273609 193989
rect 273637 193961 273671 193989
rect 273699 193961 273747 193989
rect 273437 185175 273747 193961
rect 273437 185147 273485 185175
rect 273513 185147 273547 185175
rect 273575 185147 273609 185175
rect 273637 185147 273671 185175
rect 273699 185147 273747 185175
rect 273437 185113 273747 185147
rect 273437 185085 273485 185113
rect 273513 185085 273547 185113
rect 273575 185085 273609 185113
rect 273637 185085 273671 185113
rect 273699 185085 273747 185113
rect 273437 185051 273747 185085
rect 273437 185023 273485 185051
rect 273513 185023 273547 185051
rect 273575 185023 273609 185051
rect 273637 185023 273671 185051
rect 273699 185023 273747 185051
rect 273437 184989 273747 185023
rect 273437 184961 273485 184989
rect 273513 184961 273547 184989
rect 273575 184961 273609 184989
rect 273637 184961 273671 184989
rect 273699 184961 273747 184989
rect 273437 176175 273747 184961
rect 273437 176147 273485 176175
rect 273513 176147 273547 176175
rect 273575 176147 273609 176175
rect 273637 176147 273671 176175
rect 273699 176147 273747 176175
rect 273437 176113 273747 176147
rect 273437 176085 273485 176113
rect 273513 176085 273547 176113
rect 273575 176085 273609 176113
rect 273637 176085 273671 176113
rect 273699 176085 273747 176113
rect 273437 176051 273747 176085
rect 273437 176023 273485 176051
rect 273513 176023 273547 176051
rect 273575 176023 273609 176051
rect 273637 176023 273671 176051
rect 273699 176023 273747 176051
rect 273437 175989 273747 176023
rect 273437 175961 273485 175989
rect 273513 175961 273547 175989
rect 273575 175961 273609 175989
rect 273637 175961 273671 175989
rect 273699 175961 273747 175989
rect 273437 167175 273747 175961
rect 273437 167147 273485 167175
rect 273513 167147 273547 167175
rect 273575 167147 273609 167175
rect 273637 167147 273671 167175
rect 273699 167147 273747 167175
rect 273437 167113 273747 167147
rect 273437 167085 273485 167113
rect 273513 167085 273547 167113
rect 273575 167085 273609 167113
rect 273637 167085 273671 167113
rect 273699 167085 273747 167113
rect 273437 167051 273747 167085
rect 273437 167023 273485 167051
rect 273513 167023 273547 167051
rect 273575 167023 273609 167051
rect 273637 167023 273671 167051
rect 273699 167023 273747 167051
rect 273437 166989 273747 167023
rect 273437 166961 273485 166989
rect 273513 166961 273547 166989
rect 273575 166961 273609 166989
rect 273637 166961 273671 166989
rect 273699 166961 273747 166989
rect 273437 158175 273747 166961
rect 273437 158147 273485 158175
rect 273513 158147 273547 158175
rect 273575 158147 273609 158175
rect 273637 158147 273671 158175
rect 273699 158147 273747 158175
rect 273437 158113 273747 158147
rect 273437 158085 273485 158113
rect 273513 158085 273547 158113
rect 273575 158085 273609 158113
rect 273637 158085 273671 158113
rect 273699 158085 273747 158113
rect 273437 158051 273747 158085
rect 273437 158023 273485 158051
rect 273513 158023 273547 158051
rect 273575 158023 273609 158051
rect 273637 158023 273671 158051
rect 273699 158023 273747 158051
rect 273437 157989 273747 158023
rect 273437 157961 273485 157989
rect 273513 157961 273547 157989
rect 273575 157961 273609 157989
rect 273637 157961 273671 157989
rect 273699 157961 273747 157989
rect 273437 149175 273747 157961
rect 273437 149147 273485 149175
rect 273513 149147 273547 149175
rect 273575 149147 273609 149175
rect 273637 149147 273671 149175
rect 273699 149147 273747 149175
rect 273437 149113 273747 149147
rect 273437 149085 273485 149113
rect 273513 149085 273547 149113
rect 273575 149085 273609 149113
rect 273637 149085 273671 149113
rect 273699 149085 273747 149113
rect 273437 149051 273747 149085
rect 273437 149023 273485 149051
rect 273513 149023 273547 149051
rect 273575 149023 273609 149051
rect 273637 149023 273671 149051
rect 273699 149023 273747 149051
rect 273437 148989 273747 149023
rect 273437 148961 273485 148989
rect 273513 148961 273547 148989
rect 273575 148961 273609 148989
rect 273637 148961 273671 148989
rect 273699 148961 273747 148989
rect 273437 140175 273747 148961
rect 273437 140147 273485 140175
rect 273513 140147 273547 140175
rect 273575 140147 273609 140175
rect 273637 140147 273671 140175
rect 273699 140147 273747 140175
rect 273437 140113 273747 140147
rect 273437 140085 273485 140113
rect 273513 140085 273547 140113
rect 273575 140085 273609 140113
rect 273637 140085 273671 140113
rect 273699 140085 273747 140113
rect 273437 140051 273747 140085
rect 273437 140023 273485 140051
rect 273513 140023 273547 140051
rect 273575 140023 273609 140051
rect 273637 140023 273671 140051
rect 273699 140023 273747 140051
rect 273437 139989 273747 140023
rect 273437 139961 273485 139989
rect 273513 139961 273547 139989
rect 273575 139961 273609 139989
rect 273637 139961 273671 139989
rect 273699 139961 273747 139989
rect 273437 131175 273747 139961
rect 273437 131147 273485 131175
rect 273513 131147 273547 131175
rect 273575 131147 273609 131175
rect 273637 131147 273671 131175
rect 273699 131147 273747 131175
rect 273437 131113 273747 131147
rect 273437 131085 273485 131113
rect 273513 131085 273547 131113
rect 273575 131085 273609 131113
rect 273637 131085 273671 131113
rect 273699 131085 273747 131113
rect 273437 131051 273747 131085
rect 273437 131023 273485 131051
rect 273513 131023 273547 131051
rect 273575 131023 273609 131051
rect 273637 131023 273671 131051
rect 273699 131023 273747 131051
rect 273437 130989 273747 131023
rect 273437 130961 273485 130989
rect 273513 130961 273547 130989
rect 273575 130961 273609 130989
rect 273637 130961 273671 130989
rect 273699 130961 273747 130989
rect 273437 122175 273747 130961
rect 273437 122147 273485 122175
rect 273513 122147 273547 122175
rect 273575 122147 273609 122175
rect 273637 122147 273671 122175
rect 273699 122147 273747 122175
rect 273437 122113 273747 122147
rect 273437 122085 273485 122113
rect 273513 122085 273547 122113
rect 273575 122085 273609 122113
rect 273637 122085 273671 122113
rect 273699 122085 273747 122113
rect 273437 122051 273747 122085
rect 273437 122023 273485 122051
rect 273513 122023 273547 122051
rect 273575 122023 273609 122051
rect 273637 122023 273671 122051
rect 273699 122023 273747 122051
rect 273437 121989 273747 122023
rect 273437 121961 273485 121989
rect 273513 121961 273547 121989
rect 273575 121961 273609 121989
rect 273637 121961 273671 121989
rect 273699 121961 273747 121989
rect 273437 113175 273747 121961
rect 273437 113147 273485 113175
rect 273513 113147 273547 113175
rect 273575 113147 273609 113175
rect 273637 113147 273671 113175
rect 273699 113147 273747 113175
rect 273437 113113 273747 113147
rect 273437 113085 273485 113113
rect 273513 113085 273547 113113
rect 273575 113085 273609 113113
rect 273637 113085 273671 113113
rect 273699 113085 273747 113113
rect 273437 113051 273747 113085
rect 273437 113023 273485 113051
rect 273513 113023 273547 113051
rect 273575 113023 273609 113051
rect 273637 113023 273671 113051
rect 273699 113023 273747 113051
rect 273437 112989 273747 113023
rect 273437 112961 273485 112989
rect 273513 112961 273547 112989
rect 273575 112961 273609 112989
rect 273637 112961 273671 112989
rect 273699 112961 273747 112989
rect 273437 104175 273747 112961
rect 273437 104147 273485 104175
rect 273513 104147 273547 104175
rect 273575 104147 273609 104175
rect 273637 104147 273671 104175
rect 273699 104147 273747 104175
rect 273437 104113 273747 104147
rect 273437 104085 273485 104113
rect 273513 104085 273547 104113
rect 273575 104085 273609 104113
rect 273637 104085 273671 104113
rect 273699 104085 273747 104113
rect 273437 104051 273747 104085
rect 273437 104023 273485 104051
rect 273513 104023 273547 104051
rect 273575 104023 273609 104051
rect 273637 104023 273671 104051
rect 273699 104023 273747 104051
rect 273437 103989 273747 104023
rect 273437 103961 273485 103989
rect 273513 103961 273547 103989
rect 273575 103961 273609 103989
rect 273637 103961 273671 103989
rect 273699 103961 273747 103989
rect 273437 95175 273747 103961
rect 273437 95147 273485 95175
rect 273513 95147 273547 95175
rect 273575 95147 273609 95175
rect 273637 95147 273671 95175
rect 273699 95147 273747 95175
rect 273437 95113 273747 95147
rect 273437 95085 273485 95113
rect 273513 95085 273547 95113
rect 273575 95085 273609 95113
rect 273637 95085 273671 95113
rect 273699 95085 273747 95113
rect 273437 95051 273747 95085
rect 273437 95023 273485 95051
rect 273513 95023 273547 95051
rect 273575 95023 273609 95051
rect 273637 95023 273671 95051
rect 273699 95023 273747 95051
rect 273437 94989 273747 95023
rect 273437 94961 273485 94989
rect 273513 94961 273547 94989
rect 273575 94961 273609 94989
rect 273637 94961 273671 94989
rect 273699 94961 273747 94989
rect 273437 86175 273747 94961
rect 273437 86147 273485 86175
rect 273513 86147 273547 86175
rect 273575 86147 273609 86175
rect 273637 86147 273671 86175
rect 273699 86147 273747 86175
rect 273437 86113 273747 86147
rect 273437 86085 273485 86113
rect 273513 86085 273547 86113
rect 273575 86085 273609 86113
rect 273637 86085 273671 86113
rect 273699 86085 273747 86113
rect 273437 86051 273747 86085
rect 273437 86023 273485 86051
rect 273513 86023 273547 86051
rect 273575 86023 273609 86051
rect 273637 86023 273671 86051
rect 273699 86023 273747 86051
rect 273437 85989 273747 86023
rect 273437 85961 273485 85989
rect 273513 85961 273547 85989
rect 273575 85961 273609 85989
rect 273637 85961 273671 85989
rect 273699 85961 273747 85989
rect 273437 77175 273747 85961
rect 273437 77147 273485 77175
rect 273513 77147 273547 77175
rect 273575 77147 273609 77175
rect 273637 77147 273671 77175
rect 273699 77147 273747 77175
rect 273437 77113 273747 77147
rect 273437 77085 273485 77113
rect 273513 77085 273547 77113
rect 273575 77085 273609 77113
rect 273637 77085 273671 77113
rect 273699 77085 273747 77113
rect 273437 77051 273747 77085
rect 273437 77023 273485 77051
rect 273513 77023 273547 77051
rect 273575 77023 273609 77051
rect 273637 77023 273671 77051
rect 273699 77023 273747 77051
rect 273437 76989 273747 77023
rect 273437 76961 273485 76989
rect 273513 76961 273547 76989
rect 273575 76961 273609 76989
rect 273637 76961 273671 76989
rect 273699 76961 273747 76989
rect 273437 68175 273747 76961
rect 273437 68147 273485 68175
rect 273513 68147 273547 68175
rect 273575 68147 273609 68175
rect 273637 68147 273671 68175
rect 273699 68147 273747 68175
rect 273437 68113 273747 68147
rect 273437 68085 273485 68113
rect 273513 68085 273547 68113
rect 273575 68085 273609 68113
rect 273637 68085 273671 68113
rect 273699 68085 273747 68113
rect 273437 68051 273747 68085
rect 273437 68023 273485 68051
rect 273513 68023 273547 68051
rect 273575 68023 273609 68051
rect 273637 68023 273671 68051
rect 273699 68023 273747 68051
rect 273437 67989 273747 68023
rect 273437 67961 273485 67989
rect 273513 67961 273547 67989
rect 273575 67961 273609 67989
rect 273637 67961 273671 67989
rect 273699 67961 273747 67989
rect 273437 59175 273747 67961
rect 273437 59147 273485 59175
rect 273513 59147 273547 59175
rect 273575 59147 273609 59175
rect 273637 59147 273671 59175
rect 273699 59147 273747 59175
rect 273437 59113 273747 59147
rect 273437 59085 273485 59113
rect 273513 59085 273547 59113
rect 273575 59085 273609 59113
rect 273637 59085 273671 59113
rect 273699 59085 273747 59113
rect 273437 59051 273747 59085
rect 273437 59023 273485 59051
rect 273513 59023 273547 59051
rect 273575 59023 273609 59051
rect 273637 59023 273671 59051
rect 273699 59023 273747 59051
rect 273437 58989 273747 59023
rect 273437 58961 273485 58989
rect 273513 58961 273547 58989
rect 273575 58961 273609 58989
rect 273637 58961 273671 58989
rect 273699 58961 273747 58989
rect 273437 50175 273747 58961
rect 273437 50147 273485 50175
rect 273513 50147 273547 50175
rect 273575 50147 273609 50175
rect 273637 50147 273671 50175
rect 273699 50147 273747 50175
rect 273437 50113 273747 50147
rect 273437 50085 273485 50113
rect 273513 50085 273547 50113
rect 273575 50085 273609 50113
rect 273637 50085 273671 50113
rect 273699 50085 273747 50113
rect 273437 50051 273747 50085
rect 273437 50023 273485 50051
rect 273513 50023 273547 50051
rect 273575 50023 273609 50051
rect 273637 50023 273671 50051
rect 273699 50023 273747 50051
rect 273437 49989 273747 50023
rect 273437 49961 273485 49989
rect 273513 49961 273547 49989
rect 273575 49961 273609 49989
rect 273637 49961 273671 49989
rect 273699 49961 273747 49989
rect 273437 41175 273747 49961
rect 273437 41147 273485 41175
rect 273513 41147 273547 41175
rect 273575 41147 273609 41175
rect 273637 41147 273671 41175
rect 273699 41147 273747 41175
rect 273437 41113 273747 41147
rect 273437 41085 273485 41113
rect 273513 41085 273547 41113
rect 273575 41085 273609 41113
rect 273637 41085 273671 41113
rect 273699 41085 273747 41113
rect 273437 41051 273747 41085
rect 273437 41023 273485 41051
rect 273513 41023 273547 41051
rect 273575 41023 273609 41051
rect 273637 41023 273671 41051
rect 273699 41023 273747 41051
rect 273437 40989 273747 41023
rect 273437 40961 273485 40989
rect 273513 40961 273547 40989
rect 273575 40961 273609 40989
rect 273637 40961 273671 40989
rect 273699 40961 273747 40989
rect 273437 32175 273747 40961
rect 273437 32147 273485 32175
rect 273513 32147 273547 32175
rect 273575 32147 273609 32175
rect 273637 32147 273671 32175
rect 273699 32147 273747 32175
rect 273437 32113 273747 32147
rect 273437 32085 273485 32113
rect 273513 32085 273547 32113
rect 273575 32085 273609 32113
rect 273637 32085 273671 32113
rect 273699 32085 273747 32113
rect 273437 32051 273747 32085
rect 273437 32023 273485 32051
rect 273513 32023 273547 32051
rect 273575 32023 273609 32051
rect 273637 32023 273671 32051
rect 273699 32023 273747 32051
rect 273437 31989 273747 32023
rect 273437 31961 273485 31989
rect 273513 31961 273547 31989
rect 273575 31961 273609 31989
rect 273637 31961 273671 31989
rect 273699 31961 273747 31989
rect 273437 23175 273747 31961
rect 273437 23147 273485 23175
rect 273513 23147 273547 23175
rect 273575 23147 273609 23175
rect 273637 23147 273671 23175
rect 273699 23147 273747 23175
rect 273437 23113 273747 23147
rect 273437 23085 273485 23113
rect 273513 23085 273547 23113
rect 273575 23085 273609 23113
rect 273637 23085 273671 23113
rect 273699 23085 273747 23113
rect 273437 23051 273747 23085
rect 273437 23023 273485 23051
rect 273513 23023 273547 23051
rect 273575 23023 273609 23051
rect 273637 23023 273671 23051
rect 273699 23023 273747 23051
rect 273437 22989 273747 23023
rect 273437 22961 273485 22989
rect 273513 22961 273547 22989
rect 273575 22961 273609 22989
rect 273637 22961 273671 22989
rect 273699 22961 273747 22989
rect 273437 14175 273747 22961
rect 273437 14147 273485 14175
rect 273513 14147 273547 14175
rect 273575 14147 273609 14175
rect 273637 14147 273671 14175
rect 273699 14147 273747 14175
rect 273437 14113 273747 14147
rect 273437 14085 273485 14113
rect 273513 14085 273547 14113
rect 273575 14085 273609 14113
rect 273637 14085 273671 14113
rect 273699 14085 273747 14113
rect 273437 14051 273747 14085
rect 273437 14023 273485 14051
rect 273513 14023 273547 14051
rect 273575 14023 273609 14051
rect 273637 14023 273671 14051
rect 273699 14023 273747 14051
rect 273437 13989 273747 14023
rect 273437 13961 273485 13989
rect 273513 13961 273547 13989
rect 273575 13961 273609 13989
rect 273637 13961 273671 13989
rect 273699 13961 273747 13989
rect 273437 5175 273747 13961
rect 273437 5147 273485 5175
rect 273513 5147 273547 5175
rect 273575 5147 273609 5175
rect 273637 5147 273671 5175
rect 273699 5147 273747 5175
rect 273437 5113 273747 5147
rect 273437 5085 273485 5113
rect 273513 5085 273547 5113
rect 273575 5085 273609 5113
rect 273637 5085 273671 5113
rect 273699 5085 273747 5113
rect 273437 5051 273747 5085
rect 273437 5023 273485 5051
rect 273513 5023 273547 5051
rect 273575 5023 273609 5051
rect 273637 5023 273671 5051
rect 273699 5023 273747 5051
rect 273437 4989 273747 5023
rect 273437 4961 273485 4989
rect 273513 4961 273547 4989
rect 273575 4961 273609 4989
rect 273637 4961 273671 4989
rect 273699 4961 273747 4989
rect 273437 -560 273747 4961
rect 273437 -588 273485 -560
rect 273513 -588 273547 -560
rect 273575 -588 273609 -560
rect 273637 -588 273671 -560
rect 273699 -588 273747 -560
rect 273437 -622 273747 -588
rect 273437 -650 273485 -622
rect 273513 -650 273547 -622
rect 273575 -650 273609 -622
rect 273637 -650 273671 -622
rect 273699 -650 273747 -622
rect 273437 -684 273747 -650
rect 273437 -712 273485 -684
rect 273513 -712 273547 -684
rect 273575 -712 273609 -684
rect 273637 -712 273671 -684
rect 273699 -712 273747 -684
rect 273437 -746 273747 -712
rect 273437 -774 273485 -746
rect 273513 -774 273547 -746
rect 273575 -774 273609 -746
rect 273637 -774 273671 -746
rect 273699 -774 273747 -746
rect 273437 -822 273747 -774
rect 280577 298606 280887 299134
rect 280577 298578 280625 298606
rect 280653 298578 280687 298606
rect 280715 298578 280749 298606
rect 280777 298578 280811 298606
rect 280839 298578 280887 298606
rect 280577 298544 280887 298578
rect 280577 298516 280625 298544
rect 280653 298516 280687 298544
rect 280715 298516 280749 298544
rect 280777 298516 280811 298544
rect 280839 298516 280887 298544
rect 280577 298482 280887 298516
rect 280577 298454 280625 298482
rect 280653 298454 280687 298482
rect 280715 298454 280749 298482
rect 280777 298454 280811 298482
rect 280839 298454 280887 298482
rect 280577 298420 280887 298454
rect 280577 298392 280625 298420
rect 280653 298392 280687 298420
rect 280715 298392 280749 298420
rect 280777 298392 280811 298420
rect 280839 298392 280887 298420
rect 280577 290175 280887 298392
rect 280577 290147 280625 290175
rect 280653 290147 280687 290175
rect 280715 290147 280749 290175
rect 280777 290147 280811 290175
rect 280839 290147 280887 290175
rect 280577 290113 280887 290147
rect 280577 290085 280625 290113
rect 280653 290085 280687 290113
rect 280715 290085 280749 290113
rect 280777 290085 280811 290113
rect 280839 290085 280887 290113
rect 280577 290051 280887 290085
rect 280577 290023 280625 290051
rect 280653 290023 280687 290051
rect 280715 290023 280749 290051
rect 280777 290023 280811 290051
rect 280839 290023 280887 290051
rect 280577 289989 280887 290023
rect 280577 289961 280625 289989
rect 280653 289961 280687 289989
rect 280715 289961 280749 289989
rect 280777 289961 280811 289989
rect 280839 289961 280887 289989
rect 280577 281175 280887 289961
rect 280577 281147 280625 281175
rect 280653 281147 280687 281175
rect 280715 281147 280749 281175
rect 280777 281147 280811 281175
rect 280839 281147 280887 281175
rect 280577 281113 280887 281147
rect 280577 281085 280625 281113
rect 280653 281085 280687 281113
rect 280715 281085 280749 281113
rect 280777 281085 280811 281113
rect 280839 281085 280887 281113
rect 280577 281051 280887 281085
rect 280577 281023 280625 281051
rect 280653 281023 280687 281051
rect 280715 281023 280749 281051
rect 280777 281023 280811 281051
rect 280839 281023 280887 281051
rect 280577 280989 280887 281023
rect 280577 280961 280625 280989
rect 280653 280961 280687 280989
rect 280715 280961 280749 280989
rect 280777 280961 280811 280989
rect 280839 280961 280887 280989
rect 280577 272175 280887 280961
rect 280577 272147 280625 272175
rect 280653 272147 280687 272175
rect 280715 272147 280749 272175
rect 280777 272147 280811 272175
rect 280839 272147 280887 272175
rect 280577 272113 280887 272147
rect 280577 272085 280625 272113
rect 280653 272085 280687 272113
rect 280715 272085 280749 272113
rect 280777 272085 280811 272113
rect 280839 272085 280887 272113
rect 280577 272051 280887 272085
rect 280577 272023 280625 272051
rect 280653 272023 280687 272051
rect 280715 272023 280749 272051
rect 280777 272023 280811 272051
rect 280839 272023 280887 272051
rect 280577 271989 280887 272023
rect 280577 271961 280625 271989
rect 280653 271961 280687 271989
rect 280715 271961 280749 271989
rect 280777 271961 280811 271989
rect 280839 271961 280887 271989
rect 280577 263175 280887 271961
rect 280577 263147 280625 263175
rect 280653 263147 280687 263175
rect 280715 263147 280749 263175
rect 280777 263147 280811 263175
rect 280839 263147 280887 263175
rect 280577 263113 280887 263147
rect 280577 263085 280625 263113
rect 280653 263085 280687 263113
rect 280715 263085 280749 263113
rect 280777 263085 280811 263113
rect 280839 263085 280887 263113
rect 280577 263051 280887 263085
rect 280577 263023 280625 263051
rect 280653 263023 280687 263051
rect 280715 263023 280749 263051
rect 280777 263023 280811 263051
rect 280839 263023 280887 263051
rect 280577 262989 280887 263023
rect 280577 262961 280625 262989
rect 280653 262961 280687 262989
rect 280715 262961 280749 262989
rect 280777 262961 280811 262989
rect 280839 262961 280887 262989
rect 280577 254175 280887 262961
rect 280577 254147 280625 254175
rect 280653 254147 280687 254175
rect 280715 254147 280749 254175
rect 280777 254147 280811 254175
rect 280839 254147 280887 254175
rect 280577 254113 280887 254147
rect 280577 254085 280625 254113
rect 280653 254085 280687 254113
rect 280715 254085 280749 254113
rect 280777 254085 280811 254113
rect 280839 254085 280887 254113
rect 280577 254051 280887 254085
rect 280577 254023 280625 254051
rect 280653 254023 280687 254051
rect 280715 254023 280749 254051
rect 280777 254023 280811 254051
rect 280839 254023 280887 254051
rect 280577 253989 280887 254023
rect 280577 253961 280625 253989
rect 280653 253961 280687 253989
rect 280715 253961 280749 253989
rect 280777 253961 280811 253989
rect 280839 253961 280887 253989
rect 280577 245175 280887 253961
rect 280577 245147 280625 245175
rect 280653 245147 280687 245175
rect 280715 245147 280749 245175
rect 280777 245147 280811 245175
rect 280839 245147 280887 245175
rect 280577 245113 280887 245147
rect 280577 245085 280625 245113
rect 280653 245085 280687 245113
rect 280715 245085 280749 245113
rect 280777 245085 280811 245113
rect 280839 245085 280887 245113
rect 280577 245051 280887 245085
rect 280577 245023 280625 245051
rect 280653 245023 280687 245051
rect 280715 245023 280749 245051
rect 280777 245023 280811 245051
rect 280839 245023 280887 245051
rect 280577 244989 280887 245023
rect 280577 244961 280625 244989
rect 280653 244961 280687 244989
rect 280715 244961 280749 244989
rect 280777 244961 280811 244989
rect 280839 244961 280887 244989
rect 280577 236175 280887 244961
rect 280577 236147 280625 236175
rect 280653 236147 280687 236175
rect 280715 236147 280749 236175
rect 280777 236147 280811 236175
rect 280839 236147 280887 236175
rect 280577 236113 280887 236147
rect 280577 236085 280625 236113
rect 280653 236085 280687 236113
rect 280715 236085 280749 236113
rect 280777 236085 280811 236113
rect 280839 236085 280887 236113
rect 280577 236051 280887 236085
rect 280577 236023 280625 236051
rect 280653 236023 280687 236051
rect 280715 236023 280749 236051
rect 280777 236023 280811 236051
rect 280839 236023 280887 236051
rect 280577 235989 280887 236023
rect 280577 235961 280625 235989
rect 280653 235961 280687 235989
rect 280715 235961 280749 235989
rect 280777 235961 280811 235989
rect 280839 235961 280887 235989
rect 280577 227175 280887 235961
rect 280577 227147 280625 227175
rect 280653 227147 280687 227175
rect 280715 227147 280749 227175
rect 280777 227147 280811 227175
rect 280839 227147 280887 227175
rect 280577 227113 280887 227147
rect 280577 227085 280625 227113
rect 280653 227085 280687 227113
rect 280715 227085 280749 227113
rect 280777 227085 280811 227113
rect 280839 227085 280887 227113
rect 280577 227051 280887 227085
rect 280577 227023 280625 227051
rect 280653 227023 280687 227051
rect 280715 227023 280749 227051
rect 280777 227023 280811 227051
rect 280839 227023 280887 227051
rect 280577 226989 280887 227023
rect 280577 226961 280625 226989
rect 280653 226961 280687 226989
rect 280715 226961 280749 226989
rect 280777 226961 280811 226989
rect 280839 226961 280887 226989
rect 280577 218175 280887 226961
rect 280577 218147 280625 218175
rect 280653 218147 280687 218175
rect 280715 218147 280749 218175
rect 280777 218147 280811 218175
rect 280839 218147 280887 218175
rect 280577 218113 280887 218147
rect 280577 218085 280625 218113
rect 280653 218085 280687 218113
rect 280715 218085 280749 218113
rect 280777 218085 280811 218113
rect 280839 218085 280887 218113
rect 280577 218051 280887 218085
rect 280577 218023 280625 218051
rect 280653 218023 280687 218051
rect 280715 218023 280749 218051
rect 280777 218023 280811 218051
rect 280839 218023 280887 218051
rect 280577 217989 280887 218023
rect 280577 217961 280625 217989
rect 280653 217961 280687 217989
rect 280715 217961 280749 217989
rect 280777 217961 280811 217989
rect 280839 217961 280887 217989
rect 280577 209175 280887 217961
rect 280577 209147 280625 209175
rect 280653 209147 280687 209175
rect 280715 209147 280749 209175
rect 280777 209147 280811 209175
rect 280839 209147 280887 209175
rect 280577 209113 280887 209147
rect 280577 209085 280625 209113
rect 280653 209085 280687 209113
rect 280715 209085 280749 209113
rect 280777 209085 280811 209113
rect 280839 209085 280887 209113
rect 280577 209051 280887 209085
rect 280577 209023 280625 209051
rect 280653 209023 280687 209051
rect 280715 209023 280749 209051
rect 280777 209023 280811 209051
rect 280839 209023 280887 209051
rect 280577 208989 280887 209023
rect 280577 208961 280625 208989
rect 280653 208961 280687 208989
rect 280715 208961 280749 208989
rect 280777 208961 280811 208989
rect 280839 208961 280887 208989
rect 280577 200175 280887 208961
rect 280577 200147 280625 200175
rect 280653 200147 280687 200175
rect 280715 200147 280749 200175
rect 280777 200147 280811 200175
rect 280839 200147 280887 200175
rect 280577 200113 280887 200147
rect 280577 200085 280625 200113
rect 280653 200085 280687 200113
rect 280715 200085 280749 200113
rect 280777 200085 280811 200113
rect 280839 200085 280887 200113
rect 280577 200051 280887 200085
rect 280577 200023 280625 200051
rect 280653 200023 280687 200051
rect 280715 200023 280749 200051
rect 280777 200023 280811 200051
rect 280839 200023 280887 200051
rect 280577 199989 280887 200023
rect 280577 199961 280625 199989
rect 280653 199961 280687 199989
rect 280715 199961 280749 199989
rect 280777 199961 280811 199989
rect 280839 199961 280887 199989
rect 280577 191175 280887 199961
rect 280577 191147 280625 191175
rect 280653 191147 280687 191175
rect 280715 191147 280749 191175
rect 280777 191147 280811 191175
rect 280839 191147 280887 191175
rect 280577 191113 280887 191147
rect 280577 191085 280625 191113
rect 280653 191085 280687 191113
rect 280715 191085 280749 191113
rect 280777 191085 280811 191113
rect 280839 191085 280887 191113
rect 280577 191051 280887 191085
rect 280577 191023 280625 191051
rect 280653 191023 280687 191051
rect 280715 191023 280749 191051
rect 280777 191023 280811 191051
rect 280839 191023 280887 191051
rect 280577 190989 280887 191023
rect 280577 190961 280625 190989
rect 280653 190961 280687 190989
rect 280715 190961 280749 190989
rect 280777 190961 280811 190989
rect 280839 190961 280887 190989
rect 280577 182175 280887 190961
rect 280577 182147 280625 182175
rect 280653 182147 280687 182175
rect 280715 182147 280749 182175
rect 280777 182147 280811 182175
rect 280839 182147 280887 182175
rect 280577 182113 280887 182147
rect 280577 182085 280625 182113
rect 280653 182085 280687 182113
rect 280715 182085 280749 182113
rect 280777 182085 280811 182113
rect 280839 182085 280887 182113
rect 280577 182051 280887 182085
rect 280577 182023 280625 182051
rect 280653 182023 280687 182051
rect 280715 182023 280749 182051
rect 280777 182023 280811 182051
rect 280839 182023 280887 182051
rect 280577 181989 280887 182023
rect 280577 181961 280625 181989
rect 280653 181961 280687 181989
rect 280715 181961 280749 181989
rect 280777 181961 280811 181989
rect 280839 181961 280887 181989
rect 280577 173175 280887 181961
rect 280577 173147 280625 173175
rect 280653 173147 280687 173175
rect 280715 173147 280749 173175
rect 280777 173147 280811 173175
rect 280839 173147 280887 173175
rect 280577 173113 280887 173147
rect 280577 173085 280625 173113
rect 280653 173085 280687 173113
rect 280715 173085 280749 173113
rect 280777 173085 280811 173113
rect 280839 173085 280887 173113
rect 280577 173051 280887 173085
rect 280577 173023 280625 173051
rect 280653 173023 280687 173051
rect 280715 173023 280749 173051
rect 280777 173023 280811 173051
rect 280839 173023 280887 173051
rect 280577 172989 280887 173023
rect 280577 172961 280625 172989
rect 280653 172961 280687 172989
rect 280715 172961 280749 172989
rect 280777 172961 280811 172989
rect 280839 172961 280887 172989
rect 280577 164175 280887 172961
rect 280577 164147 280625 164175
rect 280653 164147 280687 164175
rect 280715 164147 280749 164175
rect 280777 164147 280811 164175
rect 280839 164147 280887 164175
rect 280577 164113 280887 164147
rect 280577 164085 280625 164113
rect 280653 164085 280687 164113
rect 280715 164085 280749 164113
rect 280777 164085 280811 164113
rect 280839 164085 280887 164113
rect 280577 164051 280887 164085
rect 280577 164023 280625 164051
rect 280653 164023 280687 164051
rect 280715 164023 280749 164051
rect 280777 164023 280811 164051
rect 280839 164023 280887 164051
rect 280577 163989 280887 164023
rect 280577 163961 280625 163989
rect 280653 163961 280687 163989
rect 280715 163961 280749 163989
rect 280777 163961 280811 163989
rect 280839 163961 280887 163989
rect 280577 155175 280887 163961
rect 280577 155147 280625 155175
rect 280653 155147 280687 155175
rect 280715 155147 280749 155175
rect 280777 155147 280811 155175
rect 280839 155147 280887 155175
rect 280577 155113 280887 155147
rect 280577 155085 280625 155113
rect 280653 155085 280687 155113
rect 280715 155085 280749 155113
rect 280777 155085 280811 155113
rect 280839 155085 280887 155113
rect 280577 155051 280887 155085
rect 280577 155023 280625 155051
rect 280653 155023 280687 155051
rect 280715 155023 280749 155051
rect 280777 155023 280811 155051
rect 280839 155023 280887 155051
rect 280577 154989 280887 155023
rect 280577 154961 280625 154989
rect 280653 154961 280687 154989
rect 280715 154961 280749 154989
rect 280777 154961 280811 154989
rect 280839 154961 280887 154989
rect 280577 146175 280887 154961
rect 280577 146147 280625 146175
rect 280653 146147 280687 146175
rect 280715 146147 280749 146175
rect 280777 146147 280811 146175
rect 280839 146147 280887 146175
rect 280577 146113 280887 146147
rect 280577 146085 280625 146113
rect 280653 146085 280687 146113
rect 280715 146085 280749 146113
rect 280777 146085 280811 146113
rect 280839 146085 280887 146113
rect 280577 146051 280887 146085
rect 280577 146023 280625 146051
rect 280653 146023 280687 146051
rect 280715 146023 280749 146051
rect 280777 146023 280811 146051
rect 280839 146023 280887 146051
rect 280577 145989 280887 146023
rect 280577 145961 280625 145989
rect 280653 145961 280687 145989
rect 280715 145961 280749 145989
rect 280777 145961 280811 145989
rect 280839 145961 280887 145989
rect 280577 137175 280887 145961
rect 280577 137147 280625 137175
rect 280653 137147 280687 137175
rect 280715 137147 280749 137175
rect 280777 137147 280811 137175
rect 280839 137147 280887 137175
rect 280577 137113 280887 137147
rect 280577 137085 280625 137113
rect 280653 137085 280687 137113
rect 280715 137085 280749 137113
rect 280777 137085 280811 137113
rect 280839 137085 280887 137113
rect 280577 137051 280887 137085
rect 280577 137023 280625 137051
rect 280653 137023 280687 137051
rect 280715 137023 280749 137051
rect 280777 137023 280811 137051
rect 280839 137023 280887 137051
rect 280577 136989 280887 137023
rect 280577 136961 280625 136989
rect 280653 136961 280687 136989
rect 280715 136961 280749 136989
rect 280777 136961 280811 136989
rect 280839 136961 280887 136989
rect 280577 128175 280887 136961
rect 280577 128147 280625 128175
rect 280653 128147 280687 128175
rect 280715 128147 280749 128175
rect 280777 128147 280811 128175
rect 280839 128147 280887 128175
rect 280577 128113 280887 128147
rect 280577 128085 280625 128113
rect 280653 128085 280687 128113
rect 280715 128085 280749 128113
rect 280777 128085 280811 128113
rect 280839 128085 280887 128113
rect 280577 128051 280887 128085
rect 280577 128023 280625 128051
rect 280653 128023 280687 128051
rect 280715 128023 280749 128051
rect 280777 128023 280811 128051
rect 280839 128023 280887 128051
rect 280577 127989 280887 128023
rect 280577 127961 280625 127989
rect 280653 127961 280687 127989
rect 280715 127961 280749 127989
rect 280777 127961 280811 127989
rect 280839 127961 280887 127989
rect 280577 119175 280887 127961
rect 280577 119147 280625 119175
rect 280653 119147 280687 119175
rect 280715 119147 280749 119175
rect 280777 119147 280811 119175
rect 280839 119147 280887 119175
rect 280577 119113 280887 119147
rect 280577 119085 280625 119113
rect 280653 119085 280687 119113
rect 280715 119085 280749 119113
rect 280777 119085 280811 119113
rect 280839 119085 280887 119113
rect 280577 119051 280887 119085
rect 280577 119023 280625 119051
rect 280653 119023 280687 119051
rect 280715 119023 280749 119051
rect 280777 119023 280811 119051
rect 280839 119023 280887 119051
rect 280577 118989 280887 119023
rect 280577 118961 280625 118989
rect 280653 118961 280687 118989
rect 280715 118961 280749 118989
rect 280777 118961 280811 118989
rect 280839 118961 280887 118989
rect 280577 110175 280887 118961
rect 280577 110147 280625 110175
rect 280653 110147 280687 110175
rect 280715 110147 280749 110175
rect 280777 110147 280811 110175
rect 280839 110147 280887 110175
rect 280577 110113 280887 110147
rect 280577 110085 280625 110113
rect 280653 110085 280687 110113
rect 280715 110085 280749 110113
rect 280777 110085 280811 110113
rect 280839 110085 280887 110113
rect 280577 110051 280887 110085
rect 280577 110023 280625 110051
rect 280653 110023 280687 110051
rect 280715 110023 280749 110051
rect 280777 110023 280811 110051
rect 280839 110023 280887 110051
rect 280577 109989 280887 110023
rect 280577 109961 280625 109989
rect 280653 109961 280687 109989
rect 280715 109961 280749 109989
rect 280777 109961 280811 109989
rect 280839 109961 280887 109989
rect 280577 101175 280887 109961
rect 280577 101147 280625 101175
rect 280653 101147 280687 101175
rect 280715 101147 280749 101175
rect 280777 101147 280811 101175
rect 280839 101147 280887 101175
rect 280577 101113 280887 101147
rect 280577 101085 280625 101113
rect 280653 101085 280687 101113
rect 280715 101085 280749 101113
rect 280777 101085 280811 101113
rect 280839 101085 280887 101113
rect 280577 101051 280887 101085
rect 280577 101023 280625 101051
rect 280653 101023 280687 101051
rect 280715 101023 280749 101051
rect 280777 101023 280811 101051
rect 280839 101023 280887 101051
rect 280577 100989 280887 101023
rect 280577 100961 280625 100989
rect 280653 100961 280687 100989
rect 280715 100961 280749 100989
rect 280777 100961 280811 100989
rect 280839 100961 280887 100989
rect 280577 92175 280887 100961
rect 280577 92147 280625 92175
rect 280653 92147 280687 92175
rect 280715 92147 280749 92175
rect 280777 92147 280811 92175
rect 280839 92147 280887 92175
rect 280577 92113 280887 92147
rect 280577 92085 280625 92113
rect 280653 92085 280687 92113
rect 280715 92085 280749 92113
rect 280777 92085 280811 92113
rect 280839 92085 280887 92113
rect 280577 92051 280887 92085
rect 280577 92023 280625 92051
rect 280653 92023 280687 92051
rect 280715 92023 280749 92051
rect 280777 92023 280811 92051
rect 280839 92023 280887 92051
rect 280577 91989 280887 92023
rect 280577 91961 280625 91989
rect 280653 91961 280687 91989
rect 280715 91961 280749 91989
rect 280777 91961 280811 91989
rect 280839 91961 280887 91989
rect 280577 83175 280887 91961
rect 280577 83147 280625 83175
rect 280653 83147 280687 83175
rect 280715 83147 280749 83175
rect 280777 83147 280811 83175
rect 280839 83147 280887 83175
rect 280577 83113 280887 83147
rect 280577 83085 280625 83113
rect 280653 83085 280687 83113
rect 280715 83085 280749 83113
rect 280777 83085 280811 83113
rect 280839 83085 280887 83113
rect 280577 83051 280887 83085
rect 280577 83023 280625 83051
rect 280653 83023 280687 83051
rect 280715 83023 280749 83051
rect 280777 83023 280811 83051
rect 280839 83023 280887 83051
rect 280577 82989 280887 83023
rect 280577 82961 280625 82989
rect 280653 82961 280687 82989
rect 280715 82961 280749 82989
rect 280777 82961 280811 82989
rect 280839 82961 280887 82989
rect 280577 74175 280887 82961
rect 280577 74147 280625 74175
rect 280653 74147 280687 74175
rect 280715 74147 280749 74175
rect 280777 74147 280811 74175
rect 280839 74147 280887 74175
rect 280577 74113 280887 74147
rect 280577 74085 280625 74113
rect 280653 74085 280687 74113
rect 280715 74085 280749 74113
rect 280777 74085 280811 74113
rect 280839 74085 280887 74113
rect 280577 74051 280887 74085
rect 280577 74023 280625 74051
rect 280653 74023 280687 74051
rect 280715 74023 280749 74051
rect 280777 74023 280811 74051
rect 280839 74023 280887 74051
rect 280577 73989 280887 74023
rect 280577 73961 280625 73989
rect 280653 73961 280687 73989
rect 280715 73961 280749 73989
rect 280777 73961 280811 73989
rect 280839 73961 280887 73989
rect 280577 65175 280887 73961
rect 280577 65147 280625 65175
rect 280653 65147 280687 65175
rect 280715 65147 280749 65175
rect 280777 65147 280811 65175
rect 280839 65147 280887 65175
rect 280577 65113 280887 65147
rect 280577 65085 280625 65113
rect 280653 65085 280687 65113
rect 280715 65085 280749 65113
rect 280777 65085 280811 65113
rect 280839 65085 280887 65113
rect 280577 65051 280887 65085
rect 280577 65023 280625 65051
rect 280653 65023 280687 65051
rect 280715 65023 280749 65051
rect 280777 65023 280811 65051
rect 280839 65023 280887 65051
rect 280577 64989 280887 65023
rect 280577 64961 280625 64989
rect 280653 64961 280687 64989
rect 280715 64961 280749 64989
rect 280777 64961 280811 64989
rect 280839 64961 280887 64989
rect 280577 56175 280887 64961
rect 280577 56147 280625 56175
rect 280653 56147 280687 56175
rect 280715 56147 280749 56175
rect 280777 56147 280811 56175
rect 280839 56147 280887 56175
rect 280577 56113 280887 56147
rect 280577 56085 280625 56113
rect 280653 56085 280687 56113
rect 280715 56085 280749 56113
rect 280777 56085 280811 56113
rect 280839 56085 280887 56113
rect 280577 56051 280887 56085
rect 280577 56023 280625 56051
rect 280653 56023 280687 56051
rect 280715 56023 280749 56051
rect 280777 56023 280811 56051
rect 280839 56023 280887 56051
rect 280577 55989 280887 56023
rect 280577 55961 280625 55989
rect 280653 55961 280687 55989
rect 280715 55961 280749 55989
rect 280777 55961 280811 55989
rect 280839 55961 280887 55989
rect 280577 47175 280887 55961
rect 280577 47147 280625 47175
rect 280653 47147 280687 47175
rect 280715 47147 280749 47175
rect 280777 47147 280811 47175
rect 280839 47147 280887 47175
rect 280577 47113 280887 47147
rect 280577 47085 280625 47113
rect 280653 47085 280687 47113
rect 280715 47085 280749 47113
rect 280777 47085 280811 47113
rect 280839 47085 280887 47113
rect 280577 47051 280887 47085
rect 280577 47023 280625 47051
rect 280653 47023 280687 47051
rect 280715 47023 280749 47051
rect 280777 47023 280811 47051
rect 280839 47023 280887 47051
rect 280577 46989 280887 47023
rect 280577 46961 280625 46989
rect 280653 46961 280687 46989
rect 280715 46961 280749 46989
rect 280777 46961 280811 46989
rect 280839 46961 280887 46989
rect 280577 38175 280887 46961
rect 280577 38147 280625 38175
rect 280653 38147 280687 38175
rect 280715 38147 280749 38175
rect 280777 38147 280811 38175
rect 280839 38147 280887 38175
rect 280577 38113 280887 38147
rect 280577 38085 280625 38113
rect 280653 38085 280687 38113
rect 280715 38085 280749 38113
rect 280777 38085 280811 38113
rect 280839 38085 280887 38113
rect 280577 38051 280887 38085
rect 280577 38023 280625 38051
rect 280653 38023 280687 38051
rect 280715 38023 280749 38051
rect 280777 38023 280811 38051
rect 280839 38023 280887 38051
rect 280577 37989 280887 38023
rect 280577 37961 280625 37989
rect 280653 37961 280687 37989
rect 280715 37961 280749 37989
rect 280777 37961 280811 37989
rect 280839 37961 280887 37989
rect 280577 29175 280887 37961
rect 280577 29147 280625 29175
rect 280653 29147 280687 29175
rect 280715 29147 280749 29175
rect 280777 29147 280811 29175
rect 280839 29147 280887 29175
rect 280577 29113 280887 29147
rect 280577 29085 280625 29113
rect 280653 29085 280687 29113
rect 280715 29085 280749 29113
rect 280777 29085 280811 29113
rect 280839 29085 280887 29113
rect 280577 29051 280887 29085
rect 280577 29023 280625 29051
rect 280653 29023 280687 29051
rect 280715 29023 280749 29051
rect 280777 29023 280811 29051
rect 280839 29023 280887 29051
rect 280577 28989 280887 29023
rect 280577 28961 280625 28989
rect 280653 28961 280687 28989
rect 280715 28961 280749 28989
rect 280777 28961 280811 28989
rect 280839 28961 280887 28989
rect 280577 20175 280887 28961
rect 280577 20147 280625 20175
rect 280653 20147 280687 20175
rect 280715 20147 280749 20175
rect 280777 20147 280811 20175
rect 280839 20147 280887 20175
rect 280577 20113 280887 20147
rect 280577 20085 280625 20113
rect 280653 20085 280687 20113
rect 280715 20085 280749 20113
rect 280777 20085 280811 20113
rect 280839 20085 280887 20113
rect 280577 20051 280887 20085
rect 280577 20023 280625 20051
rect 280653 20023 280687 20051
rect 280715 20023 280749 20051
rect 280777 20023 280811 20051
rect 280839 20023 280887 20051
rect 280577 19989 280887 20023
rect 280577 19961 280625 19989
rect 280653 19961 280687 19989
rect 280715 19961 280749 19989
rect 280777 19961 280811 19989
rect 280839 19961 280887 19989
rect 280577 11175 280887 19961
rect 280577 11147 280625 11175
rect 280653 11147 280687 11175
rect 280715 11147 280749 11175
rect 280777 11147 280811 11175
rect 280839 11147 280887 11175
rect 280577 11113 280887 11147
rect 280577 11085 280625 11113
rect 280653 11085 280687 11113
rect 280715 11085 280749 11113
rect 280777 11085 280811 11113
rect 280839 11085 280887 11113
rect 280577 11051 280887 11085
rect 280577 11023 280625 11051
rect 280653 11023 280687 11051
rect 280715 11023 280749 11051
rect 280777 11023 280811 11051
rect 280839 11023 280887 11051
rect 280577 10989 280887 11023
rect 280577 10961 280625 10989
rect 280653 10961 280687 10989
rect 280715 10961 280749 10989
rect 280777 10961 280811 10989
rect 280839 10961 280887 10989
rect 280577 2175 280887 10961
rect 280577 2147 280625 2175
rect 280653 2147 280687 2175
rect 280715 2147 280749 2175
rect 280777 2147 280811 2175
rect 280839 2147 280887 2175
rect 280577 2113 280887 2147
rect 280577 2085 280625 2113
rect 280653 2085 280687 2113
rect 280715 2085 280749 2113
rect 280777 2085 280811 2113
rect 280839 2085 280887 2113
rect 280577 2051 280887 2085
rect 280577 2023 280625 2051
rect 280653 2023 280687 2051
rect 280715 2023 280749 2051
rect 280777 2023 280811 2051
rect 280839 2023 280887 2051
rect 280577 1989 280887 2023
rect 280577 1961 280625 1989
rect 280653 1961 280687 1989
rect 280715 1961 280749 1989
rect 280777 1961 280811 1989
rect 280839 1961 280887 1989
rect 280577 -80 280887 1961
rect 280577 -108 280625 -80
rect 280653 -108 280687 -80
rect 280715 -108 280749 -80
rect 280777 -108 280811 -80
rect 280839 -108 280887 -80
rect 280577 -142 280887 -108
rect 280577 -170 280625 -142
rect 280653 -170 280687 -142
rect 280715 -170 280749 -142
rect 280777 -170 280811 -142
rect 280839 -170 280887 -142
rect 280577 -204 280887 -170
rect 280577 -232 280625 -204
rect 280653 -232 280687 -204
rect 280715 -232 280749 -204
rect 280777 -232 280811 -204
rect 280839 -232 280887 -204
rect 280577 -266 280887 -232
rect 280577 -294 280625 -266
rect 280653 -294 280687 -266
rect 280715 -294 280749 -266
rect 280777 -294 280811 -266
rect 280839 -294 280887 -266
rect 280577 -822 280887 -294
rect 282437 299086 282747 299134
rect 282437 299058 282485 299086
rect 282513 299058 282547 299086
rect 282575 299058 282609 299086
rect 282637 299058 282671 299086
rect 282699 299058 282747 299086
rect 282437 299024 282747 299058
rect 282437 298996 282485 299024
rect 282513 298996 282547 299024
rect 282575 298996 282609 299024
rect 282637 298996 282671 299024
rect 282699 298996 282747 299024
rect 282437 298962 282747 298996
rect 282437 298934 282485 298962
rect 282513 298934 282547 298962
rect 282575 298934 282609 298962
rect 282637 298934 282671 298962
rect 282699 298934 282747 298962
rect 282437 298900 282747 298934
rect 282437 298872 282485 298900
rect 282513 298872 282547 298900
rect 282575 298872 282609 298900
rect 282637 298872 282671 298900
rect 282699 298872 282747 298900
rect 282437 293175 282747 298872
rect 282437 293147 282485 293175
rect 282513 293147 282547 293175
rect 282575 293147 282609 293175
rect 282637 293147 282671 293175
rect 282699 293147 282747 293175
rect 282437 293113 282747 293147
rect 282437 293085 282485 293113
rect 282513 293085 282547 293113
rect 282575 293085 282609 293113
rect 282637 293085 282671 293113
rect 282699 293085 282747 293113
rect 282437 293051 282747 293085
rect 282437 293023 282485 293051
rect 282513 293023 282547 293051
rect 282575 293023 282609 293051
rect 282637 293023 282671 293051
rect 282699 293023 282747 293051
rect 282437 292989 282747 293023
rect 282437 292961 282485 292989
rect 282513 292961 282547 292989
rect 282575 292961 282609 292989
rect 282637 292961 282671 292989
rect 282699 292961 282747 292989
rect 282437 284175 282747 292961
rect 282437 284147 282485 284175
rect 282513 284147 282547 284175
rect 282575 284147 282609 284175
rect 282637 284147 282671 284175
rect 282699 284147 282747 284175
rect 282437 284113 282747 284147
rect 282437 284085 282485 284113
rect 282513 284085 282547 284113
rect 282575 284085 282609 284113
rect 282637 284085 282671 284113
rect 282699 284085 282747 284113
rect 282437 284051 282747 284085
rect 282437 284023 282485 284051
rect 282513 284023 282547 284051
rect 282575 284023 282609 284051
rect 282637 284023 282671 284051
rect 282699 284023 282747 284051
rect 282437 283989 282747 284023
rect 282437 283961 282485 283989
rect 282513 283961 282547 283989
rect 282575 283961 282609 283989
rect 282637 283961 282671 283989
rect 282699 283961 282747 283989
rect 282437 275175 282747 283961
rect 282437 275147 282485 275175
rect 282513 275147 282547 275175
rect 282575 275147 282609 275175
rect 282637 275147 282671 275175
rect 282699 275147 282747 275175
rect 282437 275113 282747 275147
rect 282437 275085 282485 275113
rect 282513 275085 282547 275113
rect 282575 275085 282609 275113
rect 282637 275085 282671 275113
rect 282699 275085 282747 275113
rect 282437 275051 282747 275085
rect 282437 275023 282485 275051
rect 282513 275023 282547 275051
rect 282575 275023 282609 275051
rect 282637 275023 282671 275051
rect 282699 275023 282747 275051
rect 282437 274989 282747 275023
rect 282437 274961 282485 274989
rect 282513 274961 282547 274989
rect 282575 274961 282609 274989
rect 282637 274961 282671 274989
rect 282699 274961 282747 274989
rect 282437 266175 282747 274961
rect 282437 266147 282485 266175
rect 282513 266147 282547 266175
rect 282575 266147 282609 266175
rect 282637 266147 282671 266175
rect 282699 266147 282747 266175
rect 282437 266113 282747 266147
rect 282437 266085 282485 266113
rect 282513 266085 282547 266113
rect 282575 266085 282609 266113
rect 282637 266085 282671 266113
rect 282699 266085 282747 266113
rect 282437 266051 282747 266085
rect 282437 266023 282485 266051
rect 282513 266023 282547 266051
rect 282575 266023 282609 266051
rect 282637 266023 282671 266051
rect 282699 266023 282747 266051
rect 282437 265989 282747 266023
rect 282437 265961 282485 265989
rect 282513 265961 282547 265989
rect 282575 265961 282609 265989
rect 282637 265961 282671 265989
rect 282699 265961 282747 265989
rect 282437 257175 282747 265961
rect 282437 257147 282485 257175
rect 282513 257147 282547 257175
rect 282575 257147 282609 257175
rect 282637 257147 282671 257175
rect 282699 257147 282747 257175
rect 282437 257113 282747 257147
rect 282437 257085 282485 257113
rect 282513 257085 282547 257113
rect 282575 257085 282609 257113
rect 282637 257085 282671 257113
rect 282699 257085 282747 257113
rect 282437 257051 282747 257085
rect 282437 257023 282485 257051
rect 282513 257023 282547 257051
rect 282575 257023 282609 257051
rect 282637 257023 282671 257051
rect 282699 257023 282747 257051
rect 282437 256989 282747 257023
rect 282437 256961 282485 256989
rect 282513 256961 282547 256989
rect 282575 256961 282609 256989
rect 282637 256961 282671 256989
rect 282699 256961 282747 256989
rect 282437 248175 282747 256961
rect 282437 248147 282485 248175
rect 282513 248147 282547 248175
rect 282575 248147 282609 248175
rect 282637 248147 282671 248175
rect 282699 248147 282747 248175
rect 282437 248113 282747 248147
rect 282437 248085 282485 248113
rect 282513 248085 282547 248113
rect 282575 248085 282609 248113
rect 282637 248085 282671 248113
rect 282699 248085 282747 248113
rect 282437 248051 282747 248085
rect 282437 248023 282485 248051
rect 282513 248023 282547 248051
rect 282575 248023 282609 248051
rect 282637 248023 282671 248051
rect 282699 248023 282747 248051
rect 282437 247989 282747 248023
rect 282437 247961 282485 247989
rect 282513 247961 282547 247989
rect 282575 247961 282609 247989
rect 282637 247961 282671 247989
rect 282699 247961 282747 247989
rect 282437 239175 282747 247961
rect 282437 239147 282485 239175
rect 282513 239147 282547 239175
rect 282575 239147 282609 239175
rect 282637 239147 282671 239175
rect 282699 239147 282747 239175
rect 282437 239113 282747 239147
rect 282437 239085 282485 239113
rect 282513 239085 282547 239113
rect 282575 239085 282609 239113
rect 282637 239085 282671 239113
rect 282699 239085 282747 239113
rect 282437 239051 282747 239085
rect 282437 239023 282485 239051
rect 282513 239023 282547 239051
rect 282575 239023 282609 239051
rect 282637 239023 282671 239051
rect 282699 239023 282747 239051
rect 282437 238989 282747 239023
rect 282437 238961 282485 238989
rect 282513 238961 282547 238989
rect 282575 238961 282609 238989
rect 282637 238961 282671 238989
rect 282699 238961 282747 238989
rect 282437 230175 282747 238961
rect 282437 230147 282485 230175
rect 282513 230147 282547 230175
rect 282575 230147 282609 230175
rect 282637 230147 282671 230175
rect 282699 230147 282747 230175
rect 282437 230113 282747 230147
rect 282437 230085 282485 230113
rect 282513 230085 282547 230113
rect 282575 230085 282609 230113
rect 282637 230085 282671 230113
rect 282699 230085 282747 230113
rect 282437 230051 282747 230085
rect 282437 230023 282485 230051
rect 282513 230023 282547 230051
rect 282575 230023 282609 230051
rect 282637 230023 282671 230051
rect 282699 230023 282747 230051
rect 282437 229989 282747 230023
rect 282437 229961 282485 229989
rect 282513 229961 282547 229989
rect 282575 229961 282609 229989
rect 282637 229961 282671 229989
rect 282699 229961 282747 229989
rect 282437 221175 282747 229961
rect 282437 221147 282485 221175
rect 282513 221147 282547 221175
rect 282575 221147 282609 221175
rect 282637 221147 282671 221175
rect 282699 221147 282747 221175
rect 282437 221113 282747 221147
rect 282437 221085 282485 221113
rect 282513 221085 282547 221113
rect 282575 221085 282609 221113
rect 282637 221085 282671 221113
rect 282699 221085 282747 221113
rect 282437 221051 282747 221085
rect 282437 221023 282485 221051
rect 282513 221023 282547 221051
rect 282575 221023 282609 221051
rect 282637 221023 282671 221051
rect 282699 221023 282747 221051
rect 282437 220989 282747 221023
rect 282437 220961 282485 220989
rect 282513 220961 282547 220989
rect 282575 220961 282609 220989
rect 282637 220961 282671 220989
rect 282699 220961 282747 220989
rect 282437 212175 282747 220961
rect 282437 212147 282485 212175
rect 282513 212147 282547 212175
rect 282575 212147 282609 212175
rect 282637 212147 282671 212175
rect 282699 212147 282747 212175
rect 282437 212113 282747 212147
rect 282437 212085 282485 212113
rect 282513 212085 282547 212113
rect 282575 212085 282609 212113
rect 282637 212085 282671 212113
rect 282699 212085 282747 212113
rect 282437 212051 282747 212085
rect 282437 212023 282485 212051
rect 282513 212023 282547 212051
rect 282575 212023 282609 212051
rect 282637 212023 282671 212051
rect 282699 212023 282747 212051
rect 282437 211989 282747 212023
rect 282437 211961 282485 211989
rect 282513 211961 282547 211989
rect 282575 211961 282609 211989
rect 282637 211961 282671 211989
rect 282699 211961 282747 211989
rect 282437 203175 282747 211961
rect 282437 203147 282485 203175
rect 282513 203147 282547 203175
rect 282575 203147 282609 203175
rect 282637 203147 282671 203175
rect 282699 203147 282747 203175
rect 282437 203113 282747 203147
rect 282437 203085 282485 203113
rect 282513 203085 282547 203113
rect 282575 203085 282609 203113
rect 282637 203085 282671 203113
rect 282699 203085 282747 203113
rect 282437 203051 282747 203085
rect 282437 203023 282485 203051
rect 282513 203023 282547 203051
rect 282575 203023 282609 203051
rect 282637 203023 282671 203051
rect 282699 203023 282747 203051
rect 282437 202989 282747 203023
rect 282437 202961 282485 202989
rect 282513 202961 282547 202989
rect 282575 202961 282609 202989
rect 282637 202961 282671 202989
rect 282699 202961 282747 202989
rect 282437 194175 282747 202961
rect 282437 194147 282485 194175
rect 282513 194147 282547 194175
rect 282575 194147 282609 194175
rect 282637 194147 282671 194175
rect 282699 194147 282747 194175
rect 282437 194113 282747 194147
rect 282437 194085 282485 194113
rect 282513 194085 282547 194113
rect 282575 194085 282609 194113
rect 282637 194085 282671 194113
rect 282699 194085 282747 194113
rect 282437 194051 282747 194085
rect 282437 194023 282485 194051
rect 282513 194023 282547 194051
rect 282575 194023 282609 194051
rect 282637 194023 282671 194051
rect 282699 194023 282747 194051
rect 282437 193989 282747 194023
rect 282437 193961 282485 193989
rect 282513 193961 282547 193989
rect 282575 193961 282609 193989
rect 282637 193961 282671 193989
rect 282699 193961 282747 193989
rect 282437 185175 282747 193961
rect 282437 185147 282485 185175
rect 282513 185147 282547 185175
rect 282575 185147 282609 185175
rect 282637 185147 282671 185175
rect 282699 185147 282747 185175
rect 282437 185113 282747 185147
rect 282437 185085 282485 185113
rect 282513 185085 282547 185113
rect 282575 185085 282609 185113
rect 282637 185085 282671 185113
rect 282699 185085 282747 185113
rect 282437 185051 282747 185085
rect 282437 185023 282485 185051
rect 282513 185023 282547 185051
rect 282575 185023 282609 185051
rect 282637 185023 282671 185051
rect 282699 185023 282747 185051
rect 282437 184989 282747 185023
rect 282437 184961 282485 184989
rect 282513 184961 282547 184989
rect 282575 184961 282609 184989
rect 282637 184961 282671 184989
rect 282699 184961 282747 184989
rect 282437 176175 282747 184961
rect 282437 176147 282485 176175
rect 282513 176147 282547 176175
rect 282575 176147 282609 176175
rect 282637 176147 282671 176175
rect 282699 176147 282747 176175
rect 282437 176113 282747 176147
rect 282437 176085 282485 176113
rect 282513 176085 282547 176113
rect 282575 176085 282609 176113
rect 282637 176085 282671 176113
rect 282699 176085 282747 176113
rect 282437 176051 282747 176085
rect 282437 176023 282485 176051
rect 282513 176023 282547 176051
rect 282575 176023 282609 176051
rect 282637 176023 282671 176051
rect 282699 176023 282747 176051
rect 282437 175989 282747 176023
rect 282437 175961 282485 175989
rect 282513 175961 282547 175989
rect 282575 175961 282609 175989
rect 282637 175961 282671 175989
rect 282699 175961 282747 175989
rect 282437 167175 282747 175961
rect 282437 167147 282485 167175
rect 282513 167147 282547 167175
rect 282575 167147 282609 167175
rect 282637 167147 282671 167175
rect 282699 167147 282747 167175
rect 282437 167113 282747 167147
rect 282437 167085 282485 167113
rect 282513 167085 282547 167113
rect 282575 167085 282609 167113
rect 282637 167085 282671 167113
rect 282699 167085 282747 167113
rect 282437 167051 282747 167085
rect 282437 167023 282485 167051
rect 282513 167023 282547 167051
rect 282575 167023 282609 167051
rect 282637 167023 282671 167051
rect 282699 167023 282747 167051
rect 282437 166989 282747 167023
rect 282437 166961 282485 166989
rect 282513 166961 282547 166989
rect 282575 166961 282609 166989
rect 282637 166961 282671 166989
rect 282699 166961 282747 166989
rect 282437 158175 282747 166961
rect 282437 158147 282485 158175
rect 282513 158147 282547 158175
rect 282575 158147 282609 158175
rect 282637 158147 282671 158175
rect 282699 158147 282747 158175
rect 282437 158113 282747 158147
rect 282437 158085 282485 158113
rect 282513 158085 282547 158113
rect 282575 158085 282609 158113
rect 282637 158085 282671 158113
rect 282699 158085 282747 158113
rect 282437 158051 282747 158085
rect 282437 158023 282485 158051
rect 282513 158023 282547 158051
rect 282575 158023 282609 158051
rect 282637 158023 282671 158051
rect 282699 158023 282747 158051
rect 282437 157989 282747 158023
rect 282437 157961 282485 157989
rect 282513 157961 282547 157989
rect 282575 157961 282609 157989
rect 282637 157961 282671 157989
rect 282699 157961 282747 157989
rect 282437 149175 282747 157961
rect 282437 149147 282485 149175
rect 282513 149147 282547 149175
rect 282575 149147 282609 149175
rect 282637 149147 282671 149175
rect 282699 149147 282747 149175
rect 282437 149113 282747 149147
rect 282437 149085 282485 149113
rect 282513 149085 282547 149113
rect 282575 149085 282609 149113
rect 282637 149085 282671 149113
rect 282699 149085 282747 149113
rect 282437 149051 282747 149085
rect 282437 149023 282485 149051
rect 282513 149023 282547 149051
rect 282575 149023 282609 149051
rect 282637 149023 282671 149051
rect 282699 149023 282747 149051
rect 282437 148989 282747 149023
rect 282437 148961 282485 148989
rect 282513 148961 282547 148989
rect 282575 148961 282609 148989
rect 282637 148961 282671 148989
rect 282699 148961 282747 148989
rect 282437 140175 282747 148961
rect 282437 140147 282485 140175
rect 282513 140147 282547 140175
rect 282575 140147 282609 140175
rect 282637 140147 282671 140175
rect 282699 140147 282747 140175
rect 282437 140113 282747 140147
rect 282437 140085 282485 140113
rect 282513 140085 282547 140113
rect 282575 140085 282609 140113
rect 282637 140085 282671 140113
rect 282699 140085 282747 140113
rect 282437 140051 282747 140085
rect 282437 140023 282485 140051
rect 282513 140023 282547 140051
rect 282575 140023 282609 140051
rect 282637 140023 282671 140051
rect 282699 140023 282747 140051
rect 282437 139989 282747 140023
rect 282437 139961 282485 139989
rect 282513 139961 282547 139989
rect 282575 139961 282609 139989
rect 282637 139961 282671 139989
rect 282699 139961 282747 139989
rect 282437 131175 282747 139961
rect 282437 131147 282485 131175
rect 282513 131147 282547 131175
rect 282575 131147 282609 131175
rect 282637 131147 282671 131175
rect 282699 131147 282747 131175
rect 282437 131113 282747 131147
rect 282437 131085 282485 131113
rect 282513 131085 282547 131113
rect 282575 131085 282609 131113
rect 282637 131085 282671 131113
rect 282699 131085 282747 131113
rect 282437 131051 282747 131085
rect 282437 131023 282485 131051
rect 282513 131023 282547 131051
rect 282575 131023 282609 131051
rect 282637 131023 282671 131051
rect 282699 131023 282747 131051
rect 282437 130989 282747 131023
rect 282437 130961 282485 130989
rect 282513 130961 282547 130989
rect 282575 130961 282609 130989
rect 282637 130961 282671 130989
rect 282699 130961 282747 130989
rect 282437 122175 282747 130961
rect 282437 122147 282485 122175
rect 282513 122147 282547 122175
rect 282575 122147 282609 122175
rect 282637 122147 282671 122175
rect 282699 122147 282747 122175
rect 282437 122113 282747 122147
rect 282437 122085 282485 122113
rect 282513 122085 282547 122113
rect 282575 122085 282609 122113
rect 282637 122085 282671 122113
rect 282699 122085 282747 122113
rect 282437 122051 282747 122085
rect 282437 122023 282485 122051
rect 282513 122023 282547 122051
rect 282575 122023 282609 122051
rect 282637 122023 282671 122051
rect 282699 122023 282747 122051
rect 282437 121989 282747 122023
rect 282437 121961 282485 121989
rect 282513 121961 282547 121989
rect 282575 121961 282609 121989
rect 282637 121961 282671 121989
rect 282699 121961 282747 121989
rect 282437 113175 282747 121961
rect 282437 113147 282485 113175
rect 282513 113147 282547 113175
rect 282575 113147 282609 113175
rect 282637 113147 282671 113175
rect 282699 113147 282747 113175
rect 282437 113113 282747 113147
rect 282437 113085 282485 113113
rect 282513 113085 282547 113113
rect 282575 113085 282609 113113
rect 282637 113085 282671 113113
rect 282699 113085 282747 113113
rect 282437 113051 282747 113085
rect 282437 113023 282485 113051
rect 282513 113023 282547 113051
rect 282575 113023 282609 113051
rect 282637 113023 282671 113051
rect 282699 113023 282747 113051
rect 282437 112989 282747 113023
rect 282437 112961 282485 112989
rect 282513 112961 282547 112989
rect 282575 112961 282609 112989
rect 282637 112961 282671 112989
rect 282699 112961 282747 112989
rect 282437 104175 282747 112961
rect 282437 104147 282485 104175
rect 282513 104147 282547 104175
rect 282575 104147 282609 104175
rect 282637 104147 282671 104175
rect 282699 104147 282747 104175
rect 282437 104113 282747 104147
rect 282437 104085 282485 104113
rect 282513 104085 282547 104113
rect 282575 104085 282609 104113
rect 282637 104085 282671 104113
rect 282699 104085 282747 104113
rect 282437 104051 282747 104085
rect 282437 104023 282485 104051
rect 282513 104023 282547 104051
rect 282575 104023 282609 104051
rect 282637 104023 282671 104051
rect 282699 104023 282747 104051
rect 282437 103989 282747 104023
rect 282437 103961 282485 103989
rect 282513 103961 282547 103989
rect 282575 103961 282609 103989
rect 282637 103961 282671 103989
rect 282699 103961 282747 103989
rect 282437 95175 282747 103961
rect 282437 95147 282485 95175
rect 282513 95147 282547 95175
rect 282575 95147 282609 95175
rect 282637 95147 282671 95175
rect 282699 95147 282747 95175
rect 282437 95113 282747 95147
rect 282437 95085 282485 95113
rect 282513 95085 282547 95113
rect 282575 95085 282609 95113
rect 282637 95085 282671 95113
rect 282699 95085 282747 95113
rect 282437 95051 282747 95085
rect 282437 95023 282485 95051
rect 282513 95023 282547 95051
rect 282575 95023 282609 95051
rect 282637 95023 282671 95051
rect 282699 95023 282747 95051
rect 282437 94989 282747 95023
rect 282437 94961 282485 94989
rect 282513 94961 282547 94989
rect 282575 94961 282609 94989
rect 282637 94961 282671 94989
rect 282699 94961 282747 94989
rect 282437 86175 282747 94961
rect 282437 86147 282485 86175
rect 282513 86147 282547 86175
rect 282575 86147 282609 86175
rect 282637 86147 282671 86175
rect 282699 86147 282747 86175
rect 282437 86113 282747 86147
rect 282437 86085 282485 86113
rect 282513 86085 282547 86113
rect 282575 86085 282609 86113
rect 282637 86085 282671 86113
rect 282699 86085 282747 86113
rect 282437 86051 282747 86085
rect 282437 86023 282485 86051
rect 282513 86023 282547 86051
rect 282575 86023 282609 86051
rect 282637 86023 282671 86051
rect 282699 86023 282747 86051
rect 282437 85989 282747 86023
rect 282437 85961 282485 85989
rect 282513 85961 282547 85989
rect 282575 85961 282609 85989
rect 282637 85961 282671 85989
rect 282699 85961 282747 85989
rect 282437 77175 282747 85961
rect 282437 77147 282485 77175
rect 282513 77147 282547 77175
rect 282575 77147 282609 77175
rect 282637 77147 282671 77175
rect 282699 77147 282747 77175
rect 282437 77113 282747 77147
rect 282437 77085 282485 77113
rect 282513 77085 282547 77113
rect 282575 77085 282609 77113
rect 282637 77085 282671 77113
rect 282699 77085 282747 77113
rect 282437 77051 282747 77085
rect 282437 77023 282485 77051
rect 282513 77023 282547 77051
rect 282575 77023 282609 77051
rect 282637 77023 282671 77051
rect 282699 77023 282747 77051
rect 282437 76989 282747 77023
rect 282437 76961 282485 76989
rect 282513 76961 282547 76989
rect 282575 76961 282609 76989
rect 282637 76961 282671 76989
rect 282699 76961 282747 76989
rect 282437 68175 282747 76961
rect 282437 68147 282485 68175
rect 282513 68147 282547 68175
rect 282575 68147 282609 68175
rect 282637 68147 282671 68175
rect 282699 68147 282747 68175
rect 282437 68113 282747 68147
rect 282437 68085 282485 68113
rect 282513 68085 282547 68113
rect 282575 68085 282609 68113
rect 282637 68085 282671 68113
rect 282699 68085 282747 68113
rect 282437 68051 282747 68085
rect 282437 68023 282485 68051
rect 282513 68023 282547 68051
rect 282575 68023 282609 68051
rect 282637 68023 282671 68051
rect 282699 68023 282747 68051
rect 282437 67989 282747 68023
rect 282437 67961 282485 67989
rect 282513 67961 282547 67989
rect 282575 67961 282609 67989
rect 282637 67961 282671 67989
rect 282699 67961 282747 67989
rect 282437 59175 282747 67961
rect 282437 59147 282485 59175
rect 282513 59147 282547 59175
rect 282575 59147 282609 59175
rect 282637 59147 282671 59175
rect 282699 59147 282747 59175
rect 282437 59113 282747 59147
rect 282437 59085 282485 59113
rect 282513 59085 282547 59113
rect 282575 59085 282609 59113
rect 282637 59085 282671 59113
rect 282699 59085 282747 59113
rect 282437 59051 282747 59085
rect 282437 59023 282485 59051
rect 282513 59023 282547 59051
rect 282575 59023 282609 59051
rect 282637 59023 282671 59051
rect 282699 59023 282747 59051
rect 282437 58989 282747 59023
rect 282437 58961 282485 58989
rect 282513 58961 282547 58989
rect 282575 58961 282609 58989
rect 282637 58961 282671 58989
rect 282699 58961 282747 58989
rect 282437 50175 282747 58961
rect 282437 50147 282485 50175
rect 282513 50147 282547 50175
rect 282575 50147 282609 50175
rect 282637 50147 282671 50175
rect 282699 50147 282747 50175
rect 282437 50113 282747 50147
rect 282437 50085 282485 50113
rect 282513 50085 282547 50113
rect 282575 50085 282609 50113
rect 282637 50085 282671 50113
rect 282699 50085 282747 50113
rect 282437 50051 282747 50085
rect 282437 50023 282485 50051
rect 282513 50023 282547 50051
rect 282575 50023 282609 50051
rect 282637 50023 282671 50051
rect 282699 50023 282747 50051
rect 282437 49989 282747 50023
rect 282437 49961 282485 49989
rect 282513 49961 282547 49989
rect 282575 49961 282609 49989
rect 282637 49961 282671 49989
rect 282699 49961 282747 49989
rect 282437 41175 282747 49961
rect 282437 41147 282485 41175
rect 282513 41147 282547 41175
rect 282575 41147 282609 41175
rect 282637 41147 282671 41175
rect 282699 41147 282747 41175
rect 282437 41113 282747 41147
rect 282437 41085 282485 41113
rect 282513 41085 282547 41113
rect 282575 41085 282609 41113
rect 282637 41085 282671 41113
rect 282699 41085 282747 41113
rect 282437 41051 282747 41085
rect 282437 41023 282485 41051
rect 282513 41023 282547 41051
rect 282575 41023 282609 41051
rect 282637 41023 282671 41051
rect 282699 41023 282747 41051
rect 282437 40989 282747 41023
rect 282437 40961 282485 40989
rect 282513 40961 282547 40989
rect 282575 40961 282609 40989
rect 282637 40961 282671 40989
rect 282699 40961 282747 40989
rect 282437 32175 282747 40961
rect 282437 32147 282485 32175
rect 282513 32147 282547 32175
rect 282575 32147 282609 32175
rect 282637 32147 282671 32175
rect 282699 32147 282747 32175
rect 282437 32113 282747 32147
rect 282437 32085 282485 32113
rect 282513 32085 282547 32113
rect 282575 32085 282609 32113
rect 282637 32085 282671 32113
rect 282699 32085 282747 32113
rect 282437 32051 282747 32085
rect 282437 32023 282485 32051
rect 282513 32023 282547 32051
rect 282575 32023 282609 32051
rect 282637 32023 282671 32051
rect 282699 32023 282747 32051
rect 282437 31989 282747 32023
rect 282437 31961 282485 31989
rect 282513 31961 282547 31989
rect 282575 31961 282609 31989
rect 282637 31961 282671 31989
rect 282699 31961 282747 31989
rect 282437 23175 282747 31961
rect 282437 23147 282485 23175
rect 282513 23147 282547 23175
rect 282575 23147 282609 23175
rect 282637 23147 282671 23175
rect 282699 23147 282747 23175
rect 282437 23113 282747 23147
rect 282437 23085 282485 23113
rect 282513 23085 282547 23113
rect 282575 23085 282609 23113
rect 282637 23085 282671 23113
rect 282699 23085 282747 23113
rect 282437 23051 282747 23085
rect 282437 23023 282485 23051
rect 282513 23023 282547 23051
rect 282575 23023 282609 23051
rect 282637 23023 282671 23051
rect 282699 23023 282747 23051
rect 282437 22989 282747 23023
rect 282437 22961 282485 22989
rect 282513 22961 282547 22989
rect 282575 22961 282609 22989
rect 282637 22961 282671 22989
rect 282699 22961 282747 22989
rect 282437 14175 282747 22961
rect 282437 14147 282485 14175
rect 282513 14147 282547 14175
rect 282575 14147 282609 14175
rect 282637 14147 282671 14175
rect 282699 14147 282747 14175
rect 282437 14113 282747 14147
rect 282437 14085 282485 14113
rect 282513 14085 282547 14113
rect 282575 14085 282609 14113
rect 282637 14085 282671 14113
rect 282699 14085 282747 14113
rect 282437 14051 282747 14085
rect 282437 14023 282485 14051
rect 282513 14023 282547 14051
rect 282575 14023 282609 14051
rect 282637 14023 282671 14051
rect 282699 14023 282747 14051
rect 282437 13989 282747 14023
rect 282437 13961 282485 13989
rect 282513 13961 282547 13989
rect 282575 13961 282609 13989
rect 282637 13961 282671 13989
rect 282699 13961 282747 13989
rect 282437 5175 282747 13961
rect 282437 5147 282485 5175
rect 282513 5147 282547 5175
rect 282575 5147 282609 5175
rect 282637 5147 282671 5175
rect 282699 5147 282747 5175
rect 282437 5113 282747 5147
rect 282437 5085 282485 5113
rect 282513 5085 282547 5113
rect 282575 5085 282609 5113
rect 282637 5085 282671 5113
rect 282699 5085 282747 5113
rect 282437 5051 282747 5085
rect 282437 5023 282485 5051
rect 282513 5023 282547 5051
rect 282575 5023 282609 5051
rect 282637 5023 282671 5051
rect 282699 5023 282747 5051
rect 282437 4989 282747 5023
rect 282437 4961 282485 4989
rect 282513 4961 282547 4989
rect 282575 4961 282609 4989
rect 282637 4961 282671 4989
rect 282699 4961 282747 4989
rect 282437 -560 282747 4961
rect 282437 -588 282485 -560
rect 282513 -588 282547 -560
rect 282575 -588 282609 -560
rect 282637 -588 282671 -560
rect 282699 -588 282747 -560
rect 282437 -622 282747 -588
rect 282437 -650 282485 -622
rect 282513 -650 282547 -622
rect 282575 -650 282609 -622
rect 282637 -650 282671 -622
rect 282699 -650 282747 -622
rect 282437 -684 282747 -650
rect 282437 -712 282485 -684
rect 282513 -712 282547 -684
rect 282575 -712 282609 -684
rect 282637 -712 282671 -684
rect 282699 -712 282747 -684
rect 282437 -746 282747 -712
rect 282437 -774 282485 -746
rect 282513 -774 282547 -746
rect 282575 -774 282609 -746
rect 282637 -774 282671 -746
rect 282699 -774 282747 -746
rect 282437 -822 282747 -774
rect 289577 298606 289887 299134
rect 289577 298578 289625 298606
rect 289653 298578 289687 298606
rect 289715 298578 289749 298606
rect 289777 298578 289811 298606
rect 289839 298578 289887 298606
rect 289577 298544 289887 298578
rect 289577 298516 289625 298544
rect 289653 298516 289687 298544
rect 289715 298516 289749 298544
rect 289777 298516 289811 298544
rect 289839 298516 289887 298544
rect 289577 298482 289887 298516
rect 289577 298454 289625 298482
rect 289653 298454 289687 298482
rect 289715 298454 289749 298482
rect 289777 298454 289811 298482
rect 289839 298454 289887 298482
rect 289577 298420 289887 298454
rect 289577 298392 289625 298420
rect 289653 298392 289687 298420
rect 289715 298392 289749 298420
rect 289777 298392 289811 298420
rect 289839 298392 289887 298420
rect 289577 290175 289887 298392
rect 289577 290147 289625 290175
rect 289653 290147 289687 290175
rect 289715 290147 289749 290175
rect 289777 290147 289811 290175
rect 289839 290147 289887 290175
rect 289577 290113 289887 290147
rect 289577 290085 289625 290113
rect 289653 290085 289687 290113
rect 289715 290085 289749 290113
rect 289777 290085 289811 290113
rect 289839 290085 289887 290113
rect 289577 290051 289887 290085
rect 289577 290023 289625 290051
rect 289653 290023 289687 290051
rect 289715 290023 289749 290051
rect 289777 290023 289811 290051
rect 289839 290023 289887 290051
rect 289577 289989 289887 290023
rect 289577 289961 289625 289989
rect 289653 289961 289687 289989
rect 289715 289961 289749 289989
rect 289777 289961 289811 289989
rect 289839 289961 289887 289989
rect 289577 281175 289887 289961
rect 289577 281147 289625 281175
rect 289653 281147 289687 281175
rect 289715 281147 289749 281175
rect 289777 281147 289811 281175
rect 289839 281147 289887 281175
rect 289577 281113 289887 281147
rect 289577 281085 289625 281113
rect 289653 281085 289687 281113
rect 289715 281085 289749 281113
rect 289777 281085 289811 281113
rect 289839 281085 289887 281113
rect 289577 281051 289887 281085
rect 289577 281023 289625 281051
rect 289653 281023 289687 281051
rect 289715 281023 289749 281051
rect 289777 281023 289811 281051
rect 289839 281023 289887 281051
rect 289577 280989 289887 281023
rect 289577 280961 289625 280989
rect 289653 280961 289687 280989
rect 289715 280961 289749 280989
rect 289777 280961 289811 280989
rect 289839 280961 289887 280989
rect 289577 272175 289887 280961
rect 289577 272147 289625 272175
rect 289653 272147 289687 272175
rect 289715 272147 289749 272175
rect 289777 272147 289811 272175
rect 289839 272147 289887 272175
rect 289577 272113 289887 272147
rect 289577 272085 289625 272113
rect 289653 272085 289687 272113
rect 289715 272085 289749 272113
rect 289777 272085 289811 272113
rect 289839 272085 289887 272113
rect 289577 272051 289887 272085
rect 289577 272023 289625 272051
rect 289653 272023 289687 272051
rect 289715 272023 289749 272051
rect 289777 272023 289811 272051
rect 289839 272023 289887 272051
rect 289577 271989 289887 272023
rect 289577 271961 289625 271989
rect 289653 271961 289687 271989
rect 289715 271961 289749 271989
rect 289777 271961 289811 271989
rect 289839 271961 289887 271989
rect 289577 263175 289887 271961
rect 289577 263147 289625 263175
rect 289653 263147 289687 263175
rect 289715 263147 289749 263175
rect 289777 263147 289811 263175
rect 289839 263147 289887 263175
rect 289577 263113 289887 263147
rect 289577 263085 289625 263113
rect 289653 263085 289687 263113
rect 289715 263085 289749 263113
rect 289777 263085 289811 263113
rect 289839 263085 289887 263113
rect 289577 263051 289887 263085
rect 289577 263023 289625 263051
rect 289653 263023 289687 263051
rect 289715 263023 289749 263051
rect 289777 263023 289811 263051
rect 289839 263023 289887 263051
rect 289577 262989 289887 263023
rect 289577 262961 289625 262989
rect 289653 262961 289687 262989
rect 289715 262961 289749 262989
rect 289777 262961 289811 262989
rect 289839 262961 289887 262989
rect 289577 254175 289887 262961
rect 289577 254147 289625 254175
rect 289653 254147 289687 254175
rect 289715 254147 289749 254175
rect 289777 254147 289811 254175
rect 289839 254147 289887 254175
rect 289577 254113 289887 254147
rect 289577 254085 289625 254113
rect 289653 254085 289687 254113
rect 289715 254085 289749 254113
rect 289777 254085 289811 254113
rect 289839 254085 289887 254113
rect 289577 254051 289887 254085
rect 289577 254023 289625 254051
rect 289653 254023 289687 254051
rect 289715 254023 289749 254051
rect 289777 254023 289811 254051
rect 289839 254023 289887 254051
rect 289577 253989 289887 254023
rect 289577 253961 289625 253989
rect 289653 253961 289687 253989
rect 289715 253961 289749 253989
rect 289777 253961 289811 253989
rect 289839 253961 289887 253989
rect 289577 245175 289887 253961
rect 289577 245147 289625 245175
rect 289653 245147 289687 245175
rect 289715 245147 289749 245175
rect 289777 245147 289811 245175
rect 289839 245147 289887 245175
rect 289577 245113 289887 245147
rect 289577 245085 289625 245113
rect 289653 245085 289687 245113
rect 289715 245085 289749 245113
rect 289777 245085 289811 245113
rect 289839 245085 289887 245113
rect 289577 245051 289887 245085
rect 289577 245023 289625 245051
rect 289653 245023 289687 245051
rect 289715 245023 289749 245051
rect 289777 245023 289811 245051
rect 289839 245023 289887 245051
rect 289577 244989 289887 245023
rect 289577 244961 289625 244989
rect 289653 244961 289687 244989
rect 289715 244961 289749 244989
rect 289777 244961 289811 244989
rect 289839 244961 289887 244989
rect 289577 236175 289887 244961
rect 289577 236147 289625 236175
rect 289653 236147 289687 236175
rect 289715 236147 289749 236175
rect 289777 236147 289811 236175
rect 289839 236147 289887 236175
rect 289577 236113 289887 236147
rect 289577 236085 289625 236113
rect 289653 236085 289687 236113
rect 289715 236085 289749 236113
rect 289777 236085 289811 236113
rect 289839 236085 289887 236113
rect 289577 236051 289887 236085
rect 289577 236023 289625 236051
rect 289653 236023 289687 236051
rect 289715 236023 289749 236051
rect 289777 236023 289811 236051
rect 289839 236023 289887 236051
rect 289577 235989 289887 236023
rect 289577 235961 289625 235989
rect 289653 235961 289687 235989
rect 289715 235961 289749 235989
rect 289777 235961 289811 235989
rect 289839 235961 289887 235989
rect 289577 227175 289887 235961
rect 289577 227147 289625 227175
rect 289653 227147 289687 227175
rect 289715 227147 289749 227175
rect 289777 227147 289811 227175
rect 289839 227147 289887 227175
rect 289577 227113 289887 227147
rect 289577 227085 289625 227113
rect 289653 227085 289687 227113
rect 289715 227085 289749 227113
rect 289777 227085 289811 227113
rect 289839 227085 289887 227113
rect 289577 227051 289887 227085
rect 289577 227023 289625 227051
rect 289653 227023 289687 227051
rect 289715 227023 289749 227051
rect 289777 227023 289811 227051
rect 289839 227023 289887 227051
rect 289577 226989 289887 227023
rect 289577 226961 289625 226989
rect 289653 226961 289687 226989
rect 289715 226961 289749 226989
rect 289777 226961 289811 226989
rect 289839 226961 289887 226989
rect 289577 218175 289887 226961
rect 289577 218147 289625 218175
rect 289653 218147 289687 218175
rect 289715 218147 289749 218175
rect 289777 218147 289811 218175
rect 289839 218147 289887 218175
rect 289577 218113 289887 218147
rect 289577 218085 289625 218113
rect 289653 218085 289687 218113
rect 289715 218085 289749 218113
rect 289777 218085 289811 218113
rect 289839 218085 289887 218113
rect 289577 218051 289887 218085
rect 289577 218023 289625 218051
rect 289653 218023 289687 218051
rect 289715 218023 289749 218051
rect 289777 218023 289811 218051
rect 289839 218023 289887 218051
rect 289577 217989 289887 218023
rect 289577 217961 289625 217989
rect 289653 217961 289687 217989
rect 289715 217961 289749 217989
rect 289777 217961 289811 217989
rect 289839 217961 289887 217989
rect 289577 209175 289887 217961
rect 289577 209147 289625 209175
rect 289653 209147 289687 209175
rect 289715 209147 289749 209175
rect 289777 209147 289811 209175
rect 289839 209147 289887 209175
rect 289577 209113 289887 209147
rect 289577 209085 289625 209113
rect 289653 209085 289687 209113
rect 289715 209085 289749 209113
rect 289777 209085 289811 209113
rect 289839 209085 289887 209113
rect 289577 209051 289887 209085
rect 289577 209023 289625 209051
rect 289653 209023 289687 209051
rect 289715 209023 289749 209051
rect 289777 209023 289811 209051
rect 289839 209023 289887 209051
rect 289577 208989 289887 209023
rect 289577 208961 289625 208989
rect 289653 208961 289687 208989
rect 289715 208961 289749 208989
rect 289777 208961 289811 208989
rect 289839 208961 289887 208989
rect 289577 200175 289887 208961
rect 289577 200147 289625 200175
rect 289653 200147 289687 200175
rect 289715 200147 289749 200175
rect 289777 200147 289811 200175
rect 289839 200147 289887 200175
rect 289577 200113 289887 200147
rect 289577 200085 289625 200113
rect 289653 200085 289687 200113
rect 289715 200085 289749 200113
rect 289777 200085 289811 200113
rect 289839 200085 289887 200113
rect 289577 200051 289887 200085
rect 289577 200023 289625 200051
rect 289653 200023 289687 200051
rect 289715 200023 289749 200051
rect 289777 200023 289811 200051
rect 289839 200023 289887 200051
rect 289577 199989 289887 200023
rect 289577 199961 289625 199989
rect 289653 199961 289687 199989
rect 289715 199961 289749 199989
rect 289777 199961 289811 199989
rect 289839 199961 289887 199989
rect 289577 191175 289887 199961
rect 289577 191147 289625 191175
rect 289653 191147 289687 191175
rect 289715 191147 289749 191175
rect 289777 191147 289811 191175
rect 289839 191147 289887 191175
rect 289577 191113 289887 191147
rect 289577 191085 289625 191113
rect 289653 191085 289687 191113
rect 289715 191085 289749 191113
rect 289777 191085 289811 191113
rect 289839 191085 289887 191113
rect 289577 191051 289887 191085
rect 289577 191023 289625 191051
rect 289653 191023 289687 191051
rect 289715 191023 289749 191051
rect 289777 191023 289811 191051
rect 289839 191023 289887 191051
rect 289577 190989 289887 191023
rect 289577 190961 289625 190989
rect 289653 190961 289687 190989
rect 289715 190961 289749 190989
rect 289777 190961 289811 190989
rect 289839 190961 289887 190989
rect 289577 182175 289887 190961
rect 289577 182147 289625 182175
rect 289653 182147 289687 182175
rect 289715 182147 289749 182175
rect 289777 182147 289811 182175
rect 289839 182147 289887 182175
rect 289577 182113 289887 182147
rect 289577 182085 289625 182113
rect 289653 182085 289687 182113
rect 289715 182085 289749 182113
rect 289777 182085 289811 182113
rect 289839 182085 289887 182113
rect 289577 182051 289887 182085
rect 289577 182023 289625 182051
rect 289653 182023 289687 182051
rect 289715 182023 289749 182051
rect 289777 182023 289811 182051
rect 289839 182023 289887 182051
rect 289577 181989 289887 182023
rect 289577 181961 289625 181989
rect 289653 181961 289687 181989
rect 289715 181961 289749 181989
rect 289777 181961 289811 181989
rect 289839 181961 289887 181989
rect 289577 173175 289887 181961
rect 289577 173147 289625 173175
rect 289653 173147 289687 173175
rect 289715 173147 289749 173175
rect 289777 173147 289811 173175
rect 289839 173147 289887 173175
rect 289577 173113 289887 173147
rect 289577 173085 289625 173113
rect 289653 173085 289687 173113
rect 289715 173085 289749 173113
rect 289777 173085 289811 173113
rect 289839 173085 289887 173113
rect 289577 173051 289887 173085
rect 289577 173023 289625 173051
rect 289653 173023 289687 173051
rect 289715 173023 289749 173051
rect 289777 173023 289811 173051
rect 289839 173023 289887 173051
rect 289577 172989 289887 173023
rect 289577 172961 289625 172989
rect 289653 172961 289687 172989
rect 289715 172961 289749 172989
rect 289777 172961 289811 172989
rect 289839 172961 289887 172989
rect 289577 164175 289887 172961
rect 289577 164147 289625 164175
rect 289653 164147 289687 164175
rect 289715 164147 289749 164175
rect 289777 164147 289811 164175
rect 289839 164147 289887 164175
rect 289577 164113 289887 164147
rect 289577 164085 289625 164113
rect 289653 164085 289687 164113
rect 289715 164085 289749 164113
rect 289777 164085 289811 164113
rect 289839 164085 289887 164113
rect 289577 164051 289887 164085
rect 289577 164023 289625 164051
rect 289653 164023 289687 164051
rect 289715 164023 289749 164051
rect 289777 164023 289811 164051
rect 289839 164023 289887 164051
rect 289577 163989 289887 164023
rect 289577 163961 289625 163989
rect 289653 163961 289687 163989
rect 289715 163961 289749 163989
rect 289777 163961 289811 163989
rect 289839 163961 289887 163989
rect 289577 155175 289887 163961
rect 289577 155147 289625 155175
rect 289653 155147 289687 155175
rect 289715 155147 289749 155175
rect 289777 155147 289811 155175
rect 289839 155147 289887 155175
rect 289577 155113 289887 155147
rect 289577 155085 289625 155113
rect 289653 155085 289687 155113
rect 289715 155085 289749 155113
rect 289777 155085 289811 155113
rect 289839 155085 289887 155113
rect 289577 155051 289887 155085
rect 289577 155023 289625 155051
rect 289653 155023 289687 155051
rect 289715 155023 289749 155051
rect 289777 155023 289811 155051
rect 289839 155023 289887 155051
rect 289577 154989 289887 155023
rect 289577 154961 289625 154989
rect 289653 154961 289687 154989
rect 289715 154961 289749 154989
rect 289777 154961 289811 154989
rect 289839 154961 289887 154989
rect 289577 146175 289887 154961
rect 289577 146147 289625 146175
rect 289653 146147 289687 146175
rect 289715 146147 289749 146175
rect 289777 146147 289811 146175
rect 289839 146147 289887 146175
rect 289577 146113 289887 146147
rect 289577 146085 289625 146113
rect 289653 146085 289687 146113
rect 289715 146085 289749 146113
rect 289777 146085 289811 146113
rect 289839 146085 289887 146113
rect 289577 146051 289887 146085
rect 289577 146023 289625 146051
rect 289653 146023 289687 146051
rect 289715 146023 289749 146051
rect 289777 146023 289811 146051
rect 289839 146023 289887 146051
rect 289577 145989 289887 146023
rect 289577 145961 289625 145989
rect 289653 145961 289687 145989
rect 289715 145961 289749 145989
rect 289777 145961 289811 145989
rect 289839 145961 289887 145989
rect 289577 137175 289887 145961
rect 289577 137147 289625 137175
rect 289653 137147 289687 137175
rect 289715 137147 289749 137175
rect 289777 137147 289811 137175
rect 289839 137147 289887 137175
rect 289577 137113 289887 137147
rect 289577 137085 289625 137113
rect 289653 137085 289687 137113
rect 289715 137085 289749 137113
rect 289777 137085 289811 137113
rect 289839 137085 289887 137113
rect 289577 137051 289887 137085
rect 289577 137023 289625 137051
rect 289653 137023 289687 137051
rect 289715 137023 289749 137051
rect 289777 137023 289811 137051
rect 289839 137023 289887 137051
rect 289577 136989 289887 137023
rect 289577 136961 289625 136989
rect 289653 136961 289687 136989
rect 289715 136961 289749 136989
rect 289777 136961 289811 136989
rect 289839 136961 289887 136989
rect 289577 128175 289887 136961
rect 289577 128147 289625 128175
rect 289653 128147 289687 128175
rect 289715 128147 289749 128175
rect 289777 128147 289811 128175
rect 289839 128147 289887 128175
rect 289577 128113 289887 128147
rect 289577 128085 289625 128113
rect 289653 128085 289687 128113
rect 289715 128085 289749 128113
rect 289777 128085 289811 128113
rect 289839 128085 289887 128113
rect 289577 128051 289887 128085
rect 289577 128023 289625 128051
rect 289653 128023 289687 128051
rect 289715 128023 289749 128051
rect 289777 128023 289811 128051
rect 289839 128023 289887 128051
rect 289577 127989 289887 128023
rect 289577 127961 289625 127989
rect 289653 127961 289687 127989
rect 289715 127961 289749 127989
rect 289777 127961 289811 127989
rect 289839 127961 289887 127989
rect 289577 119175 289887 127961
rect 289577 119147 289625 119175
rect 289653 119147 289687 119175
rect 289715 119147 289749 119175
rect 289777 119147 289811 119175
rect 289839 119147 289887 119175
rect 289577 119113 289887 119147
rect 289577 119085 289625 119113
rect 289653 119085 289687 119113
rect 289715 119085 289749 119113
rect 289777 119085 289811 119113
rect 289839 119085 289887 119113
rect 289577 119051 289887 119085
rect 289577 119023 289625 119051
rect 289653 119023 289687 119051
rect 289715 119023 289749 119051
rect 289777 119023 289811 119051
rect 289839 119023 289887 119051
rect 289577 118989 289887 119023
rect 289577 118961 289625 118989
rect 289653 118961 289687 118989
rect 289715 118961 289749 118989
rect 289777 118961 289811 118989
rect 289839 118961 289887 118989
rect 289577 110175 289887 118961
rect 289577 110147 289625 110175
rect 289653 110147 289687 110175
rect 289715 110147 289749 110175
rect 289777 110147 289811 110175
rect 289839 110147 289887 110175
rect 289577 110113 289887 110147
rect 289577 110085 289625 110113
rect 289653 110085 289687 110113
rect 289715 110085 289749 110113
rect 289777 110085 289811 110113
rect 289839 110085 289887 110113
rect 289577 110051 289887 110085
rect 289577 110023 289625 110051
rect 289653 110023 289687 110051
rect 289715 110023 289749 110051
rect 289777 110023 289811 110051
rect 289839 110023 289887 110051
rect 289577 109989 289887 110023
rect 289577 109961 289625 109989
rect 289653 109961 289687 109989
rect 289715 109961 289749 109989
rect 289777 109961 289811 109989
rect 289839 109961 289887 109989
rect 289577 101175 289887 109961
rect 289577 101147 289625 101175
rect 289653 101147 289687 101175
rect 289715 101147 289749 101175
rect 289777 101147 289811 101175
rect 289839 101147 289887 101175
rect 289577 101113 289887 101147
rect 289577 101085 289625 101113
rect 289653 101085 289687 101113
rect 289715 101085 289749 101113
rect 289777 101085 289811 101113
rect 289839 101085 289887 101113
rect 289577 101051 289887 101085
rect 289577 101023 289625 101051
rect 289653 101023 289687 101051
rect 289715 101023 289749 101051
rect 289777 101023 289811 101051
rect 289839 101023 289887 101051
rect 289577 100989 289887 101023
rect 289577 100961 289625 100989
rect 289653 100961 289687 100989
rect 289715 100961 289749 100989
rect 289777 100961 289811 100989
rect 289839 100961 289887 100989
rect 289577 92175 289887 100961
rect 289577 92147 289625 92175
rect 289653 92147 289687 92175
rect 289715 92147 289749 92175
rect 289777 92147 289811 92175
rect 289839 92147 289887 92175
rect 289577 92113 289887 92147
rect 289577 92085 289625 92113
rect 289653 92085 289687 92113
rect 289715 92085 289749 92113
rect 289777 92085 289811 92113
rect 289839 92085 289887 92113
rect 289577 92051 289887 92085
rect 289577 92023 289625 92051
rect 289653 92023 289687 92051
rect 289715 92023 289749 92051
rect 289777 92023 289811 92051
rect 289839 92023 289887 92051
rect 289577 91989 289887 92023
rect 289577 91961 289625 91989
rect 289653 91961 289687 91989
rect 289715 91961 289749 91989
rect 289777 91961 289811 91989
rect 289839 91961 289887 91989
rect 289577 83175 289887 91961
rect 289577 83147 289625 83175
rect 289653 83147 289687 83175
rect 289715 83147 289749 83175
rect 289777 83147 289811 83175
rect 289839 83147 289887 83175
rect 289577 83113 289887 83147
rect 289577 83085 289625 83113
rect 289653 83085 289687 83113
rect 289715 83085 289749 83113
rect 289777 83085 289811 83113
rect 289839 83085 289887 83113
rect 289577 83051 289887 83085
rect 289577 83023 289625 83051
rect 289653 83023 289687 83051
rect 289715 83023 289749 83051
rect 289777 83023 289811 83051
rect 289839 83023 289887 83051
rect 289577 82989 289887 83023
rect 289577 82961 289625 82989
rect 289653 82961 289687 82989
rect 289715 82961 289749 82989
rect 289777 82961 289811 82989
rect 289839 82961 289887 82989
rect 289577 74175 289887 82961
rect 289577 74147 289625 74175
rect 289653 74147 289687 74175
rect 289715 74147 289749 74175
rect 289777 74147 289811 74175
rect 289839 74147 289887 74175
rect 289577 74113 289887 74147
rect 289577 74085 289625 74113
rect 289653 74085 289687 74113
rect 289715 74085 289749 74113
rect 289777 74085 289811 74113
rect 289839 74085 289887 74113
rect 289577 74051 289887 74085
rect 289577 74023 289625 74051
rect 289653 74023 289687 74051
rect 289715 74023 289749 74051
rect 289777 74023 289811 74051
rect 289839 74023 289887 74051
rect 289577 73989 289887 74023
rect 289577 73961 289625 73989
rect 289653 73961 289687 73989
rect 289715 73961 289749 73989
rect 289777 73961 289811 73989
rect 289839 73961 289887 73989
rect 289577 65175 289887 73961
rect 289577 65147 289625 65175
rect 289653 65147 289687 65175
rect 289715 65147 289749 65175
rect 289777 65147 289811 65175
rect 289839 65147 289887 65175
rect 289577 65113 289887 65147
rect 289577 65085 289625 65113
rect 289653 65085 289687 65113
rect 289715 65085 289749 65113
rect 289777 65085 289811 65113
rect 289839 65085 289887 65113
rect 289577 65051 289887 65085
rect 289577 65023 289625 65051
rect 289653 65023 289687 65051
rect 289715 65023 289749 65051
rect 289777 65023 289811 65051
rect 289839 65023 289887 65051
rect 289577 64989 289887 65023
rect 289577 64961 289625 64989
rect 289653 64961 289687 64989
rect 289715 64961 289749 64989
rect 289777 64961 289811 64989
rect 289839 64961 289887 64989
rect 289577 56175 289887 64961
rect 289577 56147 289625 56175
rect 289653 56147 289687 56175
rect 289715 56147 289749 56175
rect 289777 56147 289811 56175
rect 289839 56147 289887 56175
rect 289577 56113 289887 56147
rect 289577 56085 289625 56113
rect 289653 56085 289687 56113
rect 289715 56085 289749 56113
rect 289777 56085 289811 56113
rect 289839 56085 289887 56113
rect 289577 56051 289887 56085
rect 289577 56023 289625 56051
rect 289653 56023 289687 56051
rect 289715 56023 289749 56051
rect 289777 56023 289811 56051
rect 289839 56023 289887 56051
rect 289577 55989 289887 56023
rect 289577 55961 289625 55989
rect 289653 55961 289687 55989
rect 289715 55961 289749 55989
rect 289777 55961 289811 55989
rect 289839 55961 289887 55989
rect 289577 47175 289887 55961
rect 289577 47147 289625 47175
rect 289653 47147 289687 47175
rect 289715 47147 289749 47175
rect 289777 47147 289811 47175
rect 289839 47147 289887 47175
rect 289577 47113 289887 47147
rect 289577 47085 289625 47113
rect 289653 47085 289687 47113
rect 289715 47085 289749 47113
rect 289777 47085 289811 47113
rect 289839 47085 289887 47113
rect 289577 47051 289887 47085
rect 289577 47023 289625 47051
rect 289653 47023 289687 47051
rect 289715 47023 289749 47051
rect 289777 47023 289811 47051
rect 289839 47023 289887 47051
rect 289577 46989 289887 47023
rect 289577 46961 289625 46989
rect 289653 46961 289687 46989
rect 289715 46961 289749 46989
rect 289777 46961 289811 46989
rect 289839 46961 289887 46989
rect 289577 38175 289887 46961
rect 289577 38147 289625 38175
rect 289653 38147 289687 38175
rect 289715 38147 289749 38175
rect 289777 38147 289811 38175
rect 289839 38147 289887 38175
rect 289577 38113 289887 38147
rect 289577 38085 289625 38113
rect 289653 38085 289687 38113
rect 289715 38085 289749 38113
rect 289777 38085 289811 38113
rect 289839 38085 289887 38113
rect 289577 38051 289887 38085
rect 289577 38023 289625 38051
rect 289653 38023 289687 38051
rect 289715 38023 289749 38051
rect 289777 38023 289811 38051
rect 289839 38023 289887 38051
rect 289577 37989 289887 38023
rect 289577 37961 289625 37989
rect 289653 37961 289687 37989
rect 289715 37961 289749 37989
rect 289777 37961 289811 37989
rect 289839 37961 289887 37989
rect 289577 29175 289887 37961
rect 289577 29147 289625 29175
rect 289653 29147 289687 29175
rect 289715 29147 289749 29175
rect 289777 29147 289811 29175
rect 289839 29147 289887 29175
rect 289577 29113 289887 29147
rect 289577 29085 289625 29113
rect 289653 29085 289687 29113
rect 289715 29085 289749 29113
rect 289777 29085 289811 29113
rect 289839 29085 289887 29113
rect 289577 29051 289887 29085
rect 289577 29023 289625 29051
rect 289653 29023 289687 29051
rect 289715 29023 289749 29051
rect 289777 29023 289811 29051
rect 289839 29023 289887 29051
rect 289577 28989 289887 29023
rect 289577 28961 289625 28989
rect 289653 28961 289687 28989
rect 289715 28961 289749 28989
rect 289777 28961 289811 28989
rect 289839 28961 289887 28989
rect 289577 20175 289887 28961
rect 289577 20147 289625 20175
rect 289653 20147 289687 20175
rect 289715 20147 289749 20175
rect 289777 20147 289811 20175
rect 289839 20147 289887 20175
rect 289577 20113 289887 20147
rect 289577 20085 289625 20113
rect 289653 20085 289687 20113
rect 289715 20085 289749 20113
rect 289777 20085 289811 20113
rect 289839 20085 289887 20113
rect 289577 20051 289887 20085
rect 289577 20023 289625 20051
rect 289653 20023 289687 20051
rect 289715 20023 289749 20051
rect 289777 20023 289811 20051
rect 289839 20023 289887 20051
rect 289577 19989 289887 20023
rect 289577 19961 289625 19989
rect 289653 19961 289687 19989
rect 289715 19961 289749 19989
rect 289777 19961 289811 19989
rect 289839 19961 289887 19989
rect 289577 11175 289887 19961
rect 289577 11147 289625 11175
rect 289653 11147 289687 11175
rect 289715 11147 289749 11175
rect 289777 11147 289811 11175
rect 289839 11147 289887 11175
rect 289577 11113 289887 11147
rect 289577 11085 289625 11113
rect 289653 11085 289687 11113
rect 289715 11085 289749 11113
rect 289777 11085 289811 11113
rect 289839 11085 289887 11113
rect 289577 11051 289887 11085
rect 289577 11023 289625 11051
rect 289653 11023 289687 11051
rect 289715 11023 289749 11051
rect 289777 11023 289811 11051
rect 289839 11023 289887 11051
rect 289577 10989 289887 11023
rect 289577 10961 289625 10989
rect 289653 10961 289687 10989
rect 289715 10961 289749 10989
rect 289777 10961 289811 10989
rect 289839 10961 289887 10989
rect 289577 2175 289887 10961
rect 289577 2147 289625 2175
rect 289653 2147 289687 2175
rect 289715 2147 289749 2175
rect 289777 2147 289811 2175
rect 289839 2147 289887 2175
rect 289577 2113 289887 2147
rect 289577 2085 289625 2113
rect 289653 2085 289687 2113
rect 289715 2085 289749 2113
rect 289777 2085 289811 2113
rect 289839 2085 289887 2113
rect 289577 2051 289887 2085
rect 289577 2023 289625 2051
rect 289653 2023 289687 2051
rect 289715 2023 289749 2051
rect 289777 2023 289811 2051
rect 289839 2023 289887 2051
rect 289577 1989 289887 2023
rect 289577 1961 289625 1989
rect 289653 1961 289687 1989
rect 289715 1961 289749 1989
rect 289777 1961 289811 1989
rect 289839 1961 289887 1989
rect 289577 -80 289887 1961
rect 289577 -108 289625 -80
rect 289653 -108 289687 -80
rect 289715 -108 289749 -80
rect 289777 -108 289811 -80
rect 289839 -108 289887 -80
rect 289577 -142 289887 -108
rect 289577 -170 289625 -142
rect 289653 -170 289687 -142
rect 289715 -170 289749 -142
rect 289777 -170 289811 -142
rect 289839 -170 289887 -142
rect 289577 -204 289887 -170
rect 289577 -232 289625 -204
rect 289653 -232 289687 -204
rect 289715 -232 289749 -204
rect 289777 -232 289811 -204
rect 289839 -232 289887 -204
rect 289577 -266 289887 -232
rect 289577 -294 289625 -266
rect 289653 -294 289687 -266
rect 289715 -294 289749 -266
rect 289777 -294 289811 -266
rect 289839 -294 289887 -266
rect 289577 -822 289887 -294
rect 291437 299086 291747 299134
rect 291437 299058 291485 299086
rect 291513 299058 291547 299086
rect 291575 299058 291609 299086
rect 291637 299058 291671 299086
rect 291699 299058 291747 299086
rect 291437 299024 291747 299058
rect 291437 298996 291485 299024
rect 291513 298996 291547 299024
rect 291575 298996 291609 299024
rect 291637 298996 291671 299024
rect 291699 298996 291747 299024
rect 291437 298962 291747 298996
rect 291437 298934 291485 298962
rect 291513 298934 291547 298962
rect 291575 298934 291609 298962
rect 291637 298934 291671 298962
rect 291699 298934 291747 298962
rect 291437 298900 291747 298934
rect 291437 298872 291485 298900
rect 291513 298872 291547 298900
rect 291575 298872 291609 298900
rect 291637 298872 291671 298900
rect 291699 298872 291747 298900
rect 291437 293175 291747 298872
rect 298680 299086 298990 299134
rect 298680 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect 298680 299024 298990 299058
rect 298680 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect 298680 298962 298990 298996
rect 298680 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect 298680 298900 298990 298934
rect 298680 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect 291437 293147 291485 293175
rect 291513 293147 291547 293175
rect 291575 293147 291609 293175
rect 291637 293147 291671 293175
rect 291699 293147 291747 293175
rect 291437 293113 291747 293147
rect 291437 293085 291485 293113
rect 291513 293085 291547 293113
rect 291575 293085 291609 293113
rect 291637 293085 291671 293113
rect 291699 293085 291747 293113
rect 291437 293051 291747 293085
rect 291437 293023 291485 293051
rect 291513 293023 291547 293051
rect 291575 293023 291609 293051
rect 291637 293023 291671 293051
rect 291699 293023 291747 293051
rect 291437 292989 291747 293023
rect 291437 292961 291485 292989
rect 291513 292961 291547 292989
rect 291575 292961 291609 292989
rect 291637 292961 291671 292989
rect 291699 292961 291747 292989
rect 291437 284175 291747 292961
rect 291437 284147 291485 284175
rect 291513 284147 291547 284175
rect 291575 284147 291609 284175
rect 291637 284147 291671 284175
rect 291699 284147 291747 284175
rect 291437 284113 291747 284147
rect 291437 284085 291485 284113
rect 291513 284085 291547 284113
rect 291575 284085 291609 284113
rect 291637 284085 291671 284113
rect 291699 284085 291747 284113
rect 291437 284051 291747 284085
rect 291437 284023 291485 284051
rect 291513 284023 291547 284051
rect 291575 284023 291609 284051
rect 291637 284023 291671 284051
rect 291699 284023 291747 284051
rect 291437 283989 291747 284023
rect 291437 283961 291485 283989
rect 291513 283961 291547 283989
rect 291575 283961 291609 283989
rect 291637 283961 291671 283989
rect 291699 283961 291747 283989
rect 291437 275175 291747 283961
rect 291437 275147 291485 275175
rect 291513 275147 291547 275175
rect 291575 275147 291609 275175
rect 291637 275147 291671 275175
rect 291699 275147 291747 275175
rect 291437 275113 291747 275147
rect 291437 275085 291485 275113
rect 291513 275085 291547 275113
rect 291575 275085 291609 275113
rect 291637 275085 291671 275113
rect 291699 275085 291747 275113
rect 291437 275051 291747 275085
rect 291437 275023 291485 275051
rect 291513 275023 291547 275051
rect 291575 275023 291609 275051
rect 291637 275023 291671 275051
rect 291699 275023 291747 275051
rect 291437 274989 291747 275023
rect 291437 274961 291485 274989
rect 291513 274961 291547 274989
rect 291575 274961 291609 274989
rect 291637 274961 291671 274989
rect 291699 274961 291747 274989
rect 291437 266175 291747 274961
rect 291437 266147 291485 266175
rect 291513 266147 291547 266175
rect 291575 266147 291609 266175
rect 291637 266147 291671 266175
rect 291699 266147 291747 266175
rect 291437 266113 291747 266147
rect 291437 266085 291485 266113
rect 291513 266085 291547 266113
rect 291575 266085 291609 266113
rect 291637 266085 291671 266113
rect 291699 266085 291747 266113
rect 291437 266051 291747 266085
rect 291437 266023 291485 266051
rect 291513 266023 291547 266051
rect 291575 266023 291609 266051
rect 291637 266023 291671 266051
rect 291699 266023 291747 266051
rect 291437 265989 291747 266023
rect 291437 265961 291485 265989
rect 291513 265961 291547 265989
rect 291575 265961 291609 265989
rect 291637 265961 291671 265989
rect 291699 265961 291747 265989
rect 291437 257175 291747 265961
rect 291437 257147 291485 257175
rect 291513 257147 291547 257175
rect 291575 257147 291609 257175
rect 291637 257147 291671 257175
rect 291699 257147 291747 257175
rect 291437 257113 291747 257147
rect 291437 257085 291485 257113
rect 291513 257085 291547 257113
rect 291575 257085 291609 257113
rect 291637 257085 291671 257113
rect 291699 257085 291747 257113
rect 291437 257051 291747 257085
rect 291437 257023 291485 257051
rect 291513 257023 291547 257051
rect 291575 257023 291609 257051
rect 291637 257023 291671 257051
rect 291699 257023 291747 257051
rect 291437 256989 291747 257023
rect 291437 256961 291485 256989
rect 291513 256961 291547 256989
rect 291575 256961 291609 256989
rect 291637 256961 291671 256989
rect 291699 256961 291747 256989
rect 291437 248175 291747 256961
rect 291437 248147 291485 248175
rect 291513 248147 291547 248175
rect 291575 248147 291609 248175
rect 291637 248147 291671 248175
rect 291699 248147 291747 248175
rect 291437 248113 291747 248147
rect 291437 248085 291485 248113
rect 291513 248085 291547 248113
rect 291575 248085 291609 248113
rect 291637 248085 291671 248113
rect 291699 248085 291747 248113
rect 291437 248051 291747 248085
rect 291437 248023 291485 248051
rect 291513 248023 291547 248051
rect 291575 248023 291609 248051
rect 291637 248023 291671 248051
rect 291699 248023 291747 248051
rect 291437 247989 291747 248023
rect 291437 247961 291485 247989
rect 291513 247961 291547 247989
rect 291575 247961 291609 247989
rect 291637 247961 291671 247989
rect 291699 247961 291747 247989
rect 291437 239175 291747 247961
rect 291437 239147 291485 239175
rect 291513 239147 291547 239175
rect 291575 239147 291609 239175
rect 291637 239147 291671 239175
rect 291699 239147 291747 239175
rect 291437 239113 291747 239147
rect 291437 239085 291485 239113
rect 291513 239085 291547 239113
rect 291575 239085 291609 239113
rect 291637 239085 291671 239113
rect 291699 239085 291747 239113
rect 291437 239051 291747 239085
rect 291437 239023 291485 239051
rect 291513 239023 291547 239051
rect 291575 239023 291609 239051
rect 291637 239023 291671 239051
rect 291699 239023 291747 239051
rect 291437 238989 291747 239023
rect 291437 238961 291485 238989
rect 291513 238961 291547 238989
rect 291575 238961 291609 238989
rect 291637 238961 291671 238989
rect 291699 238961 291747 238989
rect 291437 230175 291747 238961
rect 291437 230147 291485 230175
rect 291513 230147 291547 230175
rect 291575 230147 291609 230175
rect 291637 230147 291671 230175
rect 291699 230147 291747 230175
rect 291437 230113 291747 230147
rect 291437 230085 291485 230113
rect 291513 230085 291547 230113
rect 291575 230085 291609 230113
rect 291637 230085 291671 230113
rect 291699 230085 291747 230113
rect 291437 230051 291747 230085
rect 291437 230023 291485 230051
rect 291513 230023 291547 230051
rect 291575 230023 291609 230051
rect 291637 230023 291671 230051
rect 291699 230023 291747 230051
rect 291437 229989 291747 230023
rect 291437 229961 291485 229989
rect 291513 229961 291547 229989
rect 291575 229961 291609 229989
rect 291637 229961 291671 229989
rect 291699 229961 291747 229989
rect 291437 221175 291747 229961
rect 291437 221147 291485 221175
rect 291513 221147 291547 221175
rect 291575 221147 291609 221175
rect 291637 221147 291671 221175
rect 291699 221147 291747 221175
rect 291437 221113 291747 221147
rect 291437 221085 291485 221113
rect 291513 221085 291547 221113
rect 291575 221085 291609 221113
rect 291637 221085 291671 221113
rect 291699 221085 291747 221113
rect 291437 221051 291747 221085
rect 291437 221023 291485 221051
rect 291513 221023 291547 221051
rect 291575 221023 291609 221051
rect 291637 221023 291671 221051
rect 291699 221023 291747 221051
rect 291437 220989 291747 221023
rect 291437 220961 291485 220989
rect 291513 220961 291547 220989
rect 291575 220961 291609 220989
rect 291637 220961 291671 220989
rect 291699 220961 291747 220989
rect 291437 212175 291747 220961
rect 291437 212147 291485 212175
rect 291513 212147 291547 212175
rect 291575 212147 291609 212175
rect 291637 212147 291671 212175
rect 291699 212147 291747 212175
rect 291437 212113 291747 212147
rect 291437 212085 291485 212113
rect 291513 212085 291547 212113
rect 291575 212085 291609 212113
rect 291637 212085 291671 212113
rect 291699 212085 291747 212113
rect 291437 212051 291747 212085
rect 291437 212023 291485 212051
rect 291513 212023 291547 212051
rect 291575 212023 291609 212051
rect 291637 212023 291671 212051
rect 291699 212023 291747 212051
rect 291437 211989 291747 212023
rect 291437 211961 291485 211989
rect 291513 211961 291547 211989
rect 291575 211961 291609 211989
rect 291637 211961 291671 211989
rect 291699 211961 291747 211989
rect 291437 203175 291747 211961
rect 291437 203147 291485 203175
rect 291513 203147 291547 203175
rect 291575 203147 291609 203175
rect 291637 203147 291671 203175
rect 291699 203147 291747 203175
rect 291437 203113 291747 203147
rect 291437 203085 291485 203113
rect 291513 203085 291547 203113
rect 291575 203085 291609 203113
rect 291637 203085 291671 203113
rect 291699 203085 291747 203113
rect 291437 203051 291747 203085
rect 291437 203023 291485 203051
rect 291513 203023 291547 203051
rect 291575 203023 291609 203051
rect 291637 203023 291671 203051
rect 291699 203023 291747 203051
rect 291437 202989 291747 203023
rect 291437 202961 291485 202989
rect 291513 202961 291547 202989
rect 291575 202961 291609 202989
rect 291637 202961 291671 202989
rect 291699 202961 291747 202989
rect 291437 194175 291747 202961
rect 291437 194147 291485 194175
rect 291513 194147 291547 194175
rect 291575 194147 291609 194175
rect 291637 194147 291671 194175
rect 291699 194147 291747 194175
rect 291437 194113 291747 194147
rect 291437 194085 291485 194113
rect 291513 194085 291547 194113
rect 291575 194085 291609 194113
rect 291637 194085 291671 194113
rect 291699 194085 291747 194113
rect 291437 194051 291747 194085
rect 291437 194023 291485 194051
rect 291513 194023 291547 194051
rect 291575 194023 291609 194051
rect 291637 194023 291671 194051
rect 291699 194023 291747 194051
rect 291437 193989 291747 194023
rect 291437 193961 291485 193989
rect 291513 193961 291547 193989
rect 291575 193961 291609 193989
rect 291637 193961 291671 193989
rect 291699 193961 291747 193989
rect 291437 185175 291747 193961
rect 291437 185147 291485 185175
rect 291513 185147 291547 185175
rect 291575 185147 291609 185175
rect 291637 185147 291671 185175
rect 291699 185147 291747 185175
rect 291437 185113 291747 185147
rect 291437 185085 291485 185113
rect 291513 185085 291547 185113
rect 291575 185085 291609 185113
rect 291637 185085 291671 185113
rect 291699 185085 291747 185113
rect 291437 185051 291747 185085
rect 291437 185023 291485 185051
rect 291513 185023 291547 185051
rect 291575 185023 291609 185051
rect 291637 185023 291671 185051
rect 291699 185023 291747 185051
rect 291437 184989 291747 185023
rect 291437 184961 291485 184989
rect 291513 184961 291547 184989
rect 291575 184961 291609 184989
rect 291637 184961 291671 184989
rect 291699 184961 291747 184989
rect 291437 176175 291747 184961
rect 291437 176147 291485 176175
rect 291513 176147 291547 176175
rect 291575 176147 291609 176175
rect 291637 176147 291671 176175
rect 291699 176147 291747 176175
rect 291437 176113 291747 176147
rect 291437 176085 291485 176113
rect 291513 176085 291547 176113
rect 291575 176085 291609 176113
rect 291637 176085 291671 176113
rect 291699 176085 291747 176113
rect 291437 176051 291747 176085
rect 291437 176023 291485 176051
rect 291513 176023 291547 176051
rect 291575 176023 291609 176051
rect 291637 176023 291671 176051
rect 291699 176023 291747 176051
rect 291437 175989 291747 176023
rect 291437 175961 291485 175989
rect 291513 175961 291547 175989
rect 291575 175961 291609 175989
rect 291637 175961 291671 175989
rect 291699 175961 291747 175989
rect 291437 167175 291747 175961
rect 291437 167147 291485 167175
rect 291513 167147 291547 167175
rect 291575 167147 291609 167175
rect 291637 167147 291671 167175
rect 291699 167147 291747 167175
rect 291437 167113 291747 167147
rect 291437 167085 291485 167113
rect 291513 167085 291547 167113
rect 291575 167085 291609 167113
rect 291637 167085 291671 167113
rect 291699 167085 291747 167113
rect 291437 167051 291747 167085
rect 291437 167023 291485 167051
rect 291513 167023 291547 167051
rect 291575 167023 291609 167051
rect 291637 167023 291671 167051
rect 291699 167023 291747 167051
rect 291437 166989 291747 167023
rect 291437 166961 291485 166989
rect 291513 166961 291547 166989
rect 291575 166961 291609 166989
rect 291637 166961 291671 166989
rect 291699 166961 291747 166989
rect 291437 158175 291747 166961
rect 291437 158147 291485 158175
rect 291513 158147 291547 158175
rect 291575 158147 291609 158175
rect 291637 158147 291671 158175
rect 291699 158147 291747 158175
rect 291437 158113 291747 158147
rect 291437 158085 291485 158113
rect 291513 158085 291547 158113
rect 291575 158085 291609 158113
rect 291637 158085 291671 158113
rect 291699 158085 291747 158113
rect 291437 158051 291747 158085
rect 291437 158023 291485 158051
rect 291513 158023 291547 158051
rect 291575 158023 291609 158051
rect 291637 158023 291671 158051
rect 291699 158023 291747 158051
rect 291437 157989 291747 158023
rect 291437 157961 291485 157989
rect 291513 157961 291547 157989
rect 291575 157961 291609 157989
rect 291637 157961 291671 157989
rect 291699 157961 291747 157989
rect 291437 149175 291747 157961
rect 291437 149147 291485 149175
rect 291513 149147 291547 149175
rect 291575 149147 291609 149175
rect 291637 149147 291671 149175
rect 291699 149147 291747 149175
rect 291437 149113 291747 149147
rect 291437 149085 291485 149113
rect 291513 149085 291547 149113
rect 291575 149085 291609 149113
rect 291637 149085 291671 149113
rect 291699 149085 291747 149113
rect 291437 149051 291747 149085
rect 291437 149023 291485 149051
rect 291513 149023 291547 149051
rect 291575 149023 291609 149051
rect 291637 149023 291671 149051
rect 291699 149023 291747 149051
rect 291437 148989 291747 149023
rect 291437 148961 291485 148989
rect 291513 148961 291547 148989
rect 291575 148961 291609 148989
rect 291637 148961 291671 148989
rect 291699 148961 291747 148989
rect 291437 140175 291747 148961
rect 291437 140147 291485 140175
rect 291513 140147 291547 140175
rect 291575 140147 291609 140175
rect 291637 140147 291671 140175
rect 291699 140147 291747 140175
rect 291437 140113 291747 140147
rect 291437 140085 291485 140113
rect 291513 140085 291547 140113
rect 291575 140085 291609 140113
rect 291637 140085 291671 140113
rect 291699 140085 291747 140113
rect 291437 140051 291747 140085
rect 291437 140023 291485 140051
rect 291513 140023 291547 140051
rect 291575 140023 291609 140051
rect 291637 140023 291671 140051
rect 291699 140023 291747 140051
rect 291437 139989 291747 140023
rect 291437 139961 291485 139989
rect 291513 139961 291547 139989
rect 291575 139961 291609 139989
rect 291637 139961 291671 139989
rect 291699 139961 291747 139989
rect 291437 131175 291747 139961
rect 291437 131147 291485 131175
rect 291513 131147 291547 131175
rect 291575 131147 291609 131175
rect 291637 131147 291671 131175
rect 291699 131147 291747 131175
rect 291437 131113 291747 131147
rect 291437 131085 291485 131113
rect 291513 131085 291547 131113
rect 291575 131085 291609 131113
rect 291637 131085 291671 131113
rect 291699 131085 291747 131113
rect 291437 131051 291747 131085
rect 291437 131023 291485 131051
rect 291513 131023 291547 131051
rect 291575 131023 291609 131051
rect 291637 131023 291671 131051
rect 291699 131023 291747 131051
rect 291437 130989 291747 131023
rect 291437 130961 291485 130989
rect 291513 130961 291547 130989
rect 291575 130961 291609 130989
rect 291637 130961 291671 130989
rect 291699 130961 291747 130989
rect 291437 122175 291747 130961
rect 291437 122147 291485 122175
rect 291513 122147 291547 122175
rect 291575 122147 291609 122175
rect 291637 122147 291671 122175
rect 291699 122147 291747 122175
rect 291437 122113 291747 122147
rect 291437 122085 291485 122113
rect 291513 122085 291547 122113
rect 291575 122085 291609 122113
rect 291637 122085 291671 122113
rect 291699 122085 291747 122113
rect 291437 122051 291747 122085
rect 291437 122023 291485 122051
rect 291513 122023 291547 122051
rect 291575 122023 291609 122051
rect 291637 122023 291671 122051
rect 291699 122023 291747 122051
rect 291437 121989 291747 122023
rect 291437 121961 291485 121989
rect 291513 121961 291547 121989
rect 291575 121961 291609 121989
rect 291637 121961 291671 121989
rect 291699 121961 291747 121989
rect 291437 113175 291747 121961
rect 291437 113147 291485 113175
rect 291513 113147 291547 113175
rect 291575 113147 291609 113175
rect 291637 113147 291671 113175
rect 291699 113147 291747 113175
rect 291437 113113 291747 113147
rect 291437 113085 291485 113113
rect 291513 113085 291547 113113
rect 291575 113085 291609 113113
rect 291637 113085 291671 113113
rect 291699 113085 291747 113113
rect 291437 113051 291747 113085
rect 291437 113023 291485 113051
rect 291513 113023 291547 113051
rect 291575 113023 291609 113051
rect 291637 113023 291671 113051
rect 291699 113023 291747 113051
rect 291437 112989 291747 113023
rect 291437 112961 291485 112989
rect 291513 112961 291547 112989
rect 291575 112961 291609 112989
rect 291637 112961 291671 112989
rect 291699 112961 291747 112989
rect 291437 104175 291747 112961
rect 291437 104147 291485 104175
rect 291513 104147 291547 104175
rect 291575 104147 291609 104175
rect 291637 104147 291671 104175
rect 291699 104147 291747 104175
rect 291437 104113 291747 104147
rect 291437 104085 291485 104113
rect 291513 104085 291547 104113
rect 291575 104085 291609 104113
rect 291637 104085 291671 104113
rect 291699 104085 291747 104113
rect 291437 104051 291747 104085
rect 291437 104023 291485 104051
rect 291513 104023 291547 104051
rect 291575 104023 291609 104051
rect 291637 104023 291671 104051
rect 291699 104023 291747 104051
rect 291437 103989 291747 104023
rect 291437 103961 291485 103989
rect 291513 103961 291547 103989
rect 291575 103961 291609 103989
rect 291637 103961 291671 103989
rect 291699 103961 291747 103989
rect 291437 95175 291747 103961
rect 291437 95147 291485 95175
rect 291513 95147 291547 95175
rect 291575 95147 291609 95175
rect 291637 95147 291671 95175
rect 291699 95147 291747 95175
rect 291437 95113 291747 95147
rect 291437 95085 291485 95113
rect 291513 95085 291547 95113
rect 291575 95085 291609 95113
rect 291637 95085 291671 95113
rect 291699 95085 291747 95113
rect 291437 95051 291747 95085
rect 291437 95023 291485 95051
rect 291513 95023 291547 95051
rect 291575 95023 291609 95051
rect 291637 95023 291671 95051
rect 291699 95023 291747 95051
rect 291437 94989 291747 95023
rect 291437 94961 291485 94989
rect 291513 94961 291547 94989
rect 291575 94961 291609 94989
rect 291637 94961 291671 94989
rect 291699 94961 291747 94989
rect 291437 86175 291747 94961
rect 291437 86147 291485 86175
rect 291513 86147 291547 86175
rect 291575 86147 291609 86175
rect 291637 86147 291671 86175
rect 291699 86147 291747 86175
rect 291437 86113 291747 86147
rect 291437 86085 291485 86113
rect 291513 86085 291547 86113
rect 291575 86085 291609 86113
rect 291637 86085 291671 86113
rect 291699 86085 291747 86113
rect 291437 86051 291747 86085
rect 291437 86023 291485 86051
rect 291513 86023 291547 86051
rect 291575 86023 291609 86051
rect 291637 86023 291671 86051
rect 291699 86023 291747 86051
rect 291437 85989 291747 86023
rect 291437 85961 291485 85989
rect 291513 85961 291547 85989
rect 291575 85961 291609 85989
rect 291637 85961 291671 85989
rect 291699 85961 291747 85989
rect 291437 77175 291747 85961
rect 291437 77147 291485 77175
rect 291513 77147 291547 77175
rect 291575 77147 291609 77175
rect 291637 77147 291671 77175
rect 291699 77147 291747 77175
rect 291437 77113 291747 77147
rect 291437 77085 291485 77113
rect 291513 77085 291547 77113
rect 291575 77085 291609 77113
rect 291637 77085 291671 77113
rect 291699 77085 291747 77113
rect 291437 77051 291747 77085
rect 291437 77023 291485 77051
rect 291513 77023 291547 77051
rect 291575 77023 291609 77051
rect 291637 77023 291671 77051
rect 291699 77023 291747 77051
rect 291437 76989 291747 77023
rect 291437 76961 291485 76989
rect 291513 76961 291547 76989
rect 291575 76961 291609 76989
rect 291637 76961 291671 76989
rect 291699 76961 291747 76989
rect 291437 68175 291747 76961
rect 291437 68147 291485 68175
rect 291513 68147 291547 68175
rect 291575 68147 291609 68175
rect 291637 68147 291671 68175
rect 291699 68147 291747 68175
rect 291437 68113 291747 68147
rect 291437 68085 291485 68113
rect 291513 68085 291547 68113
rect 291575 68085 291609 68113
rect 291637 68085 291671 68113
rect 291699 68085 291747 68113
rect 291437 68051 291747 68085
rect 291437 68023 291485 68051
rect 291513 68023 291547 68051
rect 291575 68023 291609 68051
rect 291637 68023 291671 68051
rect 291699 68023 291747 68051
rect 291437 67989 291747 68023
rect 291437 67961 291485 67989
rect 291513 67961 291547 67989
rect 291575 67961 291609 67989
rect 291637 67961 291671 67989
rect 291699 67961 291747 67989
rect 291437 59175 291747 67961
rect 291437 59147 291485 59175
rect 291513 59147 291547 59175
rect 291575 59147 291609 59175
rect 291637 59147 291671 59175
rect 291699 59147 291747 59175
rect 291437 59113 291747 59147
rect 291437 59085 291485 59113
rect 291513 59085 291547 59113
rect 291575 59085 291609 59113
rect 291637 59085 291671 59113
rect 291699 59085 291747 59113
rect 291437 59051 291747 59085
rect 291437 59023 291485 59051
rect 291513 59023 291547 59051
rect 291575 59023 291609 59051
rect 291637 59023 291671 59051
rect 291699 59023 291747 59051
rect 291437 58989 291747 59023
rect 291437 58961 291485 58989
rect 291513 58961 291547 58989
rect 291575 58961 291609 58989
rect 291637 58961 291671 58989
rect 291699 58961 291747 58989
rect 291437 50175 291747 58961
rect 291437 50147 291485 50175
rect 291513 50147 291547 50175
rect 291575 50147 291609 50175
rect 291637 50147 291671 50175
rect 291699 50147 291747 50175
rect 291437 50113 291747 50147
rect 291437 50085 291485 50113
rect 291513 50085 291547 50113
rect 291575 50085 291609 50113
rect 291637 50085 291671 50113
rect 291699 50085 291747 50113
rect 291437 50051 291747 50085
rect 291437 50023 291485 50051
rect 291513 50023 291547 50051
rect 291575 50023 291609 50051
rect 291637 50023 291671 50051
rect 291699 50023 291747 50051
rect 291437 49989 291747 50023
rect 291437 49961 291485 49989
rect 291513 49961 291547 49989
rect 291575 49961 291609 49989
rect 291637 49961 291671 49989
rect 291699 49961 291747 49989
rect 291437 41175 291747 49961
rect 291437 41147 291485 41175
rect 291513 41147 291547 41175
rect 291575 41147 291609 41175
rect 291637 41147 291671 41175
rect 291699 41147 291747 41175
rect 291437 41113 291747 41147
rect 291437 41085 291485 41113
rect 291513 41085 291547 41113
rect 291575 41085 291609 41113
rect 291637 41085 291671 41113
rect 291699 41085 291747 41113
rect 291437 41051 291747 41085
rect 291437 41023 291485 41051
rect 291513 41023 291547 41051
rect 291575 41023 291609 41051
rect 291637 41023 291671 41051
rect 291699 41023 291747 41051
rect 291437 40989 291747 41023
rect 291437 40961 291485 40989
rect 291513 40961 291547 40989
rect 291575 40961 291609 40989
rect 291637 40961 291671 40989
rect 291699 40961 291747 40989
rect 291437 32175 291747 40961
rect 291437 32147 291485 32175
rect 291513 32147 291547 32175
rect 291575 32147 291609 32175
rect 291637 32147 291671 32175
rect 291699 32147 291747 32175
rect 291437 32113 291747 32147
rect 291437 32085 291485 32113
rect 291513 32085 291547 32113
rect 291575 32085 291609 32113
rect 291637 32085 291671 32113
rect 291699 32085 291747 32113
rect 291437 32051 291747 32085
rect 291437 32023 291485 32051
rect 291513 32023 291547 32051
rect 291575 32023 291609 32051
rect 291637 32023 291671 32051
rect 291699 32023 291747 32051
rect 291437 31989 291747 32023
rect 291437 31961 291485 31989
rect 291513 31961 291547 31989
rect 291575 31961 291609 31989
rect 291637 31961 291671 31989
rect 291699 31961 291747 31989
rect 291437 23175 291747 31961
rect 291437 23147 291485 23175
rect 291513 23147 291547 23175
rect 291575 23147 291609 23175
rect 291637 23147 291671 23175
rect 291699 23147 291747 23175
rect 291437 23113 291747 23147
rect 291437 23085 291485 23113
rect 291513 23085 291547 23113
rect 291575 23085 291609 23113
rect 291637 23085 291671 23113
rect 291699 23085 291747 23113
rect 291437 23051 291747 23085
rect 291437 23023 291485 23051
rect 291513 23023 291547 23051
rect 291575 23023 291609 23051
rect 291637 23023 291671 23051
rect 291699 23023 291747 23051
rect 291437 22989 291747 23023
rect 291437 22961 291485 22989
rect 291513 22961 291547 22989
rect 291575 22961 291609 22989
rect 291637 22961 291671 22989
rect 291699 22961 291747 22989
rect 291437 14175 291747 22961
rect 291437 14147 291485 14175
rect 291513 14147 291547 14175
rect 291575 14147 291609 14175
rect 291637 14147 291671 14175
rect 291699 14147 291747 14175
rect 291437 14113 291747 14147
rect 291437 14085 291485 14113
rect 291513 14085 291547 14113
rect 291575 14085 291609 14113
rect 291637 14085 291671 14113
rect 291699 14085 291747 14113
rect 291437 14051 291747 14085
rect 291437 14023 291485 14051
rect 291513 14023 291547 14051
rect 291575 14023 291609 14051
rect 291637 14023 291671 14051
rect 291699 14023 291747 14051
rect 291437 13989 291747 14023
rect 291437 13961 291485 13989
rect 291513 13961 291547 13989
rect 291575 13961 291609 13989
rect 291637 13961 291671 13989
rect 291699 13961 291747 13989
rect 291437 5175 291747 13961
rect 291437 5147 291485 5175
rect 291513 5147 291547 5175
rect 291575 5147 291609 5175
rect 291637 5147 291671 5175
rect 291699 5147 291747 5175
rect 291437 5113 291747 5147
rect 291437 5085 291485 5113
rect 291513 5085 291547 5113
rect 291575 5085 291609 5113
rect 291637 5085 291671 5113
rect 291699 5085 291747 5113
rect 291437 5051 291747 5085
rect 291437 5023 291485 5051
rect 291513 5023 291547 5051
rect 291575 5023 291609 5051
rect 291637 5023 291671 5051
rect 291699 5023 291747 5051
rect 291437 4989 291747 5023
rect 291437 4961 291485 4989
rect 291513 4961 291547 4989
rect 291575 4961 291609 4989
rect 291637 4961 291671 4989
rect 291699 4961 291747 4989
rect 291437 -560 291747 4961
rect 298200 298606 298510 298654
rect 298200 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect 298200 298544 298510 298578
rect 298200 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect 298200 298482 298510 298516
rect 298200 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect 298200 298420 298510 298454
rect 298200 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect 298200 290175 298510 298392
rect 298200 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298510 290175
rect 298200 290113 298510 290147
rect 298200 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298510 290113
rect 298200 290051 298510 290085
rect 298200 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298510 290051
rect 298200 289989 298510 290023
rect 298200 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298510 289989
rect 298200 281175 298510 289961
rect 298200 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298510 281175
rect 298200 281113 298510 281147
rect 298200 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298510 281113
rect 298200 281051 298510 281085
rect 298200 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298510 281051
rect 298200 280989 298510 281023
rect 298200 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298510 280989
rect 298200 272175 298510 280961
rect 298200 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298510 272175
rect 298200 272113 298510 272147
rect 298200 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298510 272113
rect 298200 272051 298510 272085
rect 298200 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298510 272051
rect 298200 271989 298510 272023
rect 298200 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298510 271989
rect 298200 263175 298510 271961
rect 298200 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298510 263175
rect 298200 263113 298510 263147
rect 298200 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298510 263113
rect 298200 263051 298510 263085
rect 298200 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298510 263051
rect 298200 262989 298510 263023
rect 298200 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298510 262989
rect 298200 254175 298510 262961
rect 298200 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298510 254175
rect 298200 254113 298510 254147
rect 298200 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298510 254113
rect 298200 254051 298510 254085
rect 298200 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298510 254051
rect 298200 253989 298510 254023
rect 298200 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298510 253989
rect 298200 245175 298510 253961
rect 298200 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298510 245175
rect 298200 245113 298510 245147
rect 298200 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298510 245113
rect 298200 245051 298510 245085
rect 298200 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298510 245051
rect 298200 244989 298510 245023
rect 298200 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298510 244989
rect 298200 236175 298510 244961
rect 298200 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298510 236175
rect 298200 236113 298510 236147
rect 298200 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298510 236113
rect 298200 236051 298510 236085
rect 298200 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298510 236051
rect 298200 235989 298510 236023
rect 298200 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298510 235989
rect 298200 227175 298510 235961
rect 298200 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298510 227175
rect 298200 227113 298510 227147
rect 298200 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298510 227113
rect 298200 227051 298510 227085
rect 298200 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298510 227051
rect 298200 226989 298510 227023
rect 298200 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298510 226989
rect 298200 218175 298510 226961
rect 298200 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298510 218175
rect 298200 218113 298510 218147
rect 298200 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298510 218113
rect 298200 218051 298510 218085
rect 298200 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298510 218051
rect 298200 217989 298510 218023
rect 298200 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298510 217989
rect 298200 209175 298510 217961
rect 298200 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298510 209175
rect 298200 209113 298510 209147
rect 298200 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298510 209113
rect 298200 209051 298510 209085
rect 298200 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298510 209051
rect 298200 208989 298510 209023
rect 298200 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298510 208989
rect 298200 200175 298510 208961
rect 298200 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298510 200175
rect 298200 200113 298510 200147
rect 298200 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298510 200113
rect 298200 200051 298510 200085
rect 298200 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298510 200051
rect 298200 199989 298510 200023
rect 298200 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298510 199989
rect 298200 191175 298510 199961
rect 298200 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298510 191175
rect 298200 191113 298510 191147
rect 298200 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298510 191113
rect 298200 191051 298510 191085
rect 298200 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298510 191051
rect 298200 190989 298510 191023
rect 298200 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298510 190989
rect 298200 182175 298510 190961
rect 298200 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298510 182175
rect 298200 182113 298510 182147
rect 298200 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298510 182113
rect 298200 182051 298510 182085
rect 298200 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298510 182051
rect 298200 181989 298510 182023
rect 298200 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298510 181989
rect 298200 173175 298510 181961
rect 298200 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298510 173175
rect 298200 173113 298510 173147
rect 298200 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298510 173113
rect 298200 173051 298510 173085
rect 298200 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298510 173051
rect 298200 172989 298510 173023
rect 298200 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298510 172989
rect 298200 164175 298510 172961
rect 298200 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298510 164175
rect 298200 164113 298510 164147
rect 298200 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298510 164113
rect 298200 164051 298510 164085
rect 298200 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298510 164051
rect 298200 163989 298510 164023
rect 298200 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298510 163989
rect 298200 155175 298510 163961
rect 298200 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298510 155175
rect 298200 155113 298510 155147
rect 298200 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298510 155113
rect 298200 155051 298510 155085
rect 298200 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298510 155051
rect 298200 154989 298510 155023
rect 298200 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298510 154989
rect 298200 146175 298510 154961
rect 298200 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298510 146175
rect 298200 146113 298510 146147
rect 298200 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298510 146113
rect 298200 146051 298510 146085
rect 298200 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298510 146051
rect 298200 145989 298510 146023
rect 298200 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298510 145989
rect 298200 137175 298510 145961
rect 298200 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298510 137175
rect 298200 137113 298510 137147
rect 298200 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298510 137113
rect 298200 137051 298510 137085
rect 298200 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298510 137051
rect 298200 136989 298510 137023
rect 298200 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298510 136989
rect 298200 128175 298510 136961
rect 298200 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298510 128175
rect 298200 128113 298510 128147
rect 298200 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298510 128113
rect 298200 128051 298510 128085
rect 298200 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298510 128051
rect 298200 127989 298510 128023
rect 298200 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298510 127989
rect 298200 119175 298510 127961
rect 298200 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298510 119175
rect 298200 119113 298510 119147
rect 298200 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298510 119113
rect 298200 119051 298510 119085
rect 298200 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298510 119051
rect 298200 118989 298510 119023
rect 298200 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298510 118989
rect 298200 110175 298510 118961
rect 298200 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298510 110175
rect 298200 110113 298510 110147
rect 298200 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298510 110113
rect 298200 110051 298510 110085
rect 298200 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298510 110051
rect 298200 109989 298510 110023
rect 298200 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298510 109989
rect 298200 101175 298510 109961
rect 298200 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298510 101175
rect 298200 101113 298510 101147
rect 298200 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298510 101113
rect 298200 101051 298510 101085
rect 298200 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298510 101051
rect 298200 100989 298510 101023
rect 298200 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298510 100989
rect 298200 92175 298510 100961
rect 298200 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298510 92175
rect 298200 92113 298510 92147
rect 298200 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298510 92113
rect 298200 92051 298510 92085
rect 298200 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298510 92051
rect 298200 91989 298510 92023
rect 298200 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298510 91989
rect 298200 83175 298510 91961
rect 298200 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298510 83175
rect 298200 83113 298510 83147
rect 298200 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298510 83113
rect 298200 83051 298510 83085
rect 298200 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298510 83051
rect 298200 82989 298510 83023
rect 298200 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298510 82989
rect 298200 74175 298510 82961
rect 298200 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298510 74175
rect 298200 74113 298510 74147
rect 298200 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298510 74113
rect 298200 74051 298510 74085
rect 298200 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298510 74051
rect 298200 73989 298510 74023
rect 298200 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298510 73989
rect 298200 65175 298510 73961
rect 298200 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298510 65175
rect 298200 65113 298510 65147
rect 298200 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298510 65113
rect 298200 65051 298510 65085
rect 298200 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298510 65051
rect 298200 64989 298510 65023
rect 298200 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298510 64989
rect 298200 56175 298510 64961
rect 298200 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298510 56175
rect 298200 56113 298510 56147
rect 298200 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298510 56113
rect 298200 56051 298510 56085
rect 298200 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298510 56051
rect 298200 55989 298510 56023
rect 298200 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298510 55989
rect 298200 47175 298510 55961
rect 298200 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298510 47175
rect 298200 47113 298510 47147
rect 298200 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298510 47113
rect 298200 47051 298510 47085
rect 298200 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298510 47051
rect 298200 46989 298510 47023
rect 298200 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298510 46989
rect 298200 38175 298510 46961
rect 298200 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298510 38175
rect 298200 38113 298510 38147
rect 298200 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298510 38113
rect 298200 38051 298510 38085
rect 298200 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298510 38051
rect 298200 37989 298510 38023
rect 298200 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298510 37989
rect 298200 29175 298510 37961
rect 298200 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298510 29175
rect 298200 29113 298510 29147
rect 298200 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298510 29113
rect 298200 29051 298510 29085
rect 298200 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298510 29051
rect 298200 28989 298510 29023
rect 298200 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298510 28989
rect 298200 20175 298510 28961
rect 298200 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298510 20175
rect 298200 20113 298510 20147
rect 298200 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298510 20113
rect 298200 20051 298510 20085
rect 298200 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298510 20051
rect 298200 19989 298510 20023
rect 298200 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298510 19989
rect 298200 11175 298510 19961
rect 298200 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298510 11175
rect 298200 11113 298510 11147
rect 298200 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298510 11113
rect 298200 11051 298510 11085
rect 298200 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298510 11051
rect 298200 10989 298510 11023
rect 298200 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298510 10989
rect 298200 2175 298510 10961
rect 298200 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298510 2175
rect 298200 2113 298510 2147
rect 298200 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298510 2113
rect 298200 2051 298510 2085
rect 298200 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298510 2051
rect 298200 1989 298510 2023
rect 298200 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298510 1989
rect 298200 -80 298510 1961
rect 298200 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect 298200 -142 298510 -108
rect 298200 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect 298200 -204 298510 -170
rect 298200 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect 298200 -266 298510 -232
rect 298200 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect 298200 -342 298510 -294
rect 298680 293175 298990 298872
rect 298680 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect 298680 293113 298990 293147
rect 298680 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect 298680 293051 298990 293085
rect 298680 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect 298680 292989 298990 293023
rect 298680 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect 298680 284175 298990 292961
rect 298680 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect 298680 284113 298990 284147
rect 298680 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect 298680 284051 298990 284085
rect 298680 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect 298680 283989 298990 284023
rect 298680 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect 298680 275175 298990 283961
rect 298680 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect 298680 275113 298990 275147
rect 298680 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect 298680 275051 298990 275085
rect 298680 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect 298680 274989 298990 275023
rect 298680 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect 298680 266175 298990 274961
rect 298680 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect 298680 266113 298990 266147
rect 298680 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect 298680 266051 298990 266085
rect 298680 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect 298680 265989 298990 266023
rect 298680 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect 298680 257175 298990 265961
rect 298680 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect 298680 257113 298990 257147
rect 298680 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect 298680 257051 298990 257085
rect 298680 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect 298680 256989 298990 257023
rect 298680 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect 298680 248175 298990 256961
rect 298680 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect 298680 248113 298990 248147
rect 298680 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect 298680 248051 298990 248085
rect 298680 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect 298680 247989 298990 248023
rect 298680 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect 298680 239175 298990 247961
rect 298680 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect 298680 239113 298990 239147
rect 298680 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect 298680 239051 298990 239085
rect 298680 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect 298680 238989 298990 239023
rect 298680 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect 298680 230175 298990 238961
rect 298680 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect 298680 230113 298990 230147
rect 298680 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect 298680 230051 298990 230085
rect 298680 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect 298680 229989 298990 230023
rect 298680 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect 298680 221175 298990 229961
rect 298680 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect 298680 221113 298990 221147
rect 298680 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect 298680 221051 298990 221085
rect 298680 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect 298680 220989 298990 221023
rect 298680 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect 298680 212175 298990 220961
rect 298680 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect 298680 212113 298990 212147
rect 298680 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect 298680 212051 298990 212085
rect 298680 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect 298680 211989 298990 212023
rect 298680 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect 298680 203175 298990 211961
rect 298680 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect 298680 203113 298990 203147
rect 298680 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect 298680 203051 298990 203085
rect 298680 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect 298680 202989 298990 203023
rect 298680 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect 298680 194175 298990 202961
rect 298680 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect 298680 194113 298990 194147
rect 298680 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect 298680 194051 298990 194085
rect 298680 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect 298680 193989 298990 194023
rect 298680 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect 298680 185175 298990 193961
rect 298680 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect 298680 185113 298990 185147
rect 298680 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect 298680 185051 298990 185085
rect 298680 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect 298680 184989 298990 185023
rect 298680 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect 298680 176175 298990 184961
rect 298680 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect 298680 176113 298990 176147
rect 298680 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect 298680 176051 298990 176085
rect 298680 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect 298680 175989 298990 176023
rect 298680 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect 298680 167175 298990 175961
rect 298680 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect 298680 167113 298990 167147
rect 298680 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect 298680 167051 298990 167085
rect 298680 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect 298680 166989 298990 167023
rect 298680 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect 298680 158175 298990 166961
rect 298680 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect 298680 158113 298990 158147
rect 298680 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect 298680 158051 298990 158085
rect 298680 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect 298680 157989 298990 158023
rect 298680 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect 298680 149175 298990 157961
rect 298680 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect 298680 149113 298990 149147
rect 298680 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect 298680 149051 298990 149085
rect 298680 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect 298680 148989 298990 149023
rect 298680 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect 298680 140175 298990 148961
rect 298680 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect 298680 140113 298990 140147
rect 298680 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect 298680 140051 298990 140085
rect 298680 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect 298680 139989 298990 140023
rect 298680 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect 298680 131175 298990 139961
rect 298680 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect 298680 131113 298990 131147
rect 298680 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect 298680 131051 298990 131085
rect 298680 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect 298680 130989 298990 131023
rect 298680 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect 298680 122175 298990 130961
rect 298680 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect 298680 122113 298990 122147
rect 298680 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect 298680 122051 298990 122085
rect 298680 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect 298680 121989 298990 122023
rect 298680 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect 298680 113175 298990 121961
rect 298680 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect 298680 113113 298990 113147
rect 298680 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect 298680 113051 298990 113085
rect 298680 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect 298680 112989 298990 113023
rect 298680 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect 298680 104175 298990 112961
rect 298680 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect 298680 104113 298990 104147
rect 298680 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect 298680 104051 298990 104085
rect 298680 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect 298680 103989 298990 104023
rect 298680 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect 298680 95175 298990 103961
rect 298680 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect 298680 95113 298990 95147
rect 298680 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect 298680 95051 298990 95085
rect 298680 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect 298680 94989 298990 95023
rect 298680 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect 298680 86175 298990 94961
rect 298680 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect 298680 86113 298990 86147
rect 298680 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect 298680 86051 298990 86085
rect 298680 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect 298680 85989 298990 86023
rect 298680 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect 298680 77175 298990 85961
rect 298680 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect 298680 77113 298990 77147
rect 298680 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect 298680 77051 298990 77085
rect 298680 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect 298680 76989 298990 77023
rect 298680 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect 298680 68175 298990 76961
rect 298680 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect 298680 68113 298990 68147
rect 298680 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect 298680 68051 298990 68085
rect 298680 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect 298680 67989 298990 68023
rect 298680 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect 298680 59175 298990 67961
rect 298680 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect 298680 59113 298990 59147
rect 298680 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect 298680 59051 298990 59085
rect 298680 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect 298680 58989 298990 59023
rect 298680 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect 298680 50175 298990 58961
rect 298680 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect 298680 50113 298990 50147
rect 298680 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect 298680 50051 298990 50085
rect 298680 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect 298680 49989 298990 50023
rect 298680 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect 298680 41175 298990 49961
rect 298680 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect 298680 41113 298990 41147
rect 298680 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect 298680 41051 298990 41085
rect 298680 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect 298680 40989 298990 41023
rect 298680 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect 298680 32175 298990 40961
rect 298680 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect 298680 32113 298990 32147
rect 298680 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect 298680 32051 298990 32085
rect 298680 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect 298680 31989 298990 32023
rect 298680 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect 298680 23175 298990 31961
rect 298680 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect 298680 23113 298990 23147
rect 298680 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect 298680 23051 298990 23085
rect 298680 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect 298680 22989 298990 23023
rect 298680 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect 298680 14175 298990 22961
rect 298680 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect 298680 14113 298990 14147
rect 298680 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect 298680 14051 298990 14085
rect 298680 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect 298680 13989 298990 14023
rect 298680 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect 298680 5175 298990 13961
rect 298680 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect 298680 5113 298990 5147
rect 298680 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect 298680 5051 298990 5085
rect 298680 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect 298680 4989 298990 5023
rect 298680 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect 291437 -588 291485 -560
rect 291513 -588 291547 -560
rect 291575 -588 291609 -560
rect 291637 -588 291671 -560
rect 291699 -588 291747 -560
rect 291437 -622 291747 -588
rect 291437 -650 291485 -622
rect 291513 -650 291547 -622
rect 291575 -650 291609 -622
rect 291637 -650 291671 -622
rect 291699 -650 291747 -622
rect 291437 -684 291747 -650
rect 291437 -712 291485 -684
rect 291513 -712 291547 -684
rect 291575 -712 291609 -684
rect 291637 -712 291671 -684
rect 291699 -712 291747 -684
rect 291437 -746 291747 -712
rect 291437 -774 291485 -746
rect 291513 -774 291547 -746
rect 291575 -774 291609 -746
rect 291637 -774 291671 -746
rect 291699 -774 291747 -746
rect 291437 -822 291747 -774
rect 298680 -560 298990 4961
rect 298680 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect 298680 -622 298990 -588
rect 298680 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect 298680 -684 298990 -650
rect 298680 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect 298680 -746 298990 -712
rect 298680 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect 298680 -822 298990 -774
<< via4 >>
rect -910 299058 -882 299086
rect -848 299058 -820 299086
rect -786 299058 -758 299086
rect -724 299058 -696 299086
rect -910 298996 -882 299024
rect -848 298996 -820 299024
rect -786 298996 -758 299024
rect -724 298996 -696 299024
rect -910 298934 -882 298962
rect -848 298934 -820 298962
rect -786 298934 -758 298962
rect -724 298934 -696 298962
rect -910 298872 -882 298900
rect -848 298872 -820 298900
rect -786 298872 -758 298900
rect -724 298872 -696 298900
rect -910 293147 -882 293175
rect -848 293147 -820 293175
rect -786 293147 -758 293175
rect -724 293147 -696 293175
rect -910 293085 -882 293113
rect -848 293085 -820 293113
rect -786 293085 -758 293113
rect -724 293085 -696 293113
rect -910 293023 -882 293051
rect -848 293023 -820 293051
rect -786 293023 -758 293051
rect -724 293023 -696 293051
rect -910 292961 -882 292989
rect -848 292961 -820 292989
rect -786 292961 -758 292989
rect -724 292961 -696 292989
rect -910 284147 -882 284175
rect -848 284147 -820 284175
rect -786 284147 -758 284175
rect -724 284147 -696 284175
rect -910 284085 -882 284113
rect -848 284085 -820 284113
rect -786 284085 -758 284113
rect -724 284085 -696 284113
rect -910 284023 -882 284051
rect -848 284023 -820 284051
rect -786 284023 -758 284051
rect -724 284023 -696 284051
rect -910 283961 -882 283989
rect -848 283961 -820 283989
rect -786 283961 -758 283989
rect -724 283961 -696 283989
rect -910 275147 -882 275175
rect -848 275147 -820 275175
rect -786 275147 -758 275175
rect -724 275147 -696 275175
rect -910 275085 -882 275113
rect -848 275085 -820 275113
rect -786 275085 -758 275113
rect -724 275085 -696 275113
rect -910 275023 -882 275051
rect -848 275023 -820 275051
rect -786 275023 -758 275051
rect -724 275023 -696 275051
rect -910 274961 -882 274989
rect -848 274961 -820 274989
rect -786 274961 -758 274989
rect -724 274961 -696 274989
rect -910 266147 -882 266175
rect -848 266147 -820 266175
rect -786 266147 -758 266175
rect -724 266147 -696 266175
rect -910 266085 -882 266113
rect -848 266085 -820 266113
rect -786 266085 -758 266113
rect -724 266085 -696 266113
rect -910 266023 -882 266051
rect -848 266023 -820 266051
rect -786 266023 -758 266051
rect -724 266023 -696 266051
rect -910 265961 -882 265989
rect -848 265961 -820 265989
rect -786 265961 -758 265989
rect -724 265961 -696 265989
rect -910 257147 -882 257175
rect -848 257147 -820 257175
rect -786 257147 -758 257175
rect -724 257147 -696 257175
rect -910 257085 -882 257113
rect -848 257085 -820 257113
rect -786 257085 -758 257113
rect -724 257085 -696 257113
rect -910 257023 -882 257051
rect -848 257023 -820 257051
rect -786 257023 -758 257051
rect -724 257023 -696 257051
rect -910 256961 -882 256989
rect -848 256961 -820 256989
rect -786 256961 -758 256989
rect -724 256961 -696 256989
rect -910 248147 -882 248175
rect -848 248147 -820 248175
rect -786 248147 -758 248175
rect -724 248147 -696 248175
rect -910 248085 -882 248113
rect -848 248085 -820 248113
rect -786 248085 -758 248113
rect -724 248085 -696 248113
rect -910 248023 -882 248051
rect -848 248023 -820 248051
rect -786 248023 -758 248051
rect -724 248023 -696 248051
rect -910 247961 -882 247989
rect -848 247961 -820 247989
rect -786 247961 -758 247989
rect -724 247961 -696 247989
rect -910 239147 -882 239175
rect -848 239147 -820 239175
rect -786 239147 -758 239175
rect -724 239147 -696 239175
rect -910 239085 -882 239113
rect -848 239085 -820 239113
rect -786 239085 -758 239113
rect -724 239085 -696 239113
rect -910 239023 -882 239051
rect -848 239023 -820 239051
rect -786 239023 -758 239051
rect -724 239023 -696 239051
rect -910 238961 -882 238989
rect -848 238961 -820 238989
rect -786 238961 -758 238989
rect -724 238961 -696 238989
rect -910 230147 -882 230175
rect -848 230147 -820 230175
rect -786 230147 -758 230175
rect -724 230147 -696 230175
rect -910 230085 -882 230113
rect -848 230085 -820 230113
rect -786 230085 -758 230113
rect -724 230085 -696 230113
rect -910 230023 -882 230051
rect -848 230023 -820 230051
rect -786 230023 -758 230051
rect -724 230023 -696 230051
rect -910 229961 -882 229989
rect -848 229961 -820 229989
rect -786 229961 -758 229989
rect -724 229961 -696 229989
rect -910 221147 -882 221175
rect -848 221147 -820 221175
rect -786 221147 -758 221175
rect -724 221147 -696 221175
rect -910 221085 -882 221113
rect -848 221085 -820 221113
rect -786 221085 -758 221113
rect -724 221085 -696 221113
rect -910 221023 -882 221051
rect -848 221023 -820 221051
rect -786 221023 -758 221051
rect -724 221023 -696 221051
rect -910 220961 -882 220989
rect -848 220961 -820 220989
rect -786 220961 -758 220989
rect -724 220961 -696 220989
rect -910 212147 -882 212175
rect -848 212147 -820 212175
rect -786 212147 -758 212175
rect -724 212147 -696 212175
rect -910 212085 -882 212113
rect -848 212085 -820 212113
rect -786 212085 -758 212113
rect -724 212085 -696 212113
rect -910 212023 -882 212051
rect -848 212023 -820 212051
rect -786 212023 -758 212051
rect -724 212023 -696 212051
rect -910 211961 -882 211989
rect -848 211961 -820 211989
rect -786 211961 -758 211989
rect -724 211961 -696 211989
rect -910 203147 -882 203175
rect -848 203147 -820 203175
rect -786 203147 -758 203175
rect -724 203147 -696 203175
rect -910 203085 -882 203113
rect -848 203085 -820 203113
rect -786 203085 -758 203113
rect -724 203085 -696 203113
rect -910 203023 -882 203051
rect -848 203023 -820 203051
rect -786 203023 -758 203051
rect -724 203023 -696 203051
rect -910 202961 -882 202989
rect -848 202961 -820 202989
rect -786 202961 -758 202989
rect -724 202961 -696 202989
rect -910 194147 -882 194175
rect -848 194147 -820 194175
rect -786 194147 -758 194175
rect -724 194147 -696 194175
rect -910 194085 -882 194113
rect -848 194085 -820 194113
rect -786 194085 -758 194113
rect -724 194085 -696 194113
rect -910 194023 -882 194051
rect -848 194023 -820 194051
rect -786 194023 -758 194051
rect -724 194023 -696 194051
rect -910 193961 -882 193989
rect -848 193961 -820 193989
rect -786 193961 -758 193989
rect -724 193961 -696 193989
rect -910 185147 -882 185175
rect -848 185147 -820 185175
rect -786 185147 -758 185175
rect -724 185147 -696 185175
rect -910 185085 -882 185113
rect -848 185085 -820 185113
rect -786 185085 -758 185113
rect -724 185085 -696 185113
rect -910 185023 -882 185051
rect -848 185023 -820 185051
rect -786 185023 -758 185051
rect -724 185023 -696 185051
rect -910 184961 -882 184989
rect -848 184961 -820 184989
rect -786 184961 -758 184989
rect -724 184961 -696 184989
rect -910 176147 -882 176175
rect -848 176147 -820 176175
rect -786 176147 -758 176175
rect -724 176147 -696 176175
rect -910 176085 -882 176113
rect -848 176085 -820 176113
rect -786 176085 -758 176113
rect -724 176085 -696 176113
rect -910 176023 -882 176051
rect -848 176023 -820 176051
rect -786 176023 -758 176051
rect -724 176023 -696 176051
rect -910 175961 -882 175989
rect -848 175961 -820 175989
rect -786 175961 -758 175989
rect -724 175961 -696 175989
rect -910 167147 -882 167175
rect -848 167147 -820 167175
rect -786 167147 -758 167175
rect -724 167147 -696 167175
rect -910 167085 -882 167113
rect -848 167085 -820 167113
rect -786 167085 -758 167113
rect -724 167085 -696 167113
rect -910 167023 -882 167051
rect -848 167023 -820 167051
rect -786 167023 -758 167051
rect -724 167023 -696 167051
rect -910 166961 -882 166989
rect -848 166961 -820 166989
rect -786 166961 -758 166989
rect -724 166961 -696 166989
rect -910 158147 -882 158175
rect -848 158147 -820 158175
rect -786 158147 -758 158175
rect -724 158147 -696 158175
rect -910 158085 -882 158113
rect -848 158085 -820 158113
rect -786 158085 -758 158113
rect -724 158085 -696 158113
rect -910 158023 -882 158051
rect -848 158023 -820 158051
rect -786 158023 -758 158051
rect -724 158023 -696 158051
rect -910 157961 -882 157989
rect -848 157961 -820 157989
rect -786 157961 -758 157989
rect -724 157961 -696 157989
rect -910 149147 -882 149175
rect -848 149147 -820 149175
rect -786 149147 -758 149175
rect -724 149147 -696 149175
rect -910 149085 -882 149113
rect -848 149085 -820 149113
rect -786 149085 -758 149113
rect -724 149085 -696 149113
rect -910 149023 -882 149051
rect -848 149023 -820 149051
rect -786 149023 -758 149051
rect -724 149023 -696 149051
rect -910 148961 -882 148989
rect -848 148961 -820 148989
rect -786 148961 -758 148989
rect -724 148961 -696 148989
rect -910 140147 -882 140175
rect -848 140147 -820 140175
rect -786 140147 -758 140175
rect -724 140147 -696 140175
rect -910 140085 -882 140113
rect -848 140085 -820 140113
rect -786 140085 -758 140113
rect -724 140085 -696 140113
rect -910 140023 -882 140051
rect -848 140023 -820 140051
rect -786 140023 -758 140051
rect -724 140023 -696 140051
rect -910 139961 -882 139989
rect -848 139961 -820 139989
rect -786 139961 -758 139989
rect -724 139961 -696 139989
rect -910 131147 -882 131175
rect -848 131147 -820 131175
rect -786 131147 -758 131175
rect -724 131147 -696 131175
rect -910 131085 -882 131113
rect -848 131085 -820 131113
rect -786 131085 -758 131113
rect -724 131085 -696 131113
rect -910 131023 -882 131051
rect -848 131023 -820 131051
rect -786 131023 -758 131051
rect -724 131023 -696 131051
rect -910 130961 -882 130989
rect -848 130961 -820 130989
rect -786 130961 -758 130989
rect -724 130961 -696 130989
rect -910 122147 -882 122175
rect -848 122147 -820 122175
rect -786 122147 -758 122175
rect -724 122147 -696 122175
rect -910 122085 -882 122113
rect -848 122085 -820 122113
rect -786 122085 -758 122113
rect -724 122085 -696 122113
rect -910 122023 -882 122051
rect -848 122023 -820 122051
rect -786 122023 -758 122051
rect -724 122023 -696 122051
rect -910 121961 -882 121989
rect -848 121961 -820 121989
rect -786 121961 -758 121989
rect -724 121961 -696 121989
rect -910 113147 -882 113175
rect -848 113147 -820 113175
rect -786 113147 -758 113175
rect -724 113147 -696 113175
rect -910 113085 -882 113113
rect -848 113085 -820 113113
rect -786 113085 -758 113113
rect -724 113085 -696 113113
rect -910 113023 -882 113051
rect -848 113023 -820 113051
rect -786 113023 -758 113051
rect -724 113023 -696 113051
rect -910 112961 -882 112989
rect -848 112961 -820 112989
rect -786 112961 -758 112989
rect -724 112961 -696 112989
rect -910 104147 -882 104175
rect -848 104147 -820 104175
rect -786 104147 -758 104175
rect -724 104147 -696 104175
rect -910 104085 -882 104113
rect -848 104085 -820 104113
rect -786 104085 -758 104113
rect -724 104085 -696 104113
rect -910 104023 -882 104051
rect -848 104023 -820 104051
rect -786 104023 -758 104051
rect -724 104023 -696 104051
rect -910 103961 -882 103989
rect -848 103961 -820 103989
rect -786 103961 -758 103989
rect -724 103961 -696 103989
rect -910 95147 -882 95175
rect -848 95147 -820 95175
rect -786 95147 -758 95175
rect -724 95147 -696 95175
rect -910 95085 -882 95113
rect -848 95085 -820 95113
rect -786 95085 -758 95113
rect -724 95085 -696 95113
rect -910 95023 -882 95051
rect -848 95023 -820 95051
rect -786 95023 -758 95051
rect -724 95023 -696 95051
rect -910 94961 -882 94989
rect -848 94961 -820 94989
rect -786 94961 -758 94989
rect -724 94961 -696 94989
rect -910 86147 -882 86175
rect -848 86147 -820 86175
rect -786 86147 -758 86175
rect -724 86147 -696 86175
rect -910 86085 -882 86113
rect -848 86085 -820 86113
rect -786 86085 -758 86113
rect -724 86085 -696 86113
rect -910 86023 -882 86051
rect -848 86023 -820 86051
rect -786 86023 -758 86051
rect -724 86023 -696 86051
rect -910 85961 -882 85989
rect -848 85961 -820 85989
rect -786 85961 -758 85989
rect -724 85961 -696 85989
rect -910 77147 -882 77175
rect -848 77147 -820 77175
rect -786 77147 -758 77175
rect -724 77147 -696 77175
rect -910 77085 -882 77113
rect -848 77085 -820 77113
rect -786 77085 -758 77113
rect -724 77085 -696 77113
rect -910 77023 -882 77051
rect -848 77023 -820 77051
rect -786 77023 -758 77051
rect -724 77023 -696 77051
rect -910 76961 -882 76989
rect -848 76961 -820 76989
rect -786 76961 -758 76989
rect -724 76961 -696 76989
rect -910 68147 -882 68175
rect -848 68147 -820 68175
rect -786 68147 -758 68175
rect -724 68147 -696 68175
rect -910 68085 -882 68113
rect -848 68085 -820 68113
rect -786 68085 -758 68113
rect -724 68085 -696 68113
rect -910 68023 -882 68051
rect -848 68023 -820 68051
rect -786 68023 -758 68051
rect -724 68023 -696 68051
rect -910 67961 -882 67989
rect -848 67961 -820 67989
rect -786 67961 -758 67989
rect -724 67961 -696 67989
rect -910 59147 -882 59175
rect -848 59147 -820 59175
rect -786 59147 -758 59175
rect -724 59147 -696 59175
rect -910 59085 -882 59113
rect -848 59085 -820 59113
rect -786 59085 -758 59113
rect -724 59085 -696 59113
rect -910 59023 -882 59051
rect -848 59023 -820 59051
rect -786 59023 -758 59051
rect -724 59023 -696 59051
rect -910 58961 -882 58989
rect -848 58961 -820 58989
rect -786 58961 -758 58989
rect -724 58961 -696 58989
rect -910 50147 -882 50175
rect -848 50147 -820 50175
rect -786 50147 -758 50175
rect -724 50147 -696 50175
rect -910 50085 -882 50113
rect -848 50085 -820 50113
rect -786 50085 -758 50113
rect -724 50085 -696 50113
rect -910 50023 -882 50051
rect -848 50023 -820 50051
rect -786 50023 -758 50051
rect -724 50023 -696 50051
rect -910 49961 -882 49989
rect -848 49961 -820 49989
rect -786 49961 -758 49989
rect -724 49961 -696 49989
rect -910 41147 -882 41175
rect -848 41147 -820 41175
rect -786 41147 -758 41175
rect -724 41147 -696 41175
rect -910 41085 -882 41113
rect -848 41085 -820 41113
rect -786 41085 -758 41113
rect -724 41085 -696 41113
rect -910 41023 -882 41051
rect -848 41023 -820 41051
rect -786 41023 -758 41051
rect -724 41023 -696 41051
rect -910 40961 -882 40989
rect -848 40961 -820 40989
rect -786 40961 -758 40989
rect -724 40961 -696 40989
rect -910 32147 -882 32175
rect -848 32147 -820 32175
rect -786 32147 -758 32175
rect -724 32147 -696 32175
rect -910 32085 -882 32113
rect -848 32085 -820 32113
rect -786 32085 -758 32113
rect -724 32085 -696 32113
rect -910 32023 -882 32051
rect -848 32023 -820 32051
rect -786 32023 -758 32051
rect -724 32023 -696 32051
rect -910 31961 -882 31989
rect -848 31961 -820 31989
rect -786 31961 -758 31989
rect -724 31961 -696 31989
rect -910 23147 -882 23175
rect -848 23147 -820 23175
rect -786 23147 -758 23175
rect -724 23147 -696 23175
rect -910 23085 -882 23113
rect -848 23085 -820 23113
rect -786 23085 -758 23113
rect -724 23085 -696 23113
rect -910 23023 -882 23051
rect -848 23023 -820 23051
rect -786 23023 -758 23051
rect -724 23023 -696 23051
rect -910 22961 -882 22989
rect -848 22961 -820 22989
rect -786 22961 -758 22989
rect -724 22961 -696 22989
rect -910 14147 -882 14175
rect -848 14147 -820 14175
rect -786 14147 -758 14175
rect -724 14147 -696 14175
rect -910 14085 -882 14113
rect -848 14085 -820 14113
rect -786 14085 -758 14113
rect -724 14085 -696 14113
rect -910 14023 -882 14051
rect -848 14023 -820 14051
rect -786 14023 -758 14051
rect -724 14023 -696 14051
rect -910 13961 -882 13989
rect -848 13961 -820 13989
rect -786 13961 -758 13989
rect -724 13961 -696 13989
rect -910 5147 -882 5175
rect -848 5147 -820 5175
rect -786 5147 -758 5175
rect -724 5147 -696 5175
rect -910 5085 -882 5113
rect -848 5085 -820 5113
rect -786 5085 -758 5113
rect -724 5085 -696 5113
rect -910 5023 -882 5051
rect -848 5023 -820 5051
rect -786 5023 -758 5051
rect -724 5023 -696 5051
rect -910 4961 -882 4989
rect -848 4961 -820 4989
rect -786 4961 -758 4989
rect -724 4961 -696 4989
rect -430 298578 -402 298606
rect -368 298578 -340 298606
rect -306 298578 -278 298606
rect -244 298578 -216 298606
rect -430 298516 -402 298544
rect -368 298516 -340 298544
rect -306 298516 -278 298544
rect -244 298516 -216 298544
rect -430 298454 -402 298482
rect -368 298454 -340 298482
rect -306 298454 -278 298482
rect -244 298454 -216 298482
rect -430 298392 -402 298420
rect -368 298392 -340 298420
rect -306 298392 -278 298420
rect -244 298392 -216 298420
rect -430 290147 -402 290175
rect -368 290147 -340 290175
rect -306 290147 -278 290175
rect -244 290147 -216 290175
rect -430 290085 -402 290113
rect -368 290085 -340 290113
rect -306 290085 -278 290113
rect -244 290085 -216 290113
rect -430 290023 -402 290051
rect -368 290023 -340 290051
rect -306 290023 -278 290051
rect -244 290023 -216 290051
rect -430 289961 -402 289989
rect -368 289961 -340 289989
rect -306 289961 -278 289989
rect -244 289961 -216 289989
rect -430 281147 -402 281175
rect -368 281147 -340 281175
rect -306 281147 -278 281175
rect -244 281147 -216 281175
rect -430 281085 -402 281113
rect -368 281085 -340 281113
rect -306 281085 -278 281113
rect -244 281085 -216 281113
rect -430 281023 -402 281051
rect -368 281023 -340 281051
rect -306 281023 -278 281051
rect -244 281023 -216 281051
rect -430 280961 -402 280989
rect -368 280961 -340 280989
rect -306 280961 -278 280989
rect -244 280961 -216 280989
rect -430 272147 -402 272175
rect -368 272147 -340 272175
rect -306 272147 -278 272175
rect -244 272147 -216 272175
rect -430 272085 -402 272113
rect -368 272085 -340 272113
rect -306 272085 -278 272113
rect -244 272085 -216 272113
rect -430 272023 -402 272051
rect -368 272023 -340 272051
rect -306 272023 -278 272051
rect -244 272023 -216 272051
rect -430 271961 -402 271989
rect -368 271961 -340 271989
rect -306 271961 -278 271989
rect -244 271961 -216 271989
rect -430 263147 -402 263175
rect -368 263147 -340 263175
rect -306 263147 -278 263175
rect -244 263147 -216 263175
rect -430 263085 -402 263113
rect -368 263085 -340 263113
rect -306 263085 -278 263113
rect -244 263085 -216 263113
rect -430 263023 -402 263051
rect -368 263023 -340 263051
rect -306 263023 -278 263051
rect -244 263023 -216 263051
rect -430 262961 -402 262989
rect -368 262961 -340 262989
rect -306 262961 -278 262989
rect -244 262961 -216 262989
rect -430 254147 -402 254175
rect -368 254147 -340 254175
rect -306 254147 -278 254175
rect -244 254147 -216 254175
rect -430 254085 -402 254113
rect -368 254085 -340 254113
rect -306 254085 -278 254113
rect -244 254085 -216 254113
rect -430 254023 -402 254051
rect -368 254023 -340 254051
rect -306 254023 -278 254051
rect -244 254023 -216 254051
rect -430 253961 -402 253989
rect -368 253961 -340 253989
rect -306 253961 -278 253989
rect -244 253961 -216 253989
rect -430 245147 -402 245175
rect -368 245147 -340 245175
rect -306 245147 -278 245175
rect -244 245147 -216 245175
rect -430 245085 -402 245113
rect -368 245085 -340 245113
rect -306 245085 -278 245113
rect -244 245085 -216 245113
rect -430 245023 -402 245051
rect -368 245023 -340 245051
rect -306 245023 -278 245051
rect -244 245023 -216 245051
rect -430 244961 -402 244989
rect -368 244961 -340 244989
rect -306 244961 -278 244989
rect -244 244961 -216 244989
rect -430 236147 -402 236175
rect -368 236147 -340 236175
rect -306 236147 -278 236175
rect -244 236147 -216 236175
rect -430 236085 -402 236113
rect -368 236085 -340 236113
rect -306 236085 -278 236113
rect -244 236085 -216 236113
rect -430 236023 -402 236051
rect -368 236023 -340 236051
rect -306 236023 -278 236051
rect -244 236023 -216 236051
rect -430 235961 -402 235989
rect -368 235961 -340 235989
rect -306 235961 -278 235989
rect -244 235961 -216 235989
rect -430 227147 -402 227175
rect -368 227147 -340 227175
rect -306 227147 -278 227175
rect -244 227147 -216 227175
rect -430 227085 -402 227113
rect -368 227085 -340 227113
rect -306 227085 -278 227113
rect -244 227085 -216 227113
rect -430 227023 -402 227051
rect -368 227023 -340 227051
rect -306 227023 -278 227051
rect -244 227023 -216 227051
rect -430 226961 -402 226989
rect -368 226961 -340 226989
rect -306 226961 -278 226989
rect -244 226961 -216 226989
rect -430 218147 -402 218175
rect -368 218147 -340 218175
rect -306 218147 -278 218175
rect -244 218147 -216 218175
rect -430 218085 -402 218113
rect -368 218085 -340 218113
rect -306 218085 -278 218113
rect -244 218085 -216 218113
rect -430 218023 -402 218051
rect -368 218023 -340 218051
rect -306 218023 -278 218051
rect -244 218023 -216 218051
rect -430 217961 -402 217989
rect -368 217961 -340 217989
rect -306 217961 -278 217989
rect -244 217961 -216 217989
rect -430 209147 -402 209175
rect -368 209147 -340 209175
rect -306 209147 -278 209175
rect -244 209147 -216 209175
rect -430 209085 -402 209113
rect -368 209085 -340 209113
rect -306 209085 -278 209113
rect -244 209085 -216 209113
rect -430 209023 -402 209051
rect -368 209023 -340 209051
rect -306 209023 -278 209051
rect -244 209023 -216 209051
rect -430 208961 -402 208989
rect -368 208961 -340 208989
rect -306 208961 -278 208989
rect -244 208961 -216 208989
rect -430 200147 -402 200175
rect -368 200147 -340 200175
rect -306 200147 -278 200175
rect -244 200147 -216 200175
rect -430 200085 -402 200113
rect -368 200085 -340 200113
rect -306 200085 -278 200113
rect -244 200085 -216 200113
rect -430 200023 -402 200051
rect -368 200023 -340 200051
rect -306 200023 -278 200051
rect -244 200023 -216 200051
rect -430 199961 -402 199989
rect -368 199961 -340 199989
rect -306 199961 -278 199989
rect -244 199961 -216 199989
rect -430 191147 -402 191175
rect -368 191147 -340 191175
rect -306 191147 -278 191175
rect -244 191147 -216 191175
rect -430 191085 -402 191113
rect -368 191085 -340 191113
rect -306 191085 -278 191113
rect -244 191085 -216 191113
rect -430 191023 -402 191051
rect -368 191023 -340 191051
rect -306 191023 -278 191051
rect -244 191023 -216 191051
rect -430 190961 -402 190989
rect -368 190961 -340 190989
rect -306 190961 -278 190989
rect -244 190961 -216 190989
rect -430 182147 -402 182175
rect -368 182147 -340 182175
rect -306 182147 -278 182175
rect -244 182147 -216 182175
rect -430 182085 -402 182113
rect -368 182085 -340 182113
rect -306 182085 -278 182113
rect -244 182085 -216 182113
rect -430 182023 -402 182051
rect -368 182023 -340 182051
rect -306 182023 -278 182051
rect -244 182023 -216 182051
rect -430 181961 -402 181989
rect -368 181961 -340 181989
rect -306 181961 -278 181989
rect -244 181961 -216 181989
rect -430 173147 -402 173175
rect -368 173147 -340 173175
rect -306 173147 -278 173175
rect -244 173147 -216 173175
rect -430 173085 -402 173113
rect -368 173085 -340 173113
rect -306 173085 -278 173113
rect -244 173085 -216 173113
rect -430 173023 -402 173051
rect -368 173023 -340 173051
rect -306 173023 -278 173051
rect -244 173023 -216 173051
rect -430 172961 -402 172989
rect -368 172961 -340 172989
rect -306 172961 -278 172989
rect -244 172961 -216 172989
rect -430 164147 -402 164175
rect -368 164147 -340 164175
rect -306 164147 -278 164175
rect -244 164147 -216 164175
rect -430 164085 -402 164113
rect -368 164085 -340 164113
rect -306 164085 -278 164113
rect -244 164085 -216 164113
rect -430 164023 -402 164051
rect -368 164023 -340 164051
rect -306 164023 -278 164051
rect -244 164023 -216 164051
rect -430 163961 -402 163989
rect -368 163961 -340 163989
rect -306 163961 -278 163989
rect -244 163961 -216 163989
rect -430 155147 -402 155175
rect -368 155147 -340 155175
rect -306 155147 -278 155175
rect -244 155147 -216 155175
rect -430 155085 -402 155113
rect -368 155085 -340 155113
rect -306 155085 -278 155113
rect -244 155085 -216 155113
rect -430 155023 -402 155051
rect -368 155023 -340 155051
rect -306 155023 -278 155051
rect -244 155023 -216 155051
rect -430 154961 -402 154989
rect -368 154961 -340 154989
rect -306 154961 -278 154989
rect -244 154961 -216 154989
rect -430 146147 -402 146175
rect -368 146147 -340 146175
rect -306 146147 -278 146175
rect -244 146147 -216 146175
rect -430 146085 -402 146113
rect -368 146085 -340 146113
rect -306 146085 -278 146113
rect -244 146085 -216 146113
rect -430 146023 -402 146051
rect -368 146023 -340 146051
rect -306 146023 -278 146051
rect -244 146023 -216 146051
rect -430 145961 -402 145989
rect -368 145961 -340 145989
rect -306 145961 -278 145989
rect -244 145961 -216 145989
rect -430 137147 -402 137175
rect -368 137147 -340 137175
rect -306 137147 -278 137175
rect -244 137147 -216 137175
rect -430 137085 -402 137113
rect -368 137085 -340 137113
rect -306 137085 -278 137113
rect -244 137085 -216 137113
rect -430 137023 -402 137051
rect -368 137023 -340 137051
rect -306 137023 -278 137051
rect -244 137023 -216 137051
rect -430 136961 -402 136989
rect -368 136961 -340 136989
rect -306 136961 -278 136989
rect -244 136961 -216 136989
rect -430 128147 -402 128175
rect -368 128147 -340 128175
rect -306 128147 -278 128175
rect -244 128147 -216 128175
rect -430 128085 -402 128113
rect -368 128085 -340 128113
rect -306 128085 -278 128113
rect -244 128085 -216 128113
rect -430 128023 -402 128051
rect -368 128023 -340 128051
rect -306 128023 -278 128051
rect -244 128023 -216 128051
rect -430 127961 -402 127989
rect -368 127961 -340 127989
rect -306 127961 -278 127989
rect -244 127961 -216 127989
rect -430 119147 -402 119175
rect -368 119147 -340 119175
rect -306 119147 -278 119175
rect -244 119147 -216 119175
rect -430 119085 -402 119113
rect -368 119085 -340 119113
rect -306 119085 -278 119113
rect -244 119085 -216 119113
rect -430 119023 -402 119051
rect -368 119023 -340 119051
rect -306 119023 -278 119051
rect -244 119023 -216 119051
rect -430 118961 -402 118989
rect -368 118961 -340 118989
rect -306 118961 -278 118989
rect -244 118961 -216 118989
rect -430 110147 -402 110175
rect -368 110147 -340 110175
rect -306 110147 -278 110175
rect -244 110147 -216 110175
rect -430 110085 -402 110113
rect -368 110085 -340 110113
rect -306 110085 -278 110113
rect -244 110085 -216 110113
rect -430 110023 -402 110051
rect -368 110023 -340 110051
rect -306 110023 -278 110051
rect -244 110023 -216 110051
rect -430 109961 -402 109989
rect -368 109961 -340 109989
rect -306 109961 -278 109989
rect -244 109961 -216 109989
rect -430 101147 -402 101175
rect -368 101147 -340 101175
rect -306 101147 -278 101175
rect -244 101147 -216 101175
rect -430 101085 -402 101113
rect -368 101085 -340 101113
rect -306 101085 -278 101113
rect -244 101085 -216 101113
rect -430 101023 -402 101051
rect -368 101023 -340 101051
rect -306 101023 -278 101051
rect -244 101023 -216 101051
rect -430 100961 -402 100989
rect -368 100961 -340 100989
rect -306 100961 -278 100989
rect -244 100961 -216 100989
rect -430 92147 -402 92175
rect -368 92147 -340 92175
rect -306 92147 -278 92175
rect -244 92147 -216 92175
rect -430 92085 -402 92113
rect -368 92085 -340 92113
rect -306 92085 -278 92113
rect -244 92085 -216 92113
rect -430 92023 -402 92051
rect -368 92023 -340 92051
rect -306 92023 -278 92051
rect -244 92023 -216 92051
rect -430 91961 -402 91989
rect -368 91961 -340 91989
rect -306 91961 -278 91989
rect -244 91961 -216 91989
rect -430 83147 -402 83175
rect -368 83147 -340 83175
rect -306 83147 -278 83175
rect -244 83147 -216 83175
rect -430 83085 -402 83113
rect -368 83085 -340 83113
rect -306 83085 -278 83113
rect -244 83085 -216 83113
rect -430 83023 -402 83051
rect -368 83023 -340 83051
rect -306 83023 -278 83051
rect -244 83023 -216 83051
rect -430 82961 -402 82989
rect -368 82961 -340 82989
rect -306 82961 -278 82989
rect -244 82961 -216 82989
rect -430 74147 -402 74175
rect -368 74147 -340 74175
rect -306 74147 -278 74175
rect -244 74147 -216 74175
rect -430 74085 -402 74113
rect -368 74085 -340 74113
rect -306 74085 -278 74113
rect -244 74085 -216 74113
rect -430 74023 -402 74051
rect -368 74023 -340 74051
rect -306 74023 -278 74051
rect -244 74023 -216 74051
rect -430 73961 -402 73989
rect -368 73961 -340 73989
rect -306 73961 -278 73989
rect -244 73961 -216 73989
rect -430 65147 -402 65175
rect -368 65147 -340 65175
rect -306 65147 -278 65175
rect -244 65147 -216 65175
rect -430 65085 -402 65113
rect -368 65085 -340 65113
rect -306 65085 -278 65113
rect -244 65085 -216 65113
rect -430 65023 -402 65051
rect -368 65023 -340 65051
rect -306 65023 -278 65051
rect -244 65023 -216 65051
rect -430 64961 -402 64989
rect -368 64961 -340 64989
rect -306 64961 -278 64989
rect -244 64961 -216 64989
rect -430 56147 -402 56175
rect -368 56147 -340 56175
rect -306 56147 -278 56175
rect -244 56147 -216 56175
rect -430 56085 -402 56113
rect -368 56085 -340 56113
rect -306 56085 -278 56113
rect -244 56085 -216 56113
rect -430 56023 -402 56051
rect -368 56023 -340 56051
rect -306 56023 -278 56051
rect -244 56023 -216 56051
rect -430 55961 -402 55989
rect -368 55961 -340 55989
rect -306 55961 -278 55989
rect -244 55961 -216 55989
rect -430 47147 -402 47175
rect -368 47147 -340 47175
rect -306 47147 -278 47175
rect -244 47147 -216 47175
rect -430 47085 -402 47113
rect -368 47085 -340 47113
rect -306 47085 -278 47113
rect -244 47085 -216 47113
rect -430 47023 -402 47051
rect -368 47023 -340 47051
rect -306 47023 -278 47051
rect -244 47023 -216 47051
rect -430 46961 -402 46989
rect -368 46961 -340 46989
rect -306 46961 -278 46989
rect -244 46961 -216 46989
rect -430 38147 -402 38175
rect -368 38147 -340 38175
rect -306 38147 -278 38175
rect -244 38147 -216 38175
rect -430 38085 -402 38113
rect -368 38085 -340 38113
rect -306 38085 -278 38113
rect -244 38085 -216 38113
rect -430 38023 -402 38051
rect -368 38023 -340 38051
rect -306 38023 -278 38051
rect -244 38023 -216 38051
rect -430 37961 -402 37989
rect -368 37961 -340 37989
rect -306 37961 -278 37989
rect -244 37961 -216 37989
rect -430 29147 -402 29175
rect -368 29147 -340 29175
rect -306 29147 -278 29175
rect -244 29147 -216 29175
rect -430 29085 -402 29113
rect -368 29085 -340 29113
rect -306 29085 -278 29113
rect -244 29085 -216 29113
rect -430 29023 -402 29051
rect -368 29023 -340 29051
rect -306 29023 -278 29051
rect -244 29023 -216 29051
rect -430 28961 -402 28989
rect -368 28961 -340 28989
rect -306 28961 -278 28989
rect -244 28961 -216 28989
rect -430 20147 -402 20175
rect -368 20147 -340 20175
rect -306 20147 -278 20175
rect -244 20147 -216 20175
rect -430 20085 -402 20113
rect -368 20085 -340 20113
rect -306 20085 -278 20113
rect -244 20085 -216 20113
rect -430 20023 -402 20051
rect -368 20023 -340 20051
rect -306 20023 -278 20051
rect -244 20023 -216 20051
rect -430 19961 -402 19989
rect -368 19961 -340 19989
rect -306 19961 -278 19989
rect -244 19961 -216 19989
rect -430 11147 -402 11175
rect -368 11147 -340 11175
rect -306 11147 -278 11175
rect -244 11147 -216 11175
rect -430 11085 -402 11113
rect -368 11085 -340 11113
rect -306 11085 -278 11113
rect -244 11085 -216 11113
rect -430 11023 -402 11051
rect -368 11023 -340 11051
rect -306 11023 -278 11051
rect -244 11023 -216 11051
rect -430 10961 -402 10989
rect -368 10961 -340 10989
rect -306 10961 -278 10989
rect -244 10961 -216 10989
rect -430 2147 -402 2175
rect -368 2147 -340 2175
rect -306 2147 -278 2175
rect -244 2147 -216 2175
rect -430 2085 -402 2113
rect -368 2085 -340 2113
rect -306 2085 -278 2113
rect -244 2085 -216 2113
rect -430 2023 -402 2051
rect -368 2023 -340 2051
rect -306 2023 -278 2051
rect -244 2023 -216 2051
rect -430 1961 -402 1989
rect -368 1961 -340 1989
rect -306 1961 -278 1989
rect -244 1961 -216 1989
rect -430 -108 -402 -80
rect -368 -108 -340 -80
rect -306 -108 -278 -80
rect -244 -108 -216 -80
rect -430 -170 -402 -142
rect -368 -170 -340 -142
rect -306 -170 -278 -142
rect -244 -170 -216 -142
rect -430 -232 -402 -204
rect -368 -232 -340 -204
rect -306 -232 -278 -204
rect -244 -232 -216 -204
rect -430 -294 -402 -266
rect -368 -294 -340 -266
rect -306 -294 -278 -266
rect -244 -294 -216 -266
rect 1625 298578 1653 298606
rect 1687 298578 1715 298606
rect 1749 298578 1777 298606
rect 1811 298578 1839 298606
rect 1625 298516 1653 298544
rect 1687 298516 1715 298544
rect 1749 298516 1777 298544
rect 1811 298516 1839 298544
rect 1625 298454 1653 298482
rect 1687 298454 1715 298482
rect 1749 298454 1777 298482
rect 1811 298454 1839 298482
rect 1625 298392 1653 298420
rect 1687 298392 1715 298420
rect 1749 298392 1777 298420
rect 1811 298392 1839 298420
rect 1625 290147 1653 290175
rect 1687 290147 1715 290175
rect 1749 290147 1777 290175
rect 1811 290147 1839 290175
rect 1625 290085 1653 290113
rect 1687 290085 1715 290113
rect 1749 290085 1777 290113
rect 1811 290085 1839 290113
rect 1625 290023 1653 290051
rect 1687 290023 1715 290051
rect 1749 290023 1777 290051
rect 1811 290023 1839 290051
rect 1625 289961 1653 289989
rect 1687 289961 1715 289989
rect 1749 289961 1777 289989
rect 1811 289961 1839 289989
rect 1625 281147 1653 281175
rect 1687 281147 1715 281175
rect 1749 281147 1777 281175
rect 1811 281147 1839 281175
rect 1625 281085 1653 281113
rect 1687 281085 1715 281113
rect 1749 281085 1777 281113
rect 1811 281085 1839 281113
rect 1625 281023 1653 281051
rect 1687 281023 1715 281051
rect 1749 281023 1777 281051
rect 1811 281023 1839 281051
rect 1625 280961 1653 280989
rect 1687 280961 1715 280989
rect 1749 280961 1777 280989
rect 1811 280961 1839 280989
rect 1625 272147 1653 272175
rect 1687 272147 1715 272175
rect 1749 272147 1777 272175
rect 1811 272147 1839 272175
rect 1625 272085 1653 272113
rect 1687 272085 1715 272113
rect 1749 272085 1777 272113
rect 1811 272085 1839 272113
rect 1625 272023 1653 272051
rect 1687 272023 1715 272051
rect 1749 272023 1777 272051
rect 1811 272023 1839 272051
rect 1625 271961 1653 271989
rect 1687 271961 1715 271989
rect 1749 271961 1777 271989
rect 1811 271961 1839 271989
rect 1625 263147 1653 263175
rect 1687 263147 1715 263175
rect 1749 263147 1777 263175
rect 1811 263147 1839 263175
rect 1625 263085 1653 263113
rect 1687 263085 1715 263113
rect 1749 263085 1777 263113
rect 1811 263085 1839 263113
rect 1625 263023 1653 263051
rect 1687 263023 1715 263051
rect 1749 263023 1777 263051
rect 1811 263023 1839 263051
rect 1625 262961 1653 262989
rect 1687 262961 1715 262989
rect 1749 262961 1777 262989
rect 1811 262961 1839 262989
rect 1625 254147 1653 254175
rect 1687 254147 1715 254175
rect 1749 254147 1777 254175
rect 1811 254147 1839 254175
rect 1625 254085 1653 254113
rect 1687 254085 1715 254113
rect 1749 254085 1777 254113
rect 1811 254085 1839 254113
rect 1625 254023 1653 254051
rect 1687 254023 1715 254051
rect 1749 254023 1777 254051
rect 1811 254023 1839 254051
rect 1625 253961 1653 253989
rect 1687 253961 1715 253989
rect 1749 253961 1777 253989
rect 1811 253961 1839 253989
rect 1625 245147 1653 245175
rect 1687 245147 1715 245175
rect 1749 245147 1777 245175
rect 1811 245147 1839 245175
rect 1625 245085 1653 245113
rect 1687 245085 1715 245113
rect 1749 245085 1777 245113
rect 1811 245085 1839 245113
rect 1625 245023 1653 245051
rect 1687 245023 1715 245051
rect 1749 245023 1777 245051
rect 1811 245023 1839 245051
rect 1625 244961 1653 244989
rect 1687 244961 1715 244989
rect 1749 244961 1777 244989
rect 1811 244961 1839 244989
rect 1625 236147 1653 236175
rect 1687 236147 1715 236175
rect 1749 236147 1777 236175
rect 1811 236147 1839 236175
rect 1625 236085 1653 236113
rect 1687 236085 1715 236113
rect 1749 236085 1777 236113
rect 1811 236085 1839 236113
rect 1625 236023 1653 236051
rect 1687 236023 1715 236051
rect 1749 236023 1777 236051
rect 1811 236023 1839 236051
rect 1625 235961 1653 235989
rect 1687 235961 1715 235989
rect 1749 235961 1777 235989
rect 1811 235961 1839 235989
rect 1625 227147 1653 227175
rect 1687 227147 1715 227175
rect 1749 227147 1777 227175
rect 1811 227147 1839 227175
rect 1625 227085 1653 227113
rect 1687 227085 1715 227113
rect 1749 227085 1777 227113
rect 1811 227085 1839 227113
rect 1625 227023 1653 227051
rect 1687 227023 1715 227051
rect 1749 227023 1777 227051
rect 1811 227023 1839 227051
rect 1625 226961 1653 226989
rect 1687 226961 1715 226989
rect 1749 226961 1777 226989
rect 1811 226961 1839 226989
rect 1625 218147 1653 218175
rect 1687 218147 1715 218175
rect 1749 218147 1777 218175
rect 1811 218147 1839 218175
rect 1625 218085 1653 218113
rect 1687 218085 1715 218113
rect 1749 218085 1777 218113
rect 1811 218085 1839 218113
rect 1625 218023 1653 218051
rect 1687 218023 1715 218051
rect 1749 218023 1777 218051
rect 1811 218023 1839 218051
rect 1625 217961 1653 217989
rect 1687 217961 1715 217989
rect 1749 217961 1777 217989
rect 1811 217961 1839 217989
rect 1625 209147 1653 209175
rect 1687 209147 1715 209175
rect 1749 209147 1777 209175
rect 1811 209147 1839 209175
rect 1625 209085 1653 209113
rect 1687 209085 1715 209113
rect 1749 209085 1777 209113
rect 1811 209085 1839 209113
rect 1625 209023 1653 209051
rect 1687 209023 1715 209051
rect 1749 209023 1777 209051
rect 1811 209023 1839 209051
rect 1625 208961 1653 208989
rect 1687 208961 1715 208989
rect 1749 208961 1777 208989
rect 1811 208961 1839 208989
rect 1625 200147 1653 200175
rect 1687 200147 1715 200175
rect 1749 200147 1777 200175
rect 1811 200147 1839 200175
rect 1625 200085 1653 200113
rect 1687 200085 1715 200113
rect 1749 200085 1777 200113
rect 1811 200085 1839 200113
rect 1625 200023 1653 200051
rect 1687 200023 1715 200051
rect 1749 200023 1777 200051
rect 1811 200023 1839 200051
rect 1625 199961 1653 199989
rect 1687 199961 1715 199989
rect 1749 199961 1777 199989
rect 1811 199961 1839 199989
rect 1625 191147 1653 191175
rect 1687 191147 1715 191175
rect 1749 191147 1777 191175
rect 1811 191147 1839 191175
rect 1625 191085 1653 191113
rect 1687 191085 1715 191113
rect 1749 191085 1777 191113
rect 1811 191085 1839 191113
rect 1625 191023 1653 191051
rect 1687 191023 1715 191051
rect 1749 191023 1777 191051
rect 1811 191023 1839 191051
rect 1625 190961 1653 190989
rect 1687 190961 1715 190989
rect 1749 190961 1777 190989
rect 1811 190961 1839 190989
rect 1625 182147 1653 182175
rect 1687 182147 1715 182175
rect 1749 182147 1777 182175
rect 1811 182147 1839 182175
rect 1625 182085 1653 182113
rect 1687 182085 1715 182113
rect 1749 182085 1777 182113
rect 1811 182085 1839 182113
rect 1625 182023 1653 182051
rect 1687 182023 1715 182051
rect 1749 182023 1777 182051
rect 1811 182023 1839 182051
rect 1625 181961 1653 181989
rect 1687 181961 1715 181989
rect 1749 181961 1777 181989
rect 1811 181961 1839 181989
rect 1625 173147 1653 173175
rect 1687 173147 1715 173175
rect 1749 173147 1777 173175
rect 1811 173147 1839 173175
rect 1625 173085 1653 173113
rect 1687 173085 1715 173113
rect 1749 173085 1777 173113
rect 1811 173085 1839 173113
rect 1625 173023 1653 173051
rect 1687 173023 1715 173051
rect 1749 173023 1777 173051
rect 1811 173023 1839 173051
rect 1625 172961 1653 172989
rect 1687 172961 1715 172989
rect 1749 172961 1777 172989
rect 1811 172961 1839 172989
rect 1625 164147 1653 164175
rect 1687 164147 1715 164175
rect 1749 164147 1777 164175
rect 1811 164147 1839 164175
rect 1625 164085 1653 164113
rect 1687 164085 1715 164113
rect 1749 164085 1777 164113
rect 1811 164085 1839 164113
rect 1625 164023 1653 164051
rect 1687 164023 1715 164051
rect 1749 164023 1777 164051
rect 1811 164023 1839 164051
rect 1625 163961 1653 163989
rect 1687 163961 1715 163989
rect 1749 163961 1777 163989
rect 1811 163961 1839 163989
rect 1625 155147 1653 155175
rect 1687 155147 1715 155175
rect 1749 155147 1777 155175
rect 1811 155147 1839 155175
rect 1625 155085 1653 155113
rect 1687 155085 1715 155113
rect 1749 155085 1777 155113
rect 1811 155085 1839 155113
rect 1625 155023 1653 155051
rect 1687 155023 1715 155051
rect 1749 155023 1777 155051
rect 1811 155023 1839 155051
rect 1625 154961 1653 154989
rect 1687 154961 1715 154989
rect 1749 154961 1777 154989
rect 1811 154961 1839 154989
rect 1625 146147 1653 146175
rect 1687 146147 1715 146175
rect 1749 146147 1777 146175
rect 1811 146147 1839 146175
rect 1625 146085 1653 146113
rect 1687 146085 1715 146113
rect 1749 146085 1777 146113
rect 1811 146085 1839 146113
rect 1625 146023 1653 146051
rect 1687 146023 1715 146051
rect 1749 146023 1777 146051
rect 1811 146023 1839 146051
rect 1625 145961 1653 145989
rect 1687 145961 1715 145989
rect 1749 145961 1777 145989
rect 1811 145961 1839 145989
rect 1625 137147 1653 137175
rect 1687 137147 1715 137175
rect 1749 137147 1777 137175
rect 1811 137147 1839 137175
rect 1625 137085 1653 137113
rect 1687 137085 1715 137113
rect 1749 137085 1777 137113
rect 1811 137085 1839 137113
rect 1625 137023 1653 137051
rect 1687 137023 1715 137051
rect 1749 137023 1777 137051
rect 1811 137023 1839 137051
rect 1625 136961 1653 136989
rect 1687 136961 1715 136989
rect 1749 136961 1777 136989
rect 1811 136961 1839 136989
rect 1625 128147 1653 128175
rect 1687 128147 1715 128175
rect 1749 128147 1777 128175
rect 1811 128147 1839 128175
rect 1625 128085 1653 128113
rect 1687 128085 1715 128113
rect 1749 128085 1777 128113
rect 1811 128085 1839 128113
rect 1625 128023 1653 128051
rect 1687 128023 1715 128051
rect 1749 128023 1777 128051
rect 1811 128023 1839 128051
rect 1625 127961 1653 127989
rect 1687 127961 1715 127989
rect 1749 127961 1777 127989
rect 1811 127961 1839 127989
rect 1625 119147 1653 119175
rect 1687 119147 1715 119175
rect 1749 119147 1777 119175
rect 1811 119147 1839 119175
rect 1625 119085 1653 119113
rect 1687 119085 1715 119113
rect 1749 119085 1777 119113
rect 1811 119085 1839 119113
rect 1625 119023 1653 119051
rect 1687 119023 1715 119051
rect 1749 119023 1777 119051
rect 1811 119023 1839 119051
rect 1625 118961 1653 118989
rect 1687 118961 1715 118989
rect 1749 118961 1777 118989
rect 1811 118961 1839 118989
rect 1625 110147 1653 110175
rect 1687 110147 1715 110175
rect 1749 110147 1777 110175
rect 1811 110147 1839 110175
rect 1625 110085 1653 110113
rect 1687 110085 1715 110113
rect 1749 110085 1777 110113
rect 1811 110085 1839 110113
rect 1625 110023 1653 110051
rect 1687 110023 1715 110051
rect 1749 110023 1777 110051
rect 1811 110023 1839 110051
rect 1625 109961 1653 109989
rect 1687 109961 1715 109989
rect 1749 109961 1777 109989
rect 1811 109961 1839 109989
rect 1625 101147 1653 101175
rect 1687 101147 1715 101175
rect 1749 101147 1777 101175
rect 1811 101147 1839 101175
rect 1625 101085 1653 101113
rect 1687 101085 1715 101113
rect 1749 101085 1777 101113
rect 1811 101085 1839 101113
rect 1625 101023 1653 101051
rect 1687 101023 1715 101051
rect 1749 101023 1777 101051
rect 1811 101023 1839 101051
rect 1625 100961 1653 100989
rect 1687 100961 1715 100989
rect 1749 100961 1777 100989
rect 1811 100961 1839 100989
rect 1625 92147 1653 92175
rect 1687 92147 1715 92175
rect 1749 92147 1777 92175
rect 1811 92147 1839 92175
rect 1625 92085 1653 92113
rect 1687 92085 1715 92113
rect 1749 92085 1777 92113
rect 1811 92085 1839 92113
rect 1625 92023 1653 92051
rect 1687 92023 1715 92051
rect 1749 92023 1777 92051
rect 1811 92023 1839 92051
rect 1625 91961 1653 91989
rect 1687 91961 1715 91989
rect 1749 91961 1777 91989
rect 1811 91961 1839 91989
rect 1625 83147 1653 83175
rect 1687 83147 1715 83175
rect 1749 83147 1777 83175
rect 1811 83147 1839 83175
rect 1625 83085 1653 83113
rect 1687 83085 1715 83113
rect 1749 83085 1777 83113
rect 1811 83085 1839 83113
rect 1625 83023 1653 83051
rect 1687 83023 1715 83051
rect 1749 83023 1777 83051
rect 1811 83023 1839 83051
rect 1625 82961 1653 82989
rect 1687 82961 1715 82989
rect 1749 82961 1777 82989
rect 1811 82961 1839 82989
rect 1625 74147 1653 74175
rect 1687 74147 1715 74175
rect 1749 74147 1777 74175
rect 1811 74147 1839 74175
rect 1625 74085 1653 74113
rect 1687 74085 1715 74113
rect 1749 74085 1777 74113
rect 1811 74085 1839 74113
rect 1625 74023 1653 74051
rect 1687 74023 1715 74051
rect 1749 74023 1777 74051
rect 1811 74023 1839 74051
rect 1625 73961 1653 73989
rect 1687 73961 1715 73989
rect 1749 73961 1777 73989
rect 1811 73961 1839 73989
rect 1625 65147 1653 65175
rect 1687 65147 1715 65175
rect 1749 65147 1777 65175
rect 1811 65147 1839 65175
rect 1625 65085 1653 65113
rect 1687 65085 1715 65113
rect 1749 65085 1777 65113
rect 1811 65085 1839 65113
rect 1625 65023 1653 65051
rect 1687 65023 1715 65051
rect 1749 65023 1777 65051
rect 1811 65023 1839 65051
rect 1625 64961 1653 64989
rect 1687 64961 1715 64989
rect 1749 64961 1777 64989
rect 1811 64961 1839 64989
rect 1625 56147 1653 56175
rect 1687 56147 1715 56175
rect 1749 56147 1777 56175
rect 1811 56147 1839 56175
rect 1625 56085 1653 56113
rect 1687 56085 1715 56113
rect 1749 56085 1777 56113
rect 1811 56085 1839 56113
rect 1625 56023 1653 56051
rect 1687 56023 1715 56051
rect 1749 56023 1777 56051
rect 1811 56023 1839 56051
rect 1625 55961 1653 55989
rect 1687 55961 1715 55989
rect 1749 55961 1777 55989
rect 1811 55961 1839 55989
rect 1625 47147 1653 47175
rect 1687 47147 1715 47175
rect 1749 47147 1777 47175
rect 1811 47147 1839 47175
rect 1625 47085 1653 47113
rect 1687 47085 1715 47113
rect 1749 47085 1777 47113
rect 1811 47085 1839 47113
rect 1625 47023 1653 47051
rect 1687 47023 1715 47051
rect 1749 47023 1777 47051
rect 1811 47023 1839 47051
rect 1625 46961 1653 46989
rect 1687 46961 1715 46989
rect 1749 46961 1777 46989
rect 1811 46961 1839 46989
rect 1625 38147 1653 38175
rect 1687 38147 1715 38175
rect 1749 38147 1777 38175
rect 1811 38147 1839 38175
rect 1625 38085 1653 38113
rect 1687 38085 1715 38113
rect 1749 38085 1777 38113
rect 1811 38085 1839 38113
rect 1625 38023 1653 38051
rect 1687 38023 1715 38051
rect 1749 38023 1777 38051
rect 1811 38023 1839 38051
rect 1625 37961 1653 37989
rect 1687 37961 1715 37989
rect 1749 37961 1777 37989
rect 1811 37961 1839 37989
rect 1625 29147 1653 29175
rect 1687 29147 1715 29175
rect 1749 29147 1777 29175
rect 1811 29147 1839 29175
rect 1625 29085 1653 29113
rect 1687 29085 1715 29113
rect 1749 29085 1777 29113
rect 1811 29085 1839 29113
rect 1625 29023 1653 29051
rect 1687 29023 1715 29051
rect 1749 29023 1777 29051
rect 1811 29023 1839 29051
rect 1625 28961 1653 28989
rect 1687 28961 1715 28989
rect 1749 28961 1777 28989
rect 1811 28961 1839 28989
rect 1625 20147 1653 20175
rect 1687 20147 1715 20175
rect 1749 20147 1777 20175
rect 1811 20147 1839 20175
rect 1625 20085 1653 20113
rect 1687 20085 1715 20113
rect 1749 20085 1777 20113
rect 1811 20085 1839 20113
rect 1625 20023 1653 20051
rect 1687 20023 1715 20051
rect 1749 20023 1777 20051
rect 1811 20023 1839 20051
rect 1625 19961 1653 19989
rect 1687 19961 1715 19989
rect 1749 19961 1777 19989
rect 1811 19961 1839 19989
rect 1625 11147 1653 11175
rect 1687 11147 1715 11175
rect 1749 11147 1777 11175
rect 1811 11147 1839 11175
rect 1625 11085 1653 11113
rect 1687 11085 1715 11113
rect 1749 11085 1777 11113
rect 1811 11085 1839 11113
rect 1625 11023 1653 11051
rect 1687 11023 1715 11051
rect 1749 11023 1777 11051
rect 1811 11023 1839 11051
rect 1625 10961 1653 10989
rect 1687 10961 1715 10989
rect 1749 10961 1777 10989
rect 1811 10961 1839 10989
rect 1625 2147 1653 2175
rect 1687 2147 1715 2175
rect 1749 2147 1777 2175
rect 1811 2147 1839 2175
rect 1625 2085 1653 2113
rect 1687 2085 1715 2113
rect 1749 2085 1777 2113
rect 1811 2085 1839 2113
rect 1625 2023 1653 2051
rect 1687 2023 1715 2051
rect 1749 2023 1777 2051
rect 1811 2023 1839 2051
rect 1625 1961 1653 1989
rect 1687 1961 1715 1989
rect 1749 1961 1777 1989
rect 1811 1961 1839 1989
rect 1625 -108 1653 -80
rect 1687 -108 1715 -80
rect 1749 -108 1777 -80
rect 1811 -108 1839 -80
rect 1625 -170 1653 -142
rect 1687 -170 1715 -142
rect 1749 -170 1777 -142
rect 1811 -170 1839 -142
rect 1625 -232 1653 -204
rect 1687 -232 1715 -204
rect 1749 -232 1777 -204
rect 1811 -232 1839 -204
rect 1625 -294 1653 -266
rect 1687 -294 1715 -266
rect 1749 -294 1777 -266
rect 1811 -294 1839 -266
rect -910 -588 -882 -560
rect -848 -588 -820 -560
rect -786 -588 -758 -560
rect -724 -588 -696 -560
rect -910 -650 -882 -622
rect -848 -650 -820 -622
rect -786 -650 -758 -622
rect -724 -650 -696 -622
rect -910 -712 -882 -684
rect -848 -712 -820 -684
rect -786 -712 -758 -684
rect -724 -712 -696 -684
rect -910 -774 -882 -746
rect -848 -774 -820 -746
rect -786 -774 -758 -746
rect -724 -774 -696 -746
rect 3485 299058 3513 299086
rect 3547 299058 3575 299086
rect 3609 299058 3637 299086
rect 3671 299058 3699 299086
rect 3485 298996 3513 299024
rect 3547 298996 3575 299024
rect 3609 298996 3637 299024
rect 3671 298996 3699 299024
rect 3485 298934 3513 298962
rect 3547 298934 3575 298962
rect 3609 298934 3637 298962
rect 3671 298934 3699 298962
rect 3485 298872 3513 298900
rect 3547 298872 3575 298900
rect 3609 298872 3637 298900
rect 3671 298872 3699 298900
rect 3485 293147 3513 293175
rect 3547 293147 3575 293175
rect 3609 293147 3637 293175
rect 3671 293147 3699 293175
rect 3485 293085 3513 293113
rect 3547 293085 3575 293113
rect 3609 293085 3637 293113
rect 3671 293085 3699 293113
rect 3485 293023 3513 293051
rect 3547 293023 3575 293051
rect 3609 293023 3637 293051
rect 3671 293023 3699 293051
rect 3485 292961 3513 292989
rect 3547 292961 3575 292989
rect 3609 292961 3637 292989
rect 3671 292961 3699 292989
rect 3485 284147 3513 284175
rect 3547 284147 3575 284175
rect 3609 284147 3637 284175
rect 3671 284147 3699 284175
rect 3485 284085 3513 284113
rect 3547 284085 3575 284113
rect 3609 284085 3637 284113
rect 3671 284085 3699 284113
rect 3485 284023 3513 284051
rect 3547 284023 3575 284051
rect 3609 284023 3637 284051
rect 3671 284023 3699 284051
rect 3485 283961 3513 283989
rect 3547 283961 3575 283989
rect 3609 283961 3637 283989
rect 3671 283961 3699 283989
rect 3485 275147 3513 275175
rect 3547 275147 3575 275175
rect 3609 275147 3637 275175
rect 3671 275147 3699 275175
rect 3485 275085 3513 275113
rect 3547 275085 3575 275113
rect 3609 275085 3637 275113
rect 3671 275085 3699 275113
rect 3485 275023 3513 275051
rect 3547 275023 3575 275051
rect 3609 275023 3637 275051
rect 3671 275023 3699 275051
rect 3485 274961 3513 274989
rect 3547 274961 3575 274989
rect 3609 274961 3637 274989
rect 3671 274961 3699 274989
rect 3485 266147 3513 266175
rect 3547 266147 3575 266175
rect 3609 266147 3637 266175
rect 3671 266147 3699 266175
rect 3485 266085 3513 266113
rect 3547 266085 3575 266113
rect 3609 266085 3637 266113
rect 3671 266085 3699 266113
rect 3485 266023 3513 266051
rect 3547 266023 3575 266051
rect 3609 266023 3637 266051
rect 3671 266023 3699 266051
rect 3485 265961 3513 265989
rect 3547 265961 3575 265989
rect 3609 265961 3637 265989
rect 3671 265961 3699 265989
rect 3485 257147 3513 257175
rect 3547 257147 3575 257175
rect 3609 257147 3637 257175
rect 3671 257147 3699 257175
rect 3485 257085 3513 257113
rect 3547 257085 3575 257113
rect 3609 257085 3637 257113
rect 3671 257085 3699 257113
rect 3485 257023 3513 257051
rect 3547 257023 3575 257051
rect 3609 257023 3637 257051
rect 3671 257023 3699 257051
rect 3485 256961 3513 256989
rect 3547 256961 3575 256989
rect 3609 256961 3637 256989
rect 3671 256961 3699 256989
rect 3485 248147 3513 248175
rect 3547 248147 3575 248175
rect 3609 248147 3637 248175
rect 3671 248147 3699 248175
rect 3485 248085 3513 248113
rect 3547 248085 3575 248113
rect 3609 248085 3637 248113
rect 3671 248085 3699 248113
rect 3485 248023 3513 248051
rect 3547 248023 3575 248051
rect 3609 248023 3637 248051
rect 3671 248023 3699 248051
rect 3485 247961 3513 247989
rect 3547 247961 3575 247989
rect 3609 247961 3637 247989
rect 3671 247961 3699 247989
rect 3485 239147 3513 239175
rect 3547 239147 3575 239175
rect 3609 239147 3637 239175
rect 3671 239147 3699 239175
rect 3485 239085 3513 239113
rect 3547 239085 3575 239113
rect 3609 239085 3637 239113
rect 3671 239085 3699 239113
rect 3485 239023 3513 239051
rect 3547 239023 3575 239051
rect 3609 239023 3637 239051
rect 3671 239023 3699 239051
rect 3485 238961 3513 238989
rect 3547 238961 3575 238989
rect 3609 238961 3637 238989
rect 3671 238961 3699 238989
rect 3485 230147 3513 230175
rect 3547 230147 3575 230175
rect 3609 230147 3637 230175
rect 3671 230147 3699 230175
rect 3485 230085 3513 230113
rect 3547 230085 3575 230113
rect 3609 230085 3637 230113
rect 3671 230085 3699 230113
rect 3485 230023 3513 230051
rect 3547 230023 3575 230051
rect 3609 230023 3637 230051
rect 3671 230023 3699 230051
rect 3485 229961 3513 229989
rect 3547 229961 3575 229989
rect 3609 229961 3637 229989
rect 3671 229961 3699 229989
rect 3485 221147 3513 221175
rect 3547 221147 3575 221175
rect 3609 221147 3637 221175
rect 3671 221147 3699 221175
rect 3485 221085 3513 221113
rect 3547 221085 3575 221113
rect 3609 221085 3637 221113
rect 3671 221085 3699 221113
rect 3485 221023 3513 221051
rect 3547 221023 3575 221051
rect 3609 221023 3637 221051
rect 3671 221023 3699 221051
rect 3485 220961 3513 220989
rect 3547 220961 3575 220989
rect 3609 220961 3637 220989
rect 3671 220961 3699 220989
rect 3485 212147 3513 212175
rect 3547 212147 3575 212175
rect 3609 212147 3637 212175
rect 3671 212147 3699 212175
rect 3485 212085 3513 212113
rect 3547 212085 3575 212113
rect 3609 212085 3637 212113
rect 3671 212085 3699 212113
rect 3485 212023 3513 212051
rect 3547 212023 3575 212051
rect 3609 212023 3637 212051
rect 3671 212023 3699 212051
rect 3485 211961 3513 211989
rect 3547 211961 3575 211989
rect 3609 211961 3637 211989
rect 3671 211961 3699 211989
rect 3485 203147 3513 203175
rect 3547 203147 3575 203175
rect 3609 203147 3637 203175
rect 3671 203147 3699 203175
rect 3485 203085 3513 203113
rect 3547 203085 3575 203113
rect 3609 203085 3637 203113
rect 3671 203085 3699 203113
rect 3485 203023 3513 203051
rect 3547 203023 3575 203051
rect 3609 203023 3637 203051
rect 3671 203023 3699 203051
rect 3485 202961 3513 202989
rect 3547 202961 3575 202989
rect 3609 202961 3637 202989
rect 3671 202961 3699 202989
rect 3485 194147 3513 194175
rect 3547 194147 3575 194175
rect 3609 194147 3637 194175
rect 3671 194147 3699 194175
rect 3485 194085 3513 194113
rect 3547 194085 3575 194113
rect 3609 194085 3637 194113
rect 3671 194085 3699 194113
rect 3485 194023 3513 194051
rect 3547 194023 3575 194051
rect 3609 194023 3637 194051
rect 3671 194023 3699 194051
rect 3485 193961 3513 193989
rect 3547 193961 3575 193989
rect 3609 193961 3637 193989
rect 3671 193961 3699 193989
rect 3485 185147 3513 185175
rect 3547 185147 3575 185175
rect 3609 185147 3637 185175
rect 3671 185147 3699 185175
rect 3485 185085 3513 185113
rect 3547 185085 3575 185113
rect 3609 185085 3637 185113
rect 3671 185085 3699 185113
rect 3485 185023 3513 185051
rect 3547 185023 3575 185051
rect 3609 185023 3637 185051
rect 3671 185023 3699 185051
rect 3485 184961 3513 184989
rect 3547 184961 3575 184989
rect 3609 184961 3637 184989
rect 3671 184961 3699 184989
rect 3485 176147 3513 176175
rect 3547 176147 3575 176175
rect 3609 176147 3637 176175
rect 3671 176147 3699 176175
rect 3485 176085 3513 176113
rect 3547 176085 3575 176113
rect 3609 176085 3637 176113
rect 3671 176085 3699 176113
rect 3485 176023 3513 176051
rect 3547 176023 3575 176051
rect 3609 176023 3637 176051
rect 3671 176023 3699 176051
rect 3485 175961 3513 175989
rect 3547 175961 3575 175989
rect 3609 175961 3637 175989
rect 3671 175961 3699 175989
rect 3485 167147 3513 167175
rect 3547 167147 3575 167175
rect 3609 167147 3637 167175
rect 3671 167147 3699 167175
rect 3485 167085 3513 167113
rect 3547 167085 3575 167113
rect 3609 167085 3637 167113
rect 3671 167085 3699 167113
rect 3485 167023 3513 167051
rect 3547 167023 3575 167051
rect 3609 167023 3637 167051
rect 3671 167023 3699 167051
rect 3485 166961 3513 166989
rect 3547 166961 3575 166989
rect 3609 166961 3637 166989
rect 3671 166961 3699 166989
rect 3485 158147 3513 158175
rect 3547 158147 3575 158175
rect 3609 158147 3637 158175
rect 3671 158147 3699 158175
rect 3485 158085 3513 158113
rect 3547 158085 3575 158113
rect 3609 158085 3637 158113
rect 3671 158085 3699 158113
rect 3485 158023 3513 158051
rect 3547 158023 3575 158051
rect 3609 158023 3637 158051
rect 3671 158023 3699 158051
rect 3485 157961 3513 157989
rect 3547 157961 3575 157989
rect 3609 157961 3637 157989
rect 3671 157961 3699 157989
rect 3485 149147 3513 149175
rect 3547 149147 3575 149175
rect 3609 149147 3637 149175
rect 3671 149147 3699 149175
rect 3485 149085 3513 149113
rect 3547 149085 3575 149113
rect 3609 149085 3637 149113
rect 3671 149085 3699 149113
rect 3485 149023 3513 149051
rect 3547 149023 3575 149051
rect 3609 149023 3637 149051
rect 3671 149023 3699 149051
rect 3485 148961 3513 148989
rect 3547 148961 3575 148989
rect 3609 148961 3637 148989
rect 3671 148961 3699 148989
rect 3485 140147 3513 140175
rect 3547 140147 3575 140175
rect 3609 140147 3637 140175
rect 3671 140147 3699 140175
rect 3485 140085 3513 140113
rect 3547 140085 3575 140113
rect 3609 140085 3637 140113
rect 3671 140085 3699 140113
rect 3485 140023 3513 140051
rect 3547 140023 3575 140051
rect 3609 140023 3637 140051
rect 3671 140023 3699 140051
rect 3485 139961 3513 139989
rect 3547 139961 3575 139989
rect 3609 139961 3637 139989
rect 3671 139961 3699 139989
rect 3485 131147 3513 131175
rect 3547 131147 3575 131175
rect 3609 131147 3637 131175
rect 3671 131147 3699 131175
rect 3485 131085 3513 131113
rect 3547 131085 3575 131113
rect 3609 131085 3637 131113
rect 3671 131085 3699 131113
rect 3485 131023 3513 131051
rect 3547 131023 3575 131051
rect 3609 131023 3637 131051
rect 3671 131023 3699 131051
rect 3485 130961 3513 130989
rect 3547 130961 3575 130989
rect 3609 130961 3637 130989
rect 3671 130961 3699 130989
rect 3485 122147 3513 122175
rect 3547 122147 3575 122175
rect 3609 122147 3637 122175
rect 3671 122147 3699 122175
rect 3485 122085 3513 122113
rect 3547 122085 3575 122113
rect 3609 122085 3637 122113
rect 3671 122085 3699 122113
rect 3485 122023 3513 122051
rect 3547 122023 3575 122051
rect 3609 122023 3637 122051
rect 3671 122023 3699 122051
rect 3485 121961 3513 121989
rect 3547 121961 3575 121989
rect 3609 121961 3637 121989
rect 3671 121961 3699 121989
rect 3485 113147 3513 113175
rect 3547 113147 3575 113175
rect 3609 113147 3637 113175
rect 3671 113147 3699 113175
rect 3485 113085 3513 113113
rect 3547 113085 3575 113113
rect 3609 113085 3637 113113
rect 3671 113085 3699 113113
rect 3485 113023 3513 113051
rect 3547 113023 3575 113051
rect 3609 113023 3637 113051
rect 3671 113023 3699 113051
rect 3485 112961 3513 112989
rect 3547 112961 3575 112989
rect 3609 112961 3637 112989
rect 3671 112961 3699 112989
rect 3485 104147 3513 104175
rect 3547 104147 3575 104175
rect 3609 104147 3637 104175
rect 3671 104147 3699 104175
rect 3485 104085 3513 104113
rect 3547 104085 3575 104113
rect 3609 104085 3637 104113
rect 3671 104085 3699 104113
rect 3485 104023 3513 104051
rect 3547 104023 3575 104051
rect 3609 104023 3637 104051
rect 3671 104023 3699 104051
rect 3485 103961 3513 103989
rect 3547 103961 3575 103989
rect 3609 103961 3637 103989
rect 3671 103961 3699 103989
rect 3485 95147 3513 95175
rect 3547 95147 3575 95175
rect 3609 95147 3637 95175
rect 3671 95147 3699 95175
rect 3485 95085 3513 95113
rect 3547 95085 3575 95113
rect 3609 95085 3637 95113
rect 3671 95085 3699 95113
rect 3485 95023 3513 95051
rect 3547 95023 3575 95051
rect 3609 95023 3637 95051
rect 3671 95023 3699 95051
rect 3485 94961 3513 94989
rect 3547 94961 3575 94989
rect 3609 94961 3637 94989
rect 3671 94961 3699 94989
rect 3485 86147 3513 86175
rect 3547 86147 3575 86175
rect 3609 86147 3637 86175
rect 3671 86147 3699 86175
rect 3485 86085 3513 86113
rect 3547 86085 3575 86113
rect 3609 86085 3637 86113
rect 3671 86085 3699 86113
rect 3485 86023 3513 86051
rect 3547 86023 3575 86051
rect 3609 86023 3637 86051
rect 3671 86023 3699 86051
rect 3485 85961 3513 85989
rect 3547 85961 3575 85989
rect 3609 85961 3637 85989
rect 3671 85961 3699 85989
rect 3485 77147 3513 77175
rect 3547 77147 3575 77175
rect 3609 77147 3637 77175
rect 3671 77147 3699 77175
rect 3485 77085 3513 77113
rect 3547 77085 3575 77113
rect 3609 77085 3637 77113
rect 3671 77085 3699 77113
rect 3485 77023 3513 77051
rect 3547 77023 3575 77051
rect 3609 77023 3637 77051
rect 3671 77023 3699 77051
rect 3485 76961 3513 76989
rect 3547 76961 3575 76989
rect 3609 76961 3637 76989
rect 3671 76961 3699 76989
rect 3485 68147 3513 68175
rect 3547 68147 3575 68175
rect 3609 68147 3637 68175
rect 3671 68147 3699 68175
rect 3485 68085 3513 68113
rect 3547 68085 3575 68113
rect 3609 68085 3637 68113
rect 3671 68085 3699 68113
rect 3485 68023 3513 68051
rect 3547 68023 3575 68051
rect 3609 68023 3637 68051
rect 3671 68023 3699 68051
rect 3485 67961 3513 67989
rect 3547 67961 3575 67989
rect 3609 67961 3637 67989
rect 3671 67961 3699 67989
rect 3485 59147 3513 59175
rect 3547 59147 3575 59175
rect 3609 59147 3637 59175
rect 3671 59147 3699 59175
rect 3485 59085 3513 59113
rect 3547 59085 3575 59113
rect 3609 59085 3637 59113
rect 3671 59085 3699 59113
rect 3485 59023 3513 59051
rect 3547 59023 3575 59051
rect 3609 59023 3637 59051
rect 3671 59023 3699 59051
rect 3485 58961 3513 58989
rect 3547 58961 3575 58989
rect 3609 58961 3637 58989
rect 3671 58961 3699 58989
rect 3485 50147 3513 50175
rect 3547 50147 3575 50175
rect 3609 50147 3637 50175
rect 3671 50147 3699 50175
rect 3485 50085 3513 50113
rect 3547 50085 3575 50113
rect 3609 50085 3637 50113
rect 3671 50085 3699 50113
rect 3485 50023 3513 50051
rect 3547 50023 3575 50051
rect 3609 50023 3637 50051
rect 3671 50023 3699 50051
rect 3485 49961 3513 49989
rect 3547 49961 3575 49989
rect 3609 49961 3637 49989
rect 3671 49961 3699 49989
rect 3485 41147 3513 41175
rect 3547 41147 3575 41175
rect 3609 41147 3637 41175
rect 3671 41147 3699 41175
rect 3485 41085 3513 41113
rect 3547 41085 3575 41113
rect 3609 41085 3637 41113
rect 3671 41085 3699 41113
rect 3485 41023 3513 41051
rect 3547 41023 3575 41051
rect 3609 41023 3637 41051
rect 3671 41023 3699 41051
rect 3485 40961 3513 40989
rect 3547 40961 3575 40989
rect 3609 40961 3637 40989
rect 3671 40961 3699 40989
rect 3485 32147 3513 32175
rect 3547 32147 3575 32175
rect 3609 32147 3637 32175
rect 3671 32147 3699 32175
rect 3485 32085 3513 32113
rect 3547 32085 3575 32113
rect 3609 32085 3637 32113
rect 3671 32085 3699 32113
rect 3485 32023 3513 32051
rect 3547 32023 3575 32051
rect 3609 32023 3637 32051
rect 3671 32023 3699 32051
rect 3485 31961 3513 31989
rect 3547 31961 3575 31989
rect 3609 31961 3637 31989
rect 3671 31961 3699 31989
rect 3485 23147 3513 23175
rect 3547 23147 3575 23175
rect 3609 23147 3637 23175
rect 3671 23147 3699 23175
rect 3485 23085 3513 23113
rect 3547 23085 3575 23113
rect 3609 23085 3637 23113
rect 3671 23085 3699 23113
rect 3485 23023 3513 23051
rect 3547 23023 3575 23051
rect 3609 23023 3637 23051
rect 3671 23023 3699 23051
rect 3485 22961 3513 22989
rect 3547 22961 3575 22989
rect 3609 22961 3637 22989
rect 3671 22961 3699 22989
rect 3485 14147 3513 14175
rect 3547 14147 3575 14175
rect 3609 14147 3637 14175
rect 3671 14147 3699 14175
rect 3485 14085 3513 14113
rect 3547 14085 3575 14113
rect 3609 14085 3637 14113
rect 3671 14085 3699 14113
rect 3485 14023 3513 14051
rect 3547 14023 3575 14051
rect 3609 14023 3637 14051
rect 3671 14023 3699 14051
rect 3485 13961 3513 13989
rect 3547 13961 3575 13989
rect 3609 13961 3637 13989
rect 3671 13961 3699 13989
rect 3485 5147 3513 5175
rect 3547 5147 3575 5175
rect 3609 5147 3637 5175
rect 3671 5147 3699 5175
rect 3485 5085 3513 5113
rect 3547 5085 3575 5113
rect 3609 5085 3637 5113
rect 3671 5085 3699 5113
rect 3485 5023 3513 5051
rect 3547 5023 3575 5051
rect 3609 5023 3637 5051
rect 3671 5023 3699 5051
rect 3485 4961 3513 4989
rect 3547 4961 3575 4989
rect 3609 4961 3637 4989
rect 3671 4961 3699 4989
rect 3485 -588 3513 -560
rect 3547 -588 3575 -560
rect 3609 -588 3637 -560
rect 3671 -588 3699 -560
rect 3485 -650 3513 -622
rect 3547 -650 3575 -622
rect 3609 -650 3637 -622
rect 3671 -650 3699 -622
rect 3485 -712 3513 -684
rect 3547 -712 3575 -684
rect 3609 -712 3637 -684
rect 3671 -712 3699 -684
rect 3485 -774 3513 -746
rect 3547 -774 3575 -746
rect 3609 -774 3637 -746
rect 3671 -774 3699 -746
rect 10625 298578 10653 298606
rect 10687 298578 10715 298606
rect 10749 298578 10777 298606
rect 10811 298578 10839 298606
rect 10625 298516 10653 298544
rect 10687 298516 10715 298544
rect 10749 298516 10777 298544
rect 10811 298516 10839 298544
rect 10625 298454 10653 298482
rect 10687 298454 10715 298482
rect 10749 298454 10777 298482
rect 10811 298454 10839 298482
rect 10625 298392 10653 298420
rect 10687 298392 10715 298420
rect 10749 298392 10777 298420
rect 10811 298392 10839 298420
rect 10625 290147 10653 290175
rect 10687 290147 10715 290175
rect 10749 290147 10777 290175
rect 10811 290147 10839 290175
rect 10625 290085 10653 290113
rect 10687 290085 10715 290113
rect 10749 290085 10777 290113
rect 10811 290085 10839 290113
rect 10625 290023 10653 290051
rect 10687 290023 10715 290051
rect 10749 290023 10777 290051
rect 10811 290023 10839 290051
rect 10625 289961 10653 289989
rect 10687 289961 10715 289989
rect 10749 289961 10777 289989
rect 10811 289961 10839 289989
rect 10625 281147 10653 281175
rect 10687 281147 10715 281175
rect 10749 281147 10777 281175
rect 10811 281147 10839 281175
rect 10625 281085 10653 281113
rect 10687 281085 10715 281113
rect 10749 281085 10777 281113
rect 10811 281085 10839 281113
rect 10625 281023 10653 281051
rect 10687 281023 10715 281051
rect 10749 281023 10777 281051
rect 10811 281023 10839 281051
rect 10625 280961 10653 280989
rect 10687 280961 10715 280989
rect 10749 280961 10777 280989
rect 10811 280961 10839 280989
rect 10625 272147 10653 272175
rect 10687 272147 10715 272175
rect 10749 272147 10777 272175
rect 10811 272147 10839 272175
rect 10625 272085 10653 272113
rect 10687 272085 10715 272113
rect 10749 272085 10777 272113
rect 10811 272085 10839 272113
rect 10625 272023 10653 272051
rect 10687 272023 10715 272051
rect 10749 272023 10777 272051
rect 10811 272023 10839 272051
rect 10625 271961 10653 271989
rect 10687 271961 10715 271989
rect 10749 271961 10777 271989
rect 10811 271961 10839 271989
rect 10625 263147 10653 263175
rect 10687 263147 10715 263175
rect 10749 263147 10777 263175
rect 10811 263147 10839 263175
rect 10625 263085 10653 263113
rect 10687 263085 10715 263113
rect 10749 263085 10777 263113
rect 10811 263085 10839 263113
rect 10625 263023 10653 263051
rect 10687 263023 10715 263051
rect 10749 263023 10777 263051
rect 10811 263023 10839 263051
rect 10625 262961 10653 262989
rect 10687 262961 10715 262989
rect 10749 262961 10777 262989
rect 10811 262961 10839 262989
rect 10625 254147 10653 254175
rect 10687 254147 10715 254175
rect 10749 254147 10777 254175
rect 10811 254147 10839 254175
rect 10625 254085 10653 254113
rect 10687 254085 10715 254113
rect 10749 254085 10777 254113
rect 10811 254085 10839 254113
rect 10625 254023 10653 254051
rect 10687 254023 10715 254051
rect 10749 254023 10777 254051
rect 10811 254023 10839 254051
rect 10625 253961 10653 253989
rect 10687 253961 10715 253989
rect 10749 253961 10777 253989
rect 10811 253961 10839 253989
rect 10625 245147 10653 245175
rect 10687 245147 10715 245175
rect 10749 245147 10777 245175
rect 10811 245147 10839 245175
rect 10625 245085 10653 245113
rect 10687 245085 10715 245113
rect 10749 245085 10777 245113
rect 10811 245085 10839 245113
rect 10625 245023 10653 245051
rect 10687 245023 10715 245051
rect 10749 245023 10777 245051
rect 10811 245023 10839 245051
rect 10625 244961 10653 244989
rect 10687 244961 10715 244989
rect 10749 244961 10777 244989
rect 10811 244961 10839 244989
rect 10625 236147 10653 236175
rect 10687 236147 10715 236175
rect 10749 236147 10777 236175
rect 10811 236147 10839 236175
rect 10625 236085 10653 236113
rect 10687 236085 10715 236113
rect 10749 236085 10777 236113
rect 10811 236085 10839 236113
rect 10625 236023 10653 236051
rect 10687 236023 10715 236051
rect 10749 236023 10777 236051
rect 10811 236023 10839 236051
rect 10625 235961 10653 235989
rect 10687 235961 10715 235989
rect 10749 235961 10777 235989
rect 10811 235961 10839 235989
rect 10625 227147 10653 227175
rect 10687 227147 10715 227175
rect 10749 227147 10777 227175
rect 10811 227147 10839 227175
rect 10625 227085 10653 227113
rect 10687 227085 10715 227113
rect 10749 227085 10777 227113
rect 10811 227085 10839 227113
rect 10625 227023 10653 227051
rect 10687 227023 10715 227051
rect 10749 227023 10777 227051
rect 10811 227023 10839 227051
rect 10625 226961 10653 226989
rect 10687 226961 10715 226989
rect 10749 226961 10777 226989
rect 10811 226961 10839 226989
rect 10625 218147 10653 218175
rect 10687 218147 10715 218175
rect 10749 218147 10777 218175
rect 10811 218147 10839 218175
rect 10625 218085 10653 218113
rect 10687 218085 10715 218113
rect 10749 218085 10777 218113
rect 10811 218085 10839 218113
rect 10625 218023 10653 218051
rect 10687 218023 10715 218051
rect 10749 218023 10777 218051
rect 10811 218023 10839 218051
rect 10625 217961 10653 217989
rect 10687 217961 10715 217989
rect 10749 217961 10777 217989
rect 10811 217961 10839 217989
rect 10625 209147 10653 209175
rect 10687 209147 10715 209175
rect 10749 209147 10777 209175
rect 10811 209147 10839 209175
rect 10625 209085 10653 209113
rect 10687 209085 10715 209113
rect 10749 209085 10777 209113
rect 10811 209085 10839 209113
rect 10625 209023 10653 209051
rect 10687 209023 10715 209051
rect 10749 209023 10777 209051
rect 10811 209023 10839 209051
rect 10625 208961 10653 208989
rect 10687 208961 10715 208989
rect 10749 208961 10777 208989
rect 10811 208961 10839 208989
rect 10625 200147 10653 200175
rect 10687 200147 10715 200175
rect 10749 200147 10777 200175
rect 10811 200147 10839 200175
rect 10625 200085 10653 200113
rect 10687 200085 10715 200113
rect 10749 200085 10777 200113
rect 10811 200085 10839 200113
rect 10625 200023 10653 200051
rect 10687 200023 10715 200051
rect 10749 200023 10777 200051
rect 10811 200023 10839 200051
rect 10625 199961 10653 199989
rect 10687 199961 10715 199989
rect 10749 199961 10777 199989
rect 10811 199961 10839 199989
rect 10625 191147 10653 191175
rect 10687 191147 10715 191175
rect 10749 191147 10777 191175
rect 10811 191147 10839 191175
rect 10625 191085 10653 191113
rect 10687 191085 10715 191113
rect 10749 191085 10777 191113
rect 10811 191085 10839 191113
rect 10625 191023 10653 191051
rect 10687 191023 10715 191051
rect 10749 191023 10777 191051
rect 10811 191023 10839 191051
rect 10625 190961 10653 190989
rect 10687 190961 10715 190989
rect 10749 190961 10777 190989
rect 10811 190961 10839 190989
rect 10625 182147 10653 182175
rect 10687 182147 10715 182175
rect 10749 182147 10777 182175
rect 10811 182147 10839 182175
rect 10625 182085 10653 182113
rect 10687 182085 10715 182113
rect 10749 182085 10777 182113
rect 10811 182085 10839 182113
rect 10625 182023 10653 182051
rect 10687 182023 10715 182051
rect 10749 182023 10777 182051
rect 10811 182023 10839 182051
rect 10625 181961 10653 181989
rect 10687 181961 10715 181989
rect 10749 181961 10777 181989
rect 10811 181961 10839 181989
rect 10625 173147 10653 173175
rect 10687 173147 10715 173175
rect 10749 173147 10777 173175
rect 10811 173147 10839 173175
rect 10625 173085 10653 173113
rect 10687 173085 10715 173113
rect 10749 173085 10777 173113
rect 10811 173085 10839 173113
rect 10625 173023 10653 173051
rect 10687 173023 10715 173051
rect 10749 173023 10777 173051
rect 10811 173023 10839 173051
rect 10625 172961 10653 172989
rect 10687 172961 10715 172989
rect 10749 172961 10777 172989
rect 10811 172961 10839 172989
rect 10625 164147 10653 164175
rect 10687 164147 10715 164175
rect 10749 164147 10777 164175
rect 10811 164147 10839 164175
rect 10625 164085 10653 164113
rect 10687 164085 10715 164113
rect 10749 164085 10777 164113
rect 10811 164085 10839 164113
rect 10625 164023 10653 164051
rect 10687 164023 10715 164051
rect 10749 164023 10777 164051
rect 10811 164023 10839 164051
rect 10625 163961 10653 163989
rect 10687 163961 10715 163989
rect 10749 163961 10777 163989
rect 10811 163961 10839 163989
rect 10625 155147 10653 155175
rect 10687 155147 10715 155175
rect 10749 155147 10777 155175
rect 10811 155147 10839 155175
rect 10625 155085 10653 155113
rect 10687 155085 10715 155113
rect 10749 155085 10777 155113
rect 10811 155085 10839 155113
rect 10625 155023 10653 155051
rect 10687 155023 10715 155051
rect 10749 155023 10777 155051
rect 10811 155023 10839 155051
rect 10625 154961 10653 154989
rect 10687 154961 10715 154989
rect 10749 154961 10777 154989
rect 10811 154961 10839 154989
rect 10625 146147 10653 146175
rect 10687 146147 10715 146175
rect 10749 146147 10777 146175
rect 10811 146147 10839 146175
rect 10625 146085 10653 146113
rect 10687 146085 10715 146113
rect 10749 146085 10777 146113
rect 10811 146085 10839 146113
rect 10625 146023 10653 146051
rect 10687 146023 10715 146051
rect 10749 146023 10777 146051
rect 10811 146023 10839 146051
rect 10625 145961 10653 145989
rect 10687 145961 10715 145989
rect 10749 145961 10777 145989
rect 10811 145961 10839 145989
rect 10625 137147 10653 137175
rect 10687 137147 10715 137175
rect 10749 137147 10777 137175
rect 10811 137147 10839 137175
rect 10625 137085 10653 137113
rect 10687 137085 10715 137113
rect 10749 137085 10777 137113
rect 10811 137085 10839 137113
rect 10625 137023 10653 137051
rect 10687 137023 10715 137051
rect 10749 137023 10777 137051
rect 10811 137023 10839 137051
rect 10625 136961 10653 136989
rect 10687 136961 10715 136989
rect 10749 136961 10777 136989
rect 10811 136961 10839 136989
rect 10625 128147 10653 128175
rect 10687 128147 10715 128175
rect 10749 128147 10777 128175
rect 10811 128147 10839 128175
rect 10625 128085 10653 128113
rect 10687 128085 10715 128113
rect 10749 128085 10777 128113
rect 10811 128085 10839 128113
rect 10625 128023 10653 128051
rect 10687 128023 10715 128051
rect 10749 128023 10777 128051
rect 10811 128023 10839 128051
rect 10625 127961 10653 127989
rect 10687 127961 10715 127989
rect 10749 127961 10777 127989
rect 10811 127961 10839 127989
rect 10625 119147 10653 119175
rect 10687 119147 10715 119175
rect 10749 119147 10777 119175
rect 10811 119147 10839 119175
rect 10625 119085 10653 119113
rect 10687 119085 10715 119113
rect 10749 119085 10777 119113
rect 10811 119085 10839 119113
rect 10625 119023 10653 119051
rect 10687 119023 10715 119051
rect 10749 119023 10777 119051
rect 10811 119023 10839 119051
rect 10625 118961 10653 118989
rect 10687 118961 10715 118989
rect 10749 118961 10777 118989
rect 10811 118961 10839 118989
rect 10625 110147 10653 110175
rect 10687 110147 10715 110175
rect 10749 110147 10777 110175
rect 10811 110147 10839 110175
rect 10625 110085 10653 110113
rect 10687 110085 10715 110113
rect 10749 110085 10777 110113
rect 10811 110085 10839 110113
rect 10625 110023 10653 110051
rect 10687 110023 10715 110051
rect 10749 110023 10777 110051
rect 10811 110023 10839 110051
rect 10625 109961 10653 109989
rect 10687 109961 10715 109989
rect 10749 109961 10777 109989
rect 10811 109961 10839 109989
rect 10625 101147 10653 101175
rect 10687 101147 10715 101175
rect 10749 101147 10777 101175
rect 10811 101147 10839 101175
rect 10625 101085 10653 101113
rect 10687 101085 10715 101113
rect 10749 101085 10777 101113
rect 10811 101085 10839 101113
rect 10625 101023 10653 101051
rect 10687 101023 10715 101051
rect 10749 101023 10777 101051
rect 10811 101023 10839 101051
rect 10625 100961 10653 100989
rect 10687 100961 10715 100989
rect 10749 100961 10777 100989
rect 10811 100961 10839 100989
rect 10625 92147 10653 92175
rect 10687 92147 10715 92175
rect 10749 92147 10777 92175
rect 10811 92147 10839 92175
rect 10625 92085 10653 92113
rect 10687 92085 10715 92113
rect 10749 92085 10777 92113
rect 10811 92085 10839 92113
rect 10625 92023 10653 92051
rect 10687 92023 10715 92051
rect 10749 92023 10777 92051
rect 10811 92023 10839 92051
rect 10625 91961 10653 91989
rect 10687 91961 10715 91989
rect 10749 91961 10777 91989
rect 10811 91961 10839 91989
rect 10625 83147 10653 83175
rect 10687 83147 10715 83175
rect 10749 83147 10777 83175
rect 10811 83147 10839 83175
rect 10625 83085 10653 83113
rect 10687 83085 10715 83113
rect 10749 83085 10777 83113
rect 10811 83085 10839 83113
rect 10625 83023 10653 83051
rect 10687 83023 10715 83051
rect 10749 83023 10777 83051
rect 10811 83023 10839 83051
rect 10625 82961 10653 82989
rect 10687 82961 10715 82989
rect 10749 82961 10777 82989
rect 10811 82961 10839 82989
rect 10625 74147 10653 74175
rect 10687 74147 10715 74175
rect 10749 74147 10777 74175
rect 10811 74147 10839 74175
rect 10625 74085 10653 74113
rect 10687 74085 10715 74113
rect 10749 74085 10777 74113
rect 10811 74085 10839 74113
rect 10625 74023 10653 74051
rect 10687 74023 10715 74051
rect 10749 74023 10777 74051
rect 10811 74023 10839 74051
rect 10625 73961 10653 73989
rect 10687 73961 10715 73989
rect 10749 73961 10777 73989
rect 10811 73961 10839 73989
rect 10625 65147 10653 65175
rect 10687 65147 10715 65175
rect 10749 65147 10777 65175
rect 10811 65147 10839 65175
rect 10625 65085 10653 65113
rect 10687 65085 10715 65113
rect 10749 65085 10777 65113
rect 10811 65085 10839 65113
rect 10625 65023 10653 65051
rect 10687 65023 10715 65051
rect 10749 65023 10777 65051
rect 10811 65023 10839 65051
rect 10625 64961 10653 64989
rect 10687 64961 10715 64989
rect 10749 64961 10777 64989
rect 10811 64961 10839 64989
rect 10625 56147 10653 56175
rect 10687 56147 10715 56175
rect 10749 56147 10777 56175
rect 10811 56147 10839 56175
rect 10625 56085 10653 56113
rect 10687 56085 10715 56113
rect 10749 56085 10777 56113
rect 10811 56085 10839 56113
rect 10625 56023 10653 56051
rect 10687 56023 10715 56051
rect 10749 56023 10777 56051
rect 10811 56023 10839 56051
rect 10625 55961 10653 55989
rect 10687 55961 10715 55989
rect 10749 55961 10777 55989
rect 10811 55961 10839 55989
rect 10625 47147 10653 47175
rect 10687 47147 10715 47175
rect 10749 47147 10777 47175
rect 10811 47147 10839 47175
rect 10625 47085 10653 47113
rect 10687 47085 10715 47113
rect 10749 47085 10777 47113
rect 10811 47085 10839 47113
rect 10625 47023 10653 47051
rect 10687 47023 10715 47051
rect 10749 47023 10777 47051
rect 10811 47023 10839 47051
rect 10625 46961 10653 46989
rect 10687 46961 10715 46989
rect 10749 46961 10777 46989
rect 10811 46961 10839 46989
rect 10625 38147 10653 38175
rect 10687 38147 10715 38175
rect 10749 38147 10777 38175
rect 10811 38147 10839 38175
rect 10625 38085 10653 38113
rect 10687 38085 10715 38113
rect 10749 38085 10777 38113
rect 10811 38085 10839 38113
rect 10625 38023 10653 38051
rect 10687 38023 10715 38051
rect 10749 38023 10777 38051
rect 10811 38023 10839 38051
rect 10625 37961 10653 37989
rect 10687 37961 10715 37989
rect 10749 37961 10777 37989
rect 10811 37961 10839 37989
rect 10625 29147 10653 29175
rect 10687 29147 10715 29175
rect 10749 29147 10777 29175
rect 10811 29147 10839 29175
rect 10625 29085 10653 29113
rect 10687 29085 10715 29113
rect 10749 29085 10777 29113
rect 10811 29085 10839 29113
rect 10625 29023 10653 29051
rect 10687 29023 10715 29051
rect 10749 29023 10777 29051
rect 10811 29023 10839 29051
rect 10625 28961 10653 28989
rect 10687 28961 10715 28989
rect 10749 28961 10777 28989
rect 10811 28961 10839 28989
rect 10625 20147 10653 20175
rect 10687 20147 10715 20175
rect 10749 20147 10777 20175
rect 10811 20147 10839 20175
rect 10625 20085 10653 20113
rect 10687 20085 10715 20113
rect 10749 20085 10777 20113
rect 10811 20085 10839 20113
rect 10625 20023 10653 20051
rect 10687 20023 10715 20051
rect 10749 20023 10777 20051
rect 10811 20023 10839 20051
rect 10625 19961 10653 19989
rect 10687 19961 10715 19989
rect 10749 19961 10777 19989
rect 10811 19961 10839 19989
rect 10625 11147 10653 11175
rect 10687 11147 10715 11175
rect 10749 11147 10777 11175
rect 10811 11147 10839 11175
rect 10625 11085 10653 11113
rect 10687 11085 10715 11113
rect 10749 11085 10777 11113
rect 10811 11085 10839 11113
rect 10625 11023 10653 11051
rect 10687 11023 10715 11051
rect 10749 11023 10777 11051
rect 10811 11023 10839 11051
rect 10625 10961 10653 10989
rect 10687 10961 10715 10989
rect 10749 10961 10777 10989
rect 10811 10961 10839 10989
rect 10625 2147 10653 2175
rect 10687 2147 10715 2175
rect 10749 2147 10777 2175
rect 10811 2147 10839 2175
rect 10625 2085 10653 2113
rect 10687 2085 10715 2113
rect 10749 2085 10777 2113
rect 10811 2085 10839 2113
rect 10625 2023 10653 2051
rect 10687 2023 10715 2051
rect 10749 2023 10777 2051
rect 10811 2023 10839 2051
rect 10625 1961 10653 1989
rect 10687 1961 10715 1989
rect 10749 1961 10777 1989
rect 10811 1961 10839 1989
rect 10625 -108 10653 -80
rect 10687 -108 10715 -80
rect 10749 -108 10777 -80
rect 10811 -108 10839 -80
rect 10625 -170 10653 -142
rect 10687 -170 10715 -142
rect 10749 -170 10777 -142
rect 10811 -170 10839 -142
rect 10625 -232 10653 -204
rect 10687 -232 10715 -204
rect 10749 -232 10777 -204
rect 10811 -232 10839 -204
rect 10625 -294 10653 -266
rect 10687 -294 10715 -266
rect 10749 -294 10777 -266
rect 10811 -294 10839 -266
rect 12485 299058 12513 299086
rect 12547 299058 12575 299086
rect 12609 299058 12637 299086
rect 12671 299058 12699 299086
rect 12485 298996 12513 299024
rect 12547 298996 12575 299024
rect 12609 298996 12637 299024
rect 12671 298996 12699 299024
rect 12485 298934 12513 298962
rect 12547 298934 12575 298962
rect 12609 298934 12637 298962
rect 12671 298934 12699 298962
rect 12485 298872 12513 298900
rect 12547 298872 12575 298900
rect 12609 298872 12637 298900
rect 12671 298872 12699 298900
rect 12485 293147 12513 293175
rect 12547 293147 12575 293175
rect 12609 293147 12637 293175
rect 12671 293147 12699 293175
rect 12485 293085 12513 293113
rect 12547 293085 12575 293113
rect 12609 293085 12637 293113
rect 12671 293085 12699 293113
rect 12485 293023 12513 293051
rect 12547 293023 12575 293051
rect 12609 293023 12637 293051
rect 12671 293023 12699 293051
rect 12485 292961 12513 292989
rect 12547 292961 12575 292989
rect 12609 292961 12637 292989
rect 12671 292961 12699 292989
rect 12485 284147 12513 284175
rect 12547 284147 12575 284175
rect 12609 284147 12637 284175
rect 12671 284147 12699 284175
rect 12485 284085 12513 284113
rect 12547 284085 12575 284113
rect 12609 284085 12637 284113
rect 12671 284085 12699 284113
rect 12485 284023 12513 284051
rect 12547 284023 12575 284051
rect 12609 284023 12637 284051
rect 12671 284023 12699 284051
rect 12485 283961 12513 283989
rect 12547 283961 12575 283989
rect 12609 283961 12637 283989
rect 12671 283961 12699 283989
rect 12485 275147 12513 275175
rect 12547 275147 12575 275175
rect 12609 275147 12637 275175
rect 12671 275147 12699 275175
rect 12485 275085 12513 275113
rect 12547 275085 12575 275113
rect 12609 275085 12637 275113
rect 12671 275085 12699 275113
rect 12485 275023 12513 275051
rect 12547 275023 12575 275051
rect 12609 275023 12637 275051
rect 12671 275023 12699 275051
rect 12485 274961 12513 274989
rect 12547 274961 12575 274989
rect 12609 274961 12637 274989
rect 12671 274961 12699 274989
rect 12485 266147 12513 266175
rect 12547 266147 12575 266175
rect 12609 266147 12637 266175
rect 12671 266147 12699 266175
rect 12485 266085 12513 266113
rect 12547 266085 12575 266113
rect 12609 266085 12637 266113
rect 12671 266085 12699 266113
rect 12485 266023 12513 266051
rect 12547 266023 12575 266051
rect 12609 266023 12637 266051
rect 12671 266023 12699 266051
rect 12485 265961 12513 265989
rect 12547 265961 12575 265989
rect 12609 265961 12637 265989
rect 12671 265961 12699 265989
rect 12485 257147 12513 257175
rect 12547 257147 12575 257175
rect 12609 257147 12637 257175
rect 12671 257147 12699 257175
rect 12485 257085 12513 257113
rect 12547 257085 12575 257113
rect 12609 257085 12637 257113
rect 12671 257085 12699 257113
rect 12485 257023 12513 257051
rect 12547 257023 12575 257051
rect 12609 257023 12637 257051
rect 12671 257023 12699 257051
rect 12485 256961 12513 256989
rect 12547 256961 12575 256989
rect 12609 256961 12637 256989
rect 12671 256961 12699 256989
rect 12485 248147 12513 248175
rect 12547 248147 12575 248175
rect 12609 248147 12637 248175
rect 12671 248147 12699 248175
rect 12485 248085 12513 248113
rect 12547 248085 12575 248113
rect 12609 248085 12637 248113
rect 12671 248085 12699 248113
rect 12485 248023 12513 248051
rect 12547 248023 12575 248051
rect 12609 248023 12637 248051
rect 12671 248023 12699 248051
rect 12485 247961 12513 247989
rect 12547 247961 12575 247989
rect 12609 247961 12637 247989
rect 12671 247961 12699 247989
rect 12485 239147 12513 239175
rect 12547 239147 12575 239175
rect 12609 239147 12637 239175
rect 12671 239147 12699 239175
rect 12485 239085 12513 239113
rect 12547 239085 12575 239113
rect 12609 239085 12637 239113
rect 12671 239085 12699 239113
rect 12485 239023 12513 239051
rect 12547 239023 12575 239051
rect 12609 239023 12637 239051
rect 12671 239023 12699 239051
rect 12485 238961 12513 238989
rect 12547 238961 12575 238989
rect 12609 238961 12637 238989
rect 12671 238961 12699 238989
rect 12485 230147 12513 230175
rect 12547 230147 12575 230175
rect 12609 230147 12637 230175
rect 12671 230147 12699 230175
rect 12485 230085 12513 230113
rect 12547 230085 12575 230113
rect 12609 230085 12637 230113
rect 12671 230085 12699 230113
rect 12485 230023 12513 230051
rect 12547 230023 12575 230051
rect 12609 230023 12637 230051
rect 12671 230023 12699 230051
rect 12485 229961 12513 229989
rect 12547 229961 12575 229989
rect 12609 229961 12637 229989
rect 12671 229961 12699 229989
rect 12485 221147 12513 221175
rect 12547 221147 12575 221175
rect 12609 221147 12637 221175
rect 12671 221147 12699 221175
rect 12485 221085 12513 221113
rect 12547 221085 12575 221113
rect 12609 221085 12637 221113
rect 12671 221085 12699 221113
rect 12485 221023 12513 221051
rect 12547 221023 12575 221051
rect 12609 221023 12637 221051
rect 12671 221023 12699 221051
rect 12485 220961 12513 220989
rect 12547 220961 12575 220989
rect 12609 220961 12637 220989
rect 12671 220961 12699 220989
rect 12485 212147 12513 212175
rect 12547 212147 12575 212175
rect 12609 212147 12637 212175
rect 12671 212147 12699 212175
rect 12485 212085 12513 212113
rect 12547 212085 12575 212113
rect 12609 212085 12637 212113
rect 12671 212085 12699 212113
rect 12485 212023 12513 212051
rect 12547 212023 12575 212051
rect 12609 212023 12637 212051
rect 12671 212023 12699 212051
rect 12485 211961 12513 211989
rect 12547 211961 12575 211989
rect 12609 211961 12637 211989
rect 12671 211961 12699 211989
rect 12485 203147 12513 203175
rect 12547 203147 12575 203175
rect 12609 203147 12637 203175
rect 12671 203147 12699 203175
rect 12485 203085 12513 203113
rect 12547 203085 12575 203113
rect 12609 203085 12637 203113
rect 12671 203085 12699 203113
rect 12485 203023 12513 203051
rect 12547 203023 12575 203051
rect 12609 203023 12637 203051
rect 12671 203023 12699 203051
rect 12485 202961 12513 202989
rect 12547 202961 12575 202989
rect 12609 202961 12637 202989
rect 12671 202961 12699 202989
rect 12485 194147 12513 194175
rect 12547 194147 12575 194175
rect 12609 194147 12637 194175
rect 12671 194147 12699 194175
rect 12485 194085 12513 194113
rect 12547 194085 12575 194113
rect 12609 194085 12637 194113
rect 12671 194085 12699 194113
rect 12485 194023 12513 194051
rect 12547 194023 12575 194051
rect 12609 194023 12637 194051
rect 12671 194023 12699 194051
rect 12485 193961 12513 193989
rect 12547 193961 12575 193989
rect 12609 193961 12637 193989
rect 12671 193961 12699 193989
rect 12485 185147 12513 185175
rect 12547 185147 12575 185175
rect 12609 185147 12637 185175
rect 12671 185147 12699 185175
rect 12485 185085 12513 185113
rect 12547 185085 12575 185113
rect 12609 185085 12637 185113
rect 12671 185085 12699 185113
rect 12485 185023 12513 185051
rect 12547 185023 12575 185051
rect 12609 185023 12637 185051
rect 12671 185023 12699 185051
rect 12485 184961 12513 184989
rect 12547 184961 12575 184989
rect 12609 184961 12637 184989
rect 12671 184961 12699 184989
rect 12485 176147 12513 176175
rect 12547 176147 12575 176175
rect 12609 176147 12637 176175
rect 12671 176147 12699 176175
rect 12485 176085 12513 176113
rect 12547 176085 12575 176113
rect 12609 176085 12637 176113
rect 12671 176085 12699 176113
rect 12485 176023 12513 176051
rect 12547 176023 12575 176051
rect 12609 176023 12637 176051
rect 12671 176023 12699 176051
rect 12485 175961 12513 175989
rect 12547 175961 12575 175989
rect 12609 175961 12637 175989
rect 12671 175961 12699 175989
rect 12485 167147 12513 167175
rect 12547 167147 12575 167175
rect 12609 167147 12637 167175
rect 12671 167147 12699 167175
rect 12485 167085 12513 167113
rect 12547 167085 12575 167113
rect 12609 167085 12637 167113
rect 12671 167085 12699 167113
rect 12485 167023 12513 167051
rect 12547 167023 12575 167051
rect 12609 167023 12637 167051
rect 12671 167023 12699 167051
rect 12485 166961 12513 166989
rect 12547 166961 12575 166989
rect 12609 166961 12637 166989
rect 12671 166961 12699 166989
rect 12485 158147 12513 158175
rect 12547 158147 12575 158175
rect 12609 158147 12637 158175
rect 12671 158147 12699 158175
rect 12485 158085 12513 158113
rect 12547 158085 12575 158113
rect 12609 158085 12637 158113
rect 12671 158085 12699 158113
rect 12485 158023 12513 158051
rect 12547 158023 12575 158051
rect 12609 158023 12637 158051
rect 12671 158023 12699 158051
rect 12485 157961 12513 157989
rect 12547 157961 12575 157989
rect 12609 157961 12637 157989
rect 12671 157961 12699 157989
rect 12485 149147 12513 149175
rect 12547 149147 12575 149175
rect 12609 149147 12637 149175
rect 12671 149147 12699 149175
rect 12485 149085 12513 149113
rect 12547 149085 12575 149113
rect 12609 149085 12637 149113
rect 12671 149085 12699 149113
rect 12485 149023 12513 149051
rect 12547 149023 12575 149051
rect 12609 149023 12637 149051
rect 12671 149023 12699 149051
rect 12485 148961 12513 148989
rect 12547 148961 12575 148989
rect 12609 148961 12637 148989
rect 12671 148961 12699 148989
rect 12485 140147 12513 140175
rect 12547 140147 12575 140175
rect 12609 140147 12637 140175
rect 12671 140147 12699 140175
rect 12485 140085 12513 140113
rect 12547 140085 12575 140113
rect 12609 140085 12637 140113
rect 12671 140085 12699 140113
rect 12485 140023 12513 140051
rect 12547 140023 12575 140051
rect 12609 140023 12637 140051
rect 12671 140023 12699 140051
rect 12485 139961 12513 139989
rect 12547 139961 12575 139989
rect 12609 139961 12637 139989
rect 12671 139961 12699 139989
rect 12485 131147 12513 131175
rect 12547 131147 12575 131175
rect 12609 131147 12637 131175
rect 12671 131147 12699 131175
rect 12485 131085 12513 131113
rect 12547 131085 12575 131113
rect 12609 131085 12637 131113
rect 12671 131085 12699 131113
rect 12485 131023 12513 131051
rect 12547 131023 12575 131051
rect 12609 131023 12637 131051
rect 12671 131023 12699 131051
rect 12485 130961 12513 130989
rect 12547 130961 12575 130989
rect 12609 130961 12637 130989
rect 12671 130961 12699 130989
rect 12485 122147 12513 122175
rect 12547 122147 12575 122175
rect 12609 122147 12637 122175
rect 12671 122147 12699 122175
rect 12485 122085 12513 122113
rect 12547 122085 12575 122113
rect 12609 122085 12637 122113
rect 12671 122085 12699 122113
rect 12485 122023 12513 122051
rect 12547 122023 12575 122051
rect 12609 122023 12637 122051
rect 12671 122023 12699 122051
rect 12485 121961 12513 121989
rect 12547 121961 12575 121989
rect 12609 121961 12637 121989
rect 12671 121961 12699 121989
rect 12485 113147 12513 113175
rect 12547 113147 12575 113175
rect 12609 113147 12637 113175
rect 12671 113147 12699 113175
rect 12485 113085 12513 113113
rect 12547 113085 12575 113113
rect 12609 113085 12637 113113
rect 12671 113085 12699 113113
rect 12485 113023 12513 113051
rect 12547 113023 12575 113051
rect 12609 113023 12637 113051
rect 12671 113023 12699 113051
rect 12485 112961 12513 112989
rect 12547 112961 12575 112989
rect 12609 112961 12637 112989
rect 12671 112961 12699 112989
rect 12485 104147 12513 104175
rect 12547 104147 12575 104175
rect 12609 104147 12637 104175
rect 12671 104147 12699 104175
rect 12485 104085 12513 104113
rect 12547 104085 12575 104113
rect 12609 104085 12637 104113
rect 12671 104085 12699 104113
rect 12485 104023 12513 104051
rect 12547 104023 12575 104051
rect 12609 104023 12637 104051
rect 12671 104023 12699 104051
rect 12485 103961 12513 103989
rect 12547 103961 12575 103989
rect 12609 103961 12637 103989
rect 12671 103961 12699 103989
rect 12485 95147 12513 95175
rect 12547 95147 12575 95175
rect 12609 95147 12637 95175
rect 12671 95147 12699 95175
rect 12485 95085 12513 95113
rect 12547 95085 12575 95113
rect 12609 95085 12637 95113
rect 12671 95085 12699 95113
rect 12485 95023 12513 95051
rect 12547 95023 12575 95051
rect 12609 95023 12637 95051
rect 12671 95023 12699 95051
rect 12485 94961 12513 94989
rect 12547 94961 12575 94989
rect 12609 94961 12637 94989
rect 12671 94961 12699 94989
rect 12485 86147 12513 86175
rect 12547 86147 12575 86175
rect 12609 86147 12637 86175
rect 12671 86147 12699 86175
rect 12485 86085 12513 86113
rect 12547 86085 12575 86113
rect 12609 86085 12637 86113
rect 12671 86085 12699 86113
rect 12485 86023 12513 86051
rect 12547 86023 12575 86051
rect 12609 86023 12637 86051
rect 12671 86023 12699 86051
rect 12485 85961 12513 85989
rect 12547 85961 12575 85989
rect 12609 85961 12637 85989
rect 12671 85961 12699 85989
rect 12485 77147 12513 77175
rect 12547 77147 12575 77175
rect 12609 77147 12637 77175
rect 12671 77147 12699 77175
rect 12485 77085 12513 77113
rect 12547 77085 12575 77113
rect 12609 77085 12637 77113
rect 12671 77085 12699 77113
rect 12485 77023 12513 77051
rect 12547 77023 12575 77051
rect 12609 77023 12637 77051
rect 12671 77023 12699 77051
rect 12485 76961 12513 76989
rect 12547 76961 12575 76989
rect 12609 76961 12637 76989
rect 12671 76961 12699 76989
rect 12485 68147 12513 68175
rect 12547 68147 12575 68175
rect 12609 68147 12637 68175
rect 12671 68147 12699 68175
rect 12485 68085 12513 68113
rect 12547 68085 12575 68113
rect 12609 68085 12637 68113
rect 12671 68085 12699 68113
rect 12485 68023 12513 68051
rect 12547 68023 12575 68051
rect 12609 68023 12637 68051
rect 12671 68023 12699 68051
rect 12485 67961 12513 67989
rect 12547 67961 12575 67989
rect 12609 67961 12637 67989
rect 12671 67961 12699 67989
rect 12485 59147 12513 59175
rect 12547 59147 12575 59175
rect 12609 59147 12637 59175
rect 12671 59147 12699 59175
rect 12485 59085 12513 59113
rect 12547 59085 12575 59113
rect 12609 59085 12637 59113
rect 12671 59085 12699 59113
rect 12485 59023 12513 59051
rect 12547 59023 12575 59051
rect 12609 59023 12637 59051
rect 12671 59023 12699 59051
rect 12485 58961 12513 58989
rect 12547 58961 12575 58989
rect 12609 58961 12637 58989
rect 12671 58961 12699 58989
rect 12485 50147 12513 50175
rect 12547 50147 12575 50175
rect 12609 50147 12637 50175
rect 12671 50147 12699 50175
rect 12485 50085 12513 50113
rect 12547 50085 12575 50113
rect 12609 50085 12637 50113
rect 12671 50085 12699 50113
rect 12485 50023 12513 50051
rect 12547 50023 12575 50051
rect 12609 50023 12637 50051
rect 12671 50023 12699 50051
rect 12485 49961 12513 49989
rect 12547 49961 12575 49989
rect 12609 49961 12637 49989
rect 12671 49961 12699 49989
rect 12485 41147 12513 41175
rect 12547 41147 12575 41175
rect 12609 41147 12637 41175
rect 12671 41147 12699 41175
rect 12485 41085 12513 41113
rect 12547 41085 12575 41113
rect 12609 41085 12637 41113
rect 12671 41085 12699 41113
rect 12485 41023 12513 41051
rect 12547 41023 12575 41051
rect 12609 41023 12637 41051
rect 12671 41023 12699 41051
rect 12485 40961 12513 40989
rect 12547 40961 12575 40989
rect 12609 40961 12637 40989
rect 12671 40961 12699 40989
rect 12485 32147 12513 32175
rect 12547 32147 12575 32175
rect 12609 32147 12637 32175
rect 12671 32147 12699 32175
rect 12485 32085 12513 32113
rect 12547 32085 12575 32113
rect 12609 32085 12637 32113
rect 12671 32085 12699 32113
rect 12485 32023 12513 32051
rect 12547 32023 12575 32051
rect 12609 32023 12637 32051
rect 12671 32023 12699 32051
rect 12485 31961 12513 31989
rect 12547 31961 12575 31989
rect 12609 31961 12637 31989
rect 12671 31961 12699 31989
rect 12485 23147 12513 23175
rect 12547 23147 12575 23175
rect 12609 23147 12637 23175
rect 12671 23147 12699 23175
rect 12485 23085 12513 23113
rect 12547 23085 12575 23113
rect 12609 23085 12637 23113
rect 12671 23085 12699 23113
rect 12485 23023 12513 23051
rect 12547 23023 12575 23051
rect 12609 23023 12637 23051
rect 12671 23023 12699 23051
rect 12485 22961 12513 22989
rect 12547 22961 12575 22989
rect 12609 22961 12637 22989
rect 12671 22961 12699 22989
rect 12485 14147 12513 14175
rect 12547 14147 12575 14175
rect 12609 14147 12637 14175
rect 12671 14147 12699 14175
rect 12485 14085 12513 14113
rect 12547 14085 12575 14113
rect 12609 14085 12637 14113
rect 12671 14085 12699 14113
rect 12485 14023 12513 14051
rect 12547 14023 12575 14051
rect 12609 14023 12637 14051
rect 12671 14023 12699 14051
rect 12485 13961 12513 13989
rect 12547 13961 12575 13989
rect 12609 13961 12637 13989
rect 12671 13961 12699 13989
rect 12485 5147 12513 5175
rect 12547 5147 12575 5175
rect 12609 5147 12637 5175
rect 12671 5147 12699 5175
rect 12485 5085 12513 5113
rect 12547 5085 12575 5113
rect 12609 5085 12637 5113
rect 12671 5085 12699 5113
rect 12485 5023 12513 5051
rect 12547 5023 12575 5051
rect 12609 5023 12637 5051
rect 12671 5023 12699 5051
rect 12485 4961 12513 4989
rect 12547 4961 12575 4989
rect 12609 4961 12637 4989
rect 12671 4961 12699 4989
rect 12485 -588 12513 -560
rect 12547 -588 12575 -560
rect 12609 -588 12637 -560
rect 12671 -588 12699 -560
rect 12485 -650 12513 -622
rect 12547 -650 12575 -622
rect 12609 -650 12637 -622
rect 12671 -650 12699 -622
rect 12485 -712 12513 -684
rect 12547 -712 12575 -684
rect 12609 -712 12637 -684
rect 12671 -712 12699 -684
rect 12485 -774 12513 -746
rect 12547 -774 12575 -746
rect 12609 -774 12637 -746
rect 12671 -774 12699 -746
rect 19625 298578 19653 298606
rect 19687 298578 19715 298606
rect 19749 298578 19777 298606
rect 19811 298578 19839 298606
rect 19625 298516 19653 298544
rect 19687 298516 19715 298544
rect 19749 298516 19777 298544
rect 19811 298516 19839 298544
rect 19625 298454 19653 298482
rect 19687 298454 19715 298482
rect 19749 298454 19777 298482
rect 19811 298454 19839 298482
rect 19625 298392 19653 298420
rect 19687 298392 19715 298420
rect 19749 298392 19777 298420
rect 19811 298392 19839 298420
rect 19625 290147 19653 290175
rect 19687 290147 19715 290175
rect 19749 290147 19777 290175
rect 19811 290147 19839 290175
rect 19625 290085 19653 290113
rect 19687 290085 19715 290113
rect 19749 290085 19777 290113
rect 19811 290085 19839 290113
rect 19625 290023 19653 290051
rect 19687 290023 19715 290051
rect 19749 290023 19777 290051
rect 19811 290023 19839 290051
rect 19625 289961 19653 289989
rect 19687 289961 19715 289989
rect 19749 289961 19777 289989
rect 19811 289961 19839 289989
rect 19625 281147 19653 281175
rect 19687 281147 19715 281175
rect 19749 281147 19777 281175
rect 19811 281147 19839 281175
rect 19625 281085 19653 281113
rect 19687 281085 19715 281113
rect 19749 281085 19777 281113
rect 19811 281085 19839 281113
rect 19625 281023 19653 281051
rect 19687 281023 19715 281051
rect 19749 281023 19777 281051
rect 19811 281023 19839 281051
rect 19625 280961 19653 280989
rect 19687 280961 19715 280989
rect 19749 280961 19777 280989
rect 19811 280961 19839 280989
rect 19625 272147 19653 272175
rect 19687 272147 19715 272175
rect 19749 272147 19777 272175
rect 19811 272147 19839 272175
rect 19625 272085 19653 272113
rect 19687 272085 19715 272113
rect 19749 272085 19777 272113
rect 19811 272085 19839 272113
rect 19625 272023 19653 272051
rect 19687 272023 19715 272051
rect 19749 272023 19777 272051
rect 19811 272023 19839 272051
rect 19625 271961 19653 271989
rect 19687 271961 19715 271989
rect 19749 271961 19777 271989
rect 19811 271961 19839 271989
rect 19625 263147 19653 263175
rect 19687 263147 19715 263175
rect 19749 263147 19777 263175
rect 19811 263147 19839 263175
rect 19625 263085 19653 263113
rect 19687 263085 19715 263113
rect 19749 263085 19777 263113
rect 19811 263085 19839 263113
rect 19625 263023 19653 263051
rect 19687 263023 19715 263051
rect 19749 263023 19777 263051
rect 19811 263023 19839 263051
rect 19625 262961 19653 262989
rect 19687 262961 19715 262989
rect 19749 262961 19777 262989
rect 19811 262961 19839 262989
rect 19625 254147 19653 254175
rect 19687 254147 19715 254175
rect 19749 254147 19777 254175
rect 19811 254147 19839 254175
rect 19625 254085 19653 254113
rect 19687 254085 19715 254113
rect 19749 254085 19777 254113
rect 19811 254085 19839 254113
rect 19625 254023 19653 254051
rect 19687 254023 19715 254051
rect 19749 254023 19777 254051
rect 19811 254023 19839 254051
rect 19625 253961 19653 253989
rect 19687 253961 19715 253989
rect 19749 253961 19777 253989
rect 19811 253961 19839 253989
rect 19625 245147 19653 245175
rect 19687 245147 19715 245175
rect 19749 245147 19777 245175
rect 19811 245147 19839 245175
rect 19625 245085 19653 245113
rect 19687 245085 19715 245113
rect 19749 245085 19777 245113
rect 19811 245085 19839 245113
rect 19625 245023 19653 245051
rect 19687 245023 19715 245051
rect 19749 245023 19777 245051
rect 19811 245023 19839 245051
rect 19625 244961 19653 244989
rect 19687 244961 19715 244989
rect 19749 244961 19777 244989
rect 19811 244961 19839 244989
rect 19625 236147 19653 236175
rect 19687 236147 19715 236175
rect 19749 236147 19777 236175
rect 19811 236147 19839 236175
rect 19625 236085 19653 236113
rect 19687 236085 19715 236113
rect 19749 236085 19777 236113
rect 19811 236085 19839 236113
rect 19625 236023 19653 236051
rect 19687 236023 19715 236051
rect 19749 236023 19777 236051
rect 19811 236023 19839 236051
rect 19625 235961 19653 235989
rect 19687 235961 19715 235989
rect 19749 235961 19777 235989
rect 19811 235961 19839 235989
rect 19625 227147 19653 227175
rect 19687 227147 19715 227175
rect 19749 227147 19777 227175
rect 19811 227147 19839 227175
rect 19625 227085 19653 227113
rect 19687 227085 19715 227113
rect 19749 227085 19777 227113
rect 19811 227085 19839 227113
rect 19625 227023 19653 227051
rect 19687 227023 19715 227051
rect 19749 227023 19777 227051
rect 19811 227023 19839 227051
rect 19625 226961 19653 226989
rect 19687 226961 19715 226989
rect 19749 226961 19777 226989
rect 19811 226961 19839 226989
rect 19625 218147 19653 218175
rect 19687 218147 19715 218175
rect 19749 218147 19777 218175
rect 19811 218147 19839 218175
rect 19625 218085 19653 218113
rect 19687 218085 19715 218113
rect 19749 218085 19777 218113
rect 19811 218085 19839 218113
rect 19625 218023 19653 218051
rect 19687 218023 19715 218051
rect 19749 218023 19777 218051
rect 19811 218023 19839 218051
rect 19625 217961 19653 217989
rect 19687 217961 19715 217989
rect 19749 217961 19777 217989
rect 19811 217961 19839 217989
rect 19625 209147 19653 209175
rect 19687 209147 19715 209175
rect 19749 209147 19777 209175
rect 19811 209147 19839 209175
rect 19625 209085 19653 209113
rect 19687 209085 19715 209113
rect 19749 209085 19777 209113
rect 19811 209085 19839 209113
rect 19625 209023 19653 209051
rect 19687 209023 19715 209051
rect 19749 209023 19777 209051
rect 19811 209023 19839 209051
rect 19625 208961 19653 208989
rect 19687 208961 19715 208989
rect 19749 208961 19777 208989
rect 19811 208961 19839 208989
rect 19625 200147 19653 200175
rect 19687 200147 19715 200175
rect 19749 200147 19777 200175
rect 19811 200147 19839 200175
rect 19625 200085 19653 200113
rect 19687 200085 19715 200113
rect 19749 200085 19777 200113
rect 19811 200085 19839 200113
rect 19625 200023 19653 200051
rect 19687 200023 19715 200051
rect 19749 200023 19777 200051
rect 19811 200023 19839 200051
rect 19625 199961 19653 199989
rect 19687 199961 19715 199989
rect 19749 199961 19777 199989
rect 19811 199961 19839 199989
rect 19625 191147 19653 191175
rect 19687 191147 19715 191175
rect 19749 191147 19777 191175
rect 19811 191147 19839 191175
rect 19625 191085 19653 191113
rect 19687 191085 19715 191113
rect 19749 191085 19777 191113
rect 19811 191085 19839 191113
rect 19625 191023 19653 191051
rect 19687 191023 19715 191051
rect 19749 191023 19777 191051
rect 19811 191023 19839 191051
rect 19625 190961 19653 190989
rect 19687 190961 19715 190989
rect 19749 190961 19777 190989
rect 19811 190961 19839 190989
rect 19625 182147 19653 182175
rect 19687 182147 19715 182175
rect 19749 182147 19777 182175
rect 19811 182147 19839 182175
rect 19625 182085 19653 182113
rect 19687 182085 19715 182113
rect 19749 182085 19777 182113
rect 19811 182085 19839 182113
rect 19625 182023 19653 182051
rect 19687 182023 19715 182051
rect 19749 182023 19777 182051
rect 19811 182023 19839 182051
rect 19625 181961 19653 181989
rect 19687 181961 19715 181989
rect 19749 181961 19777 181989
rect 19811 181961 19839 181989
rect 19625 173147 19653 173175
rect 19687 173147 19715 173175
rect 19749 173147 19777 173175
rect 19811 173147 19839 173175
rect 19625 173085 19653 173113
rect 19687 173085 19715 173113
rect 19749 173085 19777 173113
rect 19811 173085 19839 173113
rect 19625 173023 19653 173051
rect 19687 173023 19715 173051
rect 19749 173023 19777 173051
rect 19811 173023 19839 173051
rect 19625 172961 19653 172989
rect 19687 172961 19715 172989
rect 19749 172961 19777 172989
rect 19811 172961 19839 172989
rect 19625 164147 19653 164175
rect 19687 164147 19715 164175
rect 19749 164147 19777 164175
rect 19811 164147 19839 164175
rect 19625 164085 19653 164113
rect 19687 164085 19715 164113
rect 19749 164085 19777 164113
rect 19811 164085 19839 164113
rect 19625 164023 19653 164051
rect 19687 164023 19715 164051
rect 19749 164023 19777 164051
rect 19811 164023 19839 164051
rect 19625 163961 19653 163989
rect 19687 163961 19715 163989
rect 19749 163961 19777 163989
rect 19811 163961 19839 163989
rect 19625 155147 19653 155175
rect 19687 155147 19715 155175
rect 19749 155147 19777 155175
rect 19811 155147 19839 155175
rect 19625 155085 19653 155113
rect 19687 155085 19715 155113
rect 19749 155085 19777 155113
rect 19811 155085 19839 155113
rect 19625 155023 19653 155051
rect 19687 155023 19715 155051
rect 19749 155023 19777 155051
rect 19811 155023 19839 155051
rect 19625 154961 19653 154989
rect 19687 154961 19715 154989
rect 19749 154961 19777 154989
rect 19811 154961 19839 154989
rect 19625 146147 19653 146175
rect 19687 146147 19715 146175
rect 19749 146147 19777 146175
rect 19811 146147 19839 146175
rect 19625 146085 19653 146113
rect 19687 146085 19715 146113
rect 19749 146085 19777 146113
rect 19811 146085 19839 146113
rect 19625 146023 19653 146051
rect 19687 146023 19715 146051
rect 19749 146023 19777 146051
rect 19811 146023 19839 146051
rect 19625 145961 19653 145989
rect 19687 145961 19715 145989
rect 19749 145961 19777 145989
rect 19811 145961 19839 145989
rect 19625 137147 19653 137175
rect 19687 137147 19715 137175
rect 19749 137147 19777 137175
rect 19811 137147 19839 137175
rect 19625 137085 19653 137113
rect 19687 137085 19715 137113
rect 19749 137085 19777 137113
rect 19811 137085 19839 137113
rect 19625 137023 19653 137051
rect 19687 137023 19715 137051
rect 19749 137023 19777 137051
rect 19811 137023 19839 137051
rect 19625 136961 19653 136989
rect 19687 136961 19715 136989
rect 19749 136961 19777 136989
rect 19811 136961 19839 136989
rect 19625 128147 19653 128175
rect 19687 128147 19715 128175
rect 19749 128147 19777 128175
rect 19811 128147 19839 128175
rect 19625 128085 19653 128113
rect 19687 128085 19715 128113
rect 19749 128085 19777 128113
rect 19811 128085 19839 128113
rect 19625 128023 19653 128051
rect 19687 128023 19715 128051
rect 19749 128023 19777 128051
rect 19811 128023 19839 128051
rect 19625 127961 19653 127989
rect 19687 127961 19715 127989
rect 19749 127961 19777 127989
rect 19811 127961 19839 127989
rect 19625 119147 19653 119175
rect 19687 119147 19715 119175
rect 19749 119147 19777 119175
rect 19811 119147 19839 119175
rect 19625 119085 19653 119113
rect 19687 119085 19715 119113
rect 19749 119085 19777 119113
rect 19811 119085 19839 119113
rect 19625 119023 19653 119051
rect 19687 119023 19715 119051
rect 19749 119023 19777 119051
rect 19811 119023 19839 119051
rect 19625 118961 19653 118989
rect 19687 118961 19715 118989
rect 19749 118961 19777 118989
rect 19811 118961 19839 118989
rect 19625 110147 19653 110175
rect 19687 110147 19715 110175
rect 19749 110147 19777 110175
rect 19811 110147 19839 110175
rect 19625 110085 19653 110113
rect 19687 110085 19715 110113
rect 19749 110085 19777 110113
rect 19811 110085 19839 110113
rect 19625 110023 19653 110051
rect 19687 110023 19715 110051
rect 19749 110023 19777 110051
rect 19811 110023 19839 110051
rect 19625 109961 19653 109989
rect 19687 109961 19715 109989
rect 19749 109961 19777 109989
rect 19811 109961 19839 109989
rect 19625 101147 19653 101175
rect 19687 101147 19715 101175
rect 19749 101147 19777 101175
rect 19811 101147 19839 101175
rect 19625 101085 19653 101113
rect 19687 101085 19715 101113
rect 19749 101085 19777 101113
rect 19811 101085 19839 101113
rect 19625 101023 19653 101051
rect 19687 101023 19715 101051
rect 19749 101023 19777 101051
rect 19811 101023 19839 101051
rect 19625 100961 19653 100989
rect 19687 100961 19715 100989
rect 19749 100961 19777 100989
rect 19811 100961 19839 100989
rect 19625 92147 19653 92175
rect 19687 92147 19715 92175
rect 19749 92147 19777 92175
rect 19811 92147 19839 92175
rect 19625 92085 19653 92113
rect 19687 92085 19715 92113
rect 19749 92085 19777 92113
rect 19811 92085 19839 92113
rect 19625 92023 19653 92051
rect 19687 92023 19715 92051
rect 19749 92023 19777 92051
rect 19811 92023 19839 92051
rect 19625 91961 19653 91989
rect 19687 91961 19715 91989
rect 19749 91961 19777 91989
rect 19811 91961 19839 91989
rect 19625 83147 19653 83175
rect 19687 83147 19715 83175
rect 19749 83147 19777 83175
rect 19811 83147 19839 83175
rect 19625 83085 19653 83113
rect 19687 83085 19715 83113
rect 19749 83085 19777 83113
rect 19811 83085 19839 83113
rect 19625 83023 19653 83051
rect 19687 83023 19715 83051
rect 19749 83023 19777 83051
rect 19811 83023 19839 83051
rect 19625 82961 19653 82989
rect 19687 82961 19715 82989
rect 19749 82961 19777 82989
rect 19811 82961 19839 82989
rect 19625 74147 19653 74175
rect 19687 74147 19715 74175
rect 19749 74147 19777 74175
rect 19811 74147 19839 74175
rect 19625 74085 19653 74113
rect 19687 74085 19715 74113
rect 19749 74085 19777 74113
rect 19811 74085 19839 74113
rect 19625 74023 19653 74051
rect 19687 74023 19715 74051
rect 19749 74023 19777 74051
rect 19811 74023 19839 74051
rect 19625 73961 19653 73989
rect 19687 73961 19715 73989
rect 19749 73961 19777 73989
rect 19811 73961 19839 73989
rect 19625 65147 19653 65175
rect 19687 65147 19715 65175
rect 19749 65147 19777 65175
rect 19811 65147 19839 65175
rect 19625 65085 19653 65113
rect 19687 65085 19715 65113
rect 19749 65085 19777 65113
rect 19811 65085 19839 65113
rect 19625 65023 19653 65051
rect 19687 65023 19715 65051
rect 19749 65023 19777 65051
rect 19811 65023 19839 65051
rect 19625 64961 19653 64989
rect 19687 64961 19715 64989
rect 19749 64961 19777 64989
rect 19811 64961 19839 64989
rect 19625 56147 19653 56175
rect 19687 56147 19715 56175
rect 19749 56147 19777 56175
rect 19811 56147 19839 56175
rect 19625 56085 19653 56113
rect 19687 56085 19715 56113
rect 19749 56085 19777 56113
rect 19811 56085 19839 56113
rect 19625 56023 19653 56051
rect 19687 56023 19715 56051
rect 19749 56023 19777 56051
rect 19811 56023 19839 56051
rect 19625 55961 19653 55989
rect 19687 55961 19715 55989
rect 19749 55961 19777 55989
rect 19811 55961 19839 55989
rect 19625 47147 19653 47175
rect 19687 47147 19715 47175
rect 19749 47147 19777 47175
rect 19811 47147 19839 47175
rect 19625 47085 19653 47113
rect 19687 47085 19715 47113
rect 19749 47085 19777 47113
rect 19811 47085 19839 47113
rect 19625 47023 19653 47051
rect 19687 47023 19715 47051
rect 19749 47023 19777 47051
rect 19811 47023 19839 47051
rect 19625 46961 19653 46989
rect 19687 46961 19715 46989
rect 19749 46961 19777 46989
rect 19811 46961 19839 46989
rect 19625 38147 19653 38175
rect 19687 38147 19715 38175
rect 19749 38147 19777 38175
rect 19811 38147 19839 38175
rect 19625 38085 19653 38113
rect 19687 38085 19715 38113
rect 19749 38085 19777 38113
rect 19811 38085 19839 38113
rect 19625 38023 19653 38051
rect 19687 38023 19715 38051
rect 19749 38023 19777 38051
rect 19811 38023 19839 38051
rect 19625 37961 19653 37989
rect 19687 37961 19715 37989
rect 19749 37961 19777 37989
rect 19811 37961 19839 37989
rect 19625 29147 19653 29175
rect 19687 29147 19715 29175
rect 19749 29147 19777 29175
rect 19811 29147 19839 29175
rect 19625 29085 19653 29113
rect 19687 29085 19715 29113
rect 19749 29085 19777 29113
rect 19811 29085 19839 29113
rect 19625 29023 19653 29051
rect 19687 29023 19715 29051
rect 19749 29023 19777 29051
rect 19811 29023 19839 29051
rect 19625 28961 19653 28989
rect 19687 28961 19715 28989
rect 19749 28961 19777 28989
rect 19811 28961 19839 28989
rect 19625 20147 19653 20175
rect 19687 20147 19715 20175
rect 19749 20147 19777 20175
rect 19811 20147 19839 20175
rect 19625 20085 19653 20113
rect 19687 20085 19715 20113
rect 19749 20085 19777 20113
rect 19811 20085 19839 20113
rect 19625 20023 19653 20051
rect 19687 20023 19715 20051
rect 19749 20023 19777 20051
rect 19811 20023 19839 20051
rect 19625 19961 19653 19989
rect 19687 19961 19715 19989
rect 19749 19961 19777 19989
rect 19811 19961 19839 19989
rect 19625 11147 19653 11175
rect 19687 11147 19715 11175
rect 19749 11147 19777 11175
rect 19811 11147 19839 11175
rect 19625 11085 19653 11113
rect 19687 11085 19715 11113
rect 19749 11085 19777 11113
rect 19811 11085 19839 11113
rect 19625 11023 19653 11051
rect 19687 11023 19715 11051
rect 19749 11023 19777 11051
rect 19811 11023 19839 11051
rect 19625 10961 19653 10989
rect 19687 10961 19715 10989
rect 19749 10961 19777 10989
rect 19811 10961 19839 10989
rect 19625 2147 19653 2175
rect 19687 2147 19715 2175
rect 19749 2147 19777 2175
rect 19811 2147 19839 2175
rect 19625 2085 19653 2113
rect 19687 2085 19715 2113
rect 19749 2085 19777 2113
rect 19811 2085 19839 2113
rect 19625 2023 19653 2051
rect 19687 2023 19715 2051
rect 19749 2023 19777 2051
rect 19811 2023 19839 2051
rect 19625 1961 19653 1989
rect 19687 1961 19715 1989
rect 19749 1961 19777 1989
rect 19811 1961 19839 1989
rect 19625 -108 19653 -80
rect 19687 -108 19715 -80
rect 19749 -108 19777 -80
rect 19811 -108 19839 -80
rect 19625 -170 19653 -142
rect 19687 -170 19715 -142
rect 19749 -170 19777 -142
rect 19811 -170 19839 -142
rect 19625 -232 19653 -204
rect 19687 -232 19715 -204
rect 19749 -232 19777 -204
rect 19811 -232 19839 -204
rect 19625 -294 19653 -266
rect 19687 -294 19715 -266
rect 19749 -294 19777 -266
rect 19811 -294 19839 -266
rect 21485 299058 21513 299086
rect 21547 299058 21575 299086
rect 21609 299058 21637 299086
rect 21671 299058 21699 299086
rect 21485 298996 21513 299024
rect 21547 298996 21575 299024
rect 21609 298996 21637 299024
rect 21671 298996 21699 299024
rect 21485 298934 21513 298962
rect 21547 298934 21575 298962
rect 21609 298934 21637 298962
rect 21671 298934 21699 298962
rect 21485 298872 21513 298900
rect 21547 298872 21575 298900
rect 21609 298872 21637 298900
rect 21671 298872 21699 298900
rect 21485 293147 21513 293175
rect 21547 293147 21575 293175
rect 21609 293147 21637 293175
rect 21671 293147 21699 293175
rect 21485 293085 21513 293113
rect 21547 293085 21575 293113
rect 21609 293085 21637 293113
rect 21671 293085 21699 293113
rect 21485 293023 21513 293051
rect 21547 293023 21575 293051
rect 21609 293023 21637 293051
rect 21671 293023 21699 293051
rect 21485 292961 21513 292989
rect 21547 292961 21575 292989
rect 21609 292961 21637 292989
rect 21671 292961 21699 292989
rect 21485 284147 21513 284175
rect 21547 284147 21575 284175
rect 21609 284147 21637 284175
rect 21671 284147 21699 284175
rect 21485 284085 21513 284113
rect 21547 284085 21575 284113
rect 21609 284085 21637 284113
rect 21671 284085 21699 284113
rect 21485 284023 21513 284051
rect 21547 284023 21575 284051
rect 21609 284023 21637 284051
rect 21671 284023 21699 284051
rect 21485 283961 21513 283989
rect 21547 283961 21575 283989
rect 21609 283961 21637 283989
rect 21671 283961 21699 283989
rect 21485 275147 21513 275175
rect 21547 275147 21575 275175
rect 21609 275147 21637 275175
rect 21671 275147 21699 275175
rect 21485 275085 21513 275113
rect 21547 275085 21575 275113
rect 21609 275085 21637 275113
rect 21671 275085 21699 275113
rect 21485 275023 21513 275051
rect 21547 275023 21575 275051
rect 21609 275023 21637 275051
rect 21671 275023 21699 275051
rect 21485 274961 21513 274989
rect 21547 274961 21575 274989
rect 21609 274961 21637 274989
rect 21671 274961 21699 274989
rect 21485 266147 21513 266175
rect 21547 266147 21575 266175
rect 21609 266147 21637 266175
rect 21671 266147 21699 266175
rect 21485 266085 21513 266113
rect 21547 266085 21575 266113
rect 21609 266085 21637 266113
rect 21671 266085 21699 266113
rect 21485 266023 21513 266051
rect 21547 266023 21575 266051
rect 21609 266023 21637 266051
rect 21671 266023 21699 266051
rect 21485 265961 21513 265989
rect 21547 265961 21575 265989
rect 21609 265961 21637 265989
rect 21671 265961 21699 265989
rect 21485 257147 21513 257175
rect 21547 257147 21575 257175
rect 21609 257147 21637 257175
rect 21671 257147 21699 257175
rect 21485 257085 21513 257113
rect 21547 257085 21575 257113
rect 21609 257085 21637 257113
rect 21671 257085 21699 257113
rect 21485 257023 21513 257051
rect 21547 257023 21575 257051
rect 21609 257023 21637 257051
rect 21671 257023 21699 257051
rect 21485 256961 21513 256989
rect 21547 256961 21575 256989
rect 21609 256961 21637 256989
rect 21671 256961 21699 256989
rect 21485 248147 21513 248175
rect 21547 248147 21575 248175
rect 21609 248147 21637 248175
rect 21671 248147 21699 248175
rect 21485 248085 21513 248113
rect 21547 248085 21575 248113
rect 21609 248085 21637 248113
rect 21671 248085 21699 248113
rect 21485 248023 21513 248051
rect 21547 248023 21575 248051
rect 21609 248023 21637 248051
rect 21671 248023 21699 248051
rect 21485 247961 21513 247989
rect 21547 247961 21575 247989
rect 21609 247961 21637 247989
rect 21671 247961 21699 247989
rect 21485 239147 21513 239175
rect 21547 239147 21575 239175
rect 21609 239147 21637 239175
rect 21671 239147 21699 239175
rect 21485 239085 21513 239113
rect 21547 239085 21575 239113
rect 21609 239085 21637 239113
rect 21671 239085 21699 239113
rect 21485 239023 21513 239051
rect 21547 239023 21575 239051
rect 21609 239023 21637 239051
rect 21671 239023 21699 239051
rect 21485 238961 21513 238989
rect 21547 238961 21575 238989
rect 21609 238961 21637 238989
rect 21671 238961 21699 238989
rect 21485 230147 21513 230175
rect 21547 230147 21575 230175
rect 21609 230147 21637 230175
rect 21671 230147 21699 230175
rect 21485 230085 21513 230113
rect 21547 230085 21575 230113
rect 21609 230085 21637 230113
rect 21671 230085 21699 230113
rect 21485 230023 21513 230051
rect 21547 230023 21575 230051
rect 21609 230023 21637 230051
rect 21671 230023 21699 230051
rect 21485 229961 21513 229989
rect 21547 229961 21575 229989
rect 21609 229961 21637 229989
rect 21671 229961 21699 229989
rect 21485 221147 21513 221175
rect 21547 221147 21575 221175
rect 21609 221147 21637 221175
rect 21671 221147 21699 221175
rect 21485 221085 21513 221113
rect 21547 221085 21575 221113
rect 21609 221085 21637 221113
rect 21671 221085 21699 221113
rect 21485 221023 21513 221051
rect 21547 221023 21575 221051
rect 21609 221023 21637 221051
rect 21671 221023 21699 221051
rect 21485 220961 21513 220989
rect 21547 220961 21575 220989
rect 21609 220961 21637 220989
rect 21671 220961 21699 220989
rect 21485 212147 21513 212175
rect 21547 212147 21575 212175
rect 21609 212147 21637 212175
rect 21671 212147 21699 212175
rect 21485 212085 21513 212113
rect 21547 212085 21575 212113
rect 21609 212085 21637 212113
rect 21671 212085 21699 212113
rect 21485 212023 21513 212051
rect 21547 212023 21575 212051
rect 21609 212023 21637 212051
rect 21671 212023 21699 212051
rect 21485 211961 21513 211989
rect 21547 211961 21575 211989
rect 21609 211961 21637 211989
rect 21671 211961 21699 211989
rect 21485 203147 21513 203175
rect 21547 203147 21575 203175
rect 21609 203147 21637 203175
rect 21671 203147 21699 203175
rect 21485 203085 21513 203113
rect 21547 203085 21575 203113
rect 21609 203085 21637 203113
rect 21671 203085 21699 203113
rect 21485 203023 21513 203051
rect 21547 203023 21575 203051
rect 21609 203023 21637 203051
rect 21671 203023 21699 203051
rect 21485 202961 21513 202989
rect 21547 202961 21575 202989
rect 21609 202961 21637 202989
rect 21671 202961 21699 202989
rect 21485 194147 21513 194175
rect 21547 194147 21575 194175
rect 21609 194147 21637 194175
rect 21671 194147 21699 194175
rect 21485 194085 21513 194113
rect 21547 194085 21575 194113
rect 21609 194085 21637 194113
rect 21671 194085 21699 194113
rect 21485 194023 21513 194051
rect 21547 194023 21575 194051
rect 21609 194023 21637 194051
rect 21671 194023 21699 194051
rect 21485 193961 21513 193989
rect 21547 193961 21575 193989
rect 21609 193961 21637 193989
rect 21671 193961 21699 193989
rect 21485 185147 21513 185175
rect 21547 185147 21575 185175
rect 21609 185147 21637 185175
rect 21671 185147 21699 185175
rect 21485 185085 21513 185113
rect 21547 185085 21575 185113
rect 21609 185085 21637 185113
rect 21671 185085 21699 185113
rect 21485 185023 21513 185051
rect 21547 185023 21575 185051
rect 21609 185023 21637 185051
rect 21671 185023 21699 185051
rect 21485 184961 21513 184989
rect 21547 184961 21575 184989
rect 21609 184961 21637 184989
rect 21671 184961 21699 184989
rect 21485 176147 21513 176175
rect 21547 176147 21575 176175
rect 21609 176147 21637 176175
rect 21671 176147 21699 176175
rect 21485 176085 21513 176113
rect 21547 176085 21575 176113
rect 21609 176085 21637 176113
rect 21671 176085 21699 176113
rect 21485 176023 21513 176051
rect 21547 176023 21575 176051
rect 21609 176023 21637 176051
rect 21671 176023 21699 176051
rect 21485 175961 21513 175989
rect 21547 175961 21575 175989
rect 21609 175961 21637 175989
rect 21671 175961 21699 175989
rect 21485 167147 21513 167175
rect 21547 167147 21575 167175
rect 21609 167147 21637 167175
rect 21671 167147 21699 167175
rect 21485 167085 21513 167113
rect 21547 167085 21575 167113
rect 21609 167085 21637 167113
rect 21671 167085 21699 167113
rect 21485 167023 21513 167051
rect 21547 167023 21575 167051
rect 21609 167023 21637 167051
rect 21671 167023 21699 167051
rect 21485 166961 21513 166989
rect 21547 166961 21575 166989
rect 21609 166961 21637 166989
rect 21671 166961 21699 166989
rect 21485 158147 21513 158175
rect 21547 158147 21575 158175
rect 21609 158147 21637 158175
rect 21671 158147 21699 158175
rect 21485 158085 21513 158113
rect 21547 158085 21575 158113
rect 21609 158085 21637 158113
rect 21671 158085 21699 158113
rect 21485 158023 21513 158051
rect 21547 158023 21575 158051
rect 21609 158023 21637 158051
rect 21671 158023 21699 158051
rect 21485 157961 21513 157989
rect 21547 157961 21575 157989
rect 21609 157961 21637 157989
rect 21671 157961 21699 157989
rect 21485 149147 21513 149175
rect 21547 149147 21575 149175
rect 21609 149147 21637 149175
rect 21671 149147 21699 149175
rect 21485 149085 21513 149113
rect 21547 149085 21575 149113
rect 21609 149085 21637 149113
rect 21671 149085 21699 149113
rect 21485 149023 21513 149051
rect 21547 149023 21575 149051
rect 21609 149023 21637 149051
rect 21671 149023 21699 149051
rect 21485 148961 21513 148989
rect 21547 148961 21575 148989
rect 21609 148961 21637 148989
rect 21671 148961 21699 148989
rect 21485 140147 21513 140175
rect 21547 140147 21575 140175
rect 21609 140147 21637 140175
rect 21671 140147 21699 140175
rect 21485 140085 21513 140113
rect 21547 140085 21575 140113
rect 21609 140085 21637 140113
rect 21671 140085 21699 140113
rect 21485 140023 21513 140051
rect 21547 140023 21575 140051
rect 21609 140023 21637 140051
rect 21671 140023 21699 140051
rect 21485 139961 21513 139989
rect 21547 139961 21575 139989
rect 21609 139961 21637 139989
rect 21671 139961 21699 139989
rect 21485 131147 21513 131175
rect 21547 131147 21575 131175
rect 21609 131147 21637 131175
rect 21671 131147 21699 131175
rect 21485 131085 21513 131113
rect 21547 131085 21575 131113
rect 21609 131085 21637 131113
rect 21671 131085 21699 131113
rect 21485 131023 21513 131051
rect 21547 131023 21575 131051
rect 21609 131023 21637 131051
rect 21671 131023 21699 131051
rect 21485 130961 21513 130989
rect 21547 130961 21575 130989
rect 21609 130961 21637 130989
rect 21671 130961 21699 130989
rect 21485 122147 21513 122175
rect 21547 122147 21575 122175
rect 21609 122147 21637 122175
rect 21671 122147 21699 122175
rect 21485 122085 21513 122113
rect 21547 122085 21575 122113
rect 21609 122085 21637 122113
rect 21671 122085 21699 122113
rect 21485 122023 21513 122051
rect 21547 122023 21575 122051
rect 21609 122023 21637 122051
rect 21671 122023 21699 122051
rect 21485 121961 21513 121989
rect 21547 121961 21575 121989
rect 21609 121961 21637 121989
rect 21671 121961 21699 121989
rect 21485 113147 21513 113175
rect 21547 113147 21575 113175
rect 21609 113147 21637 113175
rect 21671 113147 21699 113175
rect 21485 113085 21513 113113
rect 21547 113085 21575 113113
rect 21609 113085 21637 113113
rect 21671 113085 21699 113113
rect 21485 113023 21513 113051
rect 21547 113023 21575 113051
rect 21609 113023 21637 113051
rect 21671 113023 21699 113051
rect 21485 112961 21513 112989
rect 21547 112961 21575 112989
rect 21609 112961 21637 112989
rect 21671 112961 21699 112989
rect 21485 104147 21513 104175
rect 21547 104147 21575 104175
rect 21609 104147 21637 104175
rect 21671 104147 21699 104175
rect 21485 104085 21513 104113
rect 21547 104085 21575 104113
rect 21609 104085 21637 104113
rect 21671 104085 21699 104113
rect 21485 104023 21513 104051
rect 21547 104023 21575 104051
rect 21609 104023 21637 104051
rect 21671 104023 21699 104051
rect 21485 103961 21513 103989
rect 21547 103961 21575 103989
rect 21609 103961 21637 103989
rect 21671 103961 21699 103989
rect 21485 95147 21513 95175
rect 21547 95147 21575 95175
rect 21609 95147 21637 95175
rect 21671 95147 21699 95175
rect 21485 95085 21513 95113
rect 21547 95085 21575 95113
rect 21609 95085 21637 95113
rect 21671 95085 21699 95113
rect 21485 95023 21513 95051
rect 21547 95023 21575 95051
rect 21609 95023 21637 95051
rect 21671 95023 21699 95051
rect 21485 94961 21513 94989
rect 21547 94961 21575 94989
rect 21609 94961 21637 94989
rect 21671 94961 21699 94989
rect 21485 86147 21513 86175
rect 21547 86147 21575 86175
rect 21609 86147 21637 86175
rect 21671 86147 21699 86175
rect 21485 86085 21513 86113
rect 21547 86085 21575 86113
rect 21609 86085 21637 86113
rect 21671 86085 21699 86113
rect 21485 86023 21513 86051
rect 21547 86023 21575 86051
rect 21609 86023 21637 86051
rect 21671 86023 21699 86051
rect 21485 85961 21513 85989
rect 21547 85961 21575 85989
rect 21609 85961 21637 85989
rect 21671 85961 21699 85989
rect 21485 77147 21513 77175
rect 21547 77147 21575 77175
rect 21609 77147 21637 77175
rect 21671 77147 21699 77175
rect 21485 77085 21513 77113
rect 21547 77085 21575 77113
rect 21609 77085 21637 77113
rect 21671 77085 21699 77113
rect 21485 77023 21513 77051
rect 21547 77023 21575 77051
rect 21609 77023 21637 77051
rect 21671 77023 21699 77051
rect 21485 76961 21513 76989
rect 21547 76961 21575 76989
rect 21609 76961 21637 76989
rect 21671 76961 21699 76989
rect 21485 68147 21513 68175
rect 21547 68147 21575 68175
rect 21609 68147 21637 68175
rect 21671 68147 21699 68175
rect 21485 68085 21513 68113
rect 21547 68085 21575 68113
rect 21609 68085 21637 68113
rect 21671 68085 21699 68113
rect 21485 68023 21513 68051
rect 21547 68023 21575 68051
rect 21609 68023 21637 68051
rect 21671 68023 21699 68051
rect 21485 67961 21513 67989
rect 21547 67961 21575 67989
rect 21609 67961 21637 67989
rect 21671 67961 21699 67989
rect 21485 59147 21513 59175
rect 21547 59147 21575 59175
rect 21609 59147 21637 59175
rect 21671 59147 21699 59175
rect 21485 59085 21513 59113
rect 21547 59085 21575 59113
rect 21609 59085 21637 59113
rect 21671 59085 21699 59113
rect 21485 59023 21513 59051
rect 21547 59023 21575 59051
rect 21609 59023 21637 59051
rect 21671 59023 21699 59051
rect 21485 58961 21513 58989
rect 21547 58961 21575 58989
rect 21609 58961 21637 58989
rect 21671 58961 21699 58989
rect 21485 50147 21513 50175
rect 21547 50147 21575 50175
rect 21609 50147 21637 50175
rect 21671 50147 21699 50175
rect 21485 50085 21513 50113
rect 21547 50085 21575 50113
rect 21609 50085 21637 50113
rect 21671 50085 21699 50113
rect 21485 50023 21513 50051
rect 21547 50023 21575 50051
rect 21609 50023 21637 50051
rect 21671 50023 21699 50051
rect 21485 49961 21513 49989
rect 21547 49961 21575 49989
rect 21609 49961 21637 49989
rect 21671 49961 21699 49989
rect 21485 41147 21513 41175
rect 21547 41147 21575 41175
rect 21609 41147 21637 41175
rect 21671 41147 21699 41175
rect 21485 41085 21513 41113
rect 21547 41085 21575 41113
rect 21609 41085 21637 41113
rect 21671 41085 21699 41113
rect 21485 41023 21513 41051
rect 21547 41023 21575 41051
rect 21609 41023 21637 41051
rect 21671 41023 21699 41051
rect 21485 40961 21513 40989
rect 21547 40961 21575 40989
rect 21609 40961 21637 40989
rect 21671 40961 21699 40989
rect 21485 32147 21513 32175
rect 21547 32147 21575 32175
rect 21609 32147 21637 32175
rect 21671 32147 21699 32175
rect 21485 32085 21513 32113
rect 21547 32085 21575 32113
rect 21609 32085 21637 32113
rect 21671 32085 21699 32113
rect 21485 32023 21513 32051
rect 21547 32023 21575 32051
rect 21609 32023 21637 32051
rect 21671 32023 21699 32051
rect 21485 31961 21513 31989
rect 21547 31961 21575 31989
rect 21609 31961 21637 31989
rect 21671 31961 21699 31989
rect 21485 23147 21513 23175
rect 21547 23147 21575 23175
rect 21609 23147 21637 23175
rect 21671 23147 21699 23175
rect 21485 23085 21513 23113
rect 21547 23085 21575 23113
rect 21609 23085 21637 23113
rect 21671 23085 21699 23113
rect 21485 23023 21513 23051
rect 21547 23023 21575 23051
rect 21609 23023 21637 23051
rect 21671 23023 21699 23051
rect 21485 22961 21513 22989
rect 21547 22961 21575 22989
rect 21609 22961 21637 22989
rect 21671 22961 21699 22989
rect 21485 14147 21513 14175
rect 21547 14147 21575 14175
rect 21609 14147 21637 14175
rect 21671 14147 21699 14175
rect 21485 14085 21513 14113
rect 21547 14085 21575 14113
rect 21609 14085 21637 14113
rect 21671 14085 21699 14113
rect 21485 14023 21513 14051
rect 21547 14023 21575 14051
rect 21609 14023 21637 14051
rect 21671 14023 21699 14051
rect 21485 13961 21513 13989
rect 21547 13961 21575 13989
rect 21609 13961 21637 13989
rect 21671 13961 21699 13989
rect 21485 5147 21513 5175
rect 21547 5147 21575 5175
rect 21609 5147 21637 5175
rect 21671 5147 21699 5175
rect 21485 5085 21513 5113
rect 21547 5085 21575 5113
rect 21609 5085 21637 5113
rect 21671 5085 21699 5113
rect 21485 5023 21513 5051
rect 21547 5023 21575 5051
rect 21609 5023 21637 5051
rect 21671 5023 21699 5051
rect 21485 4961 21513 4989
rect 21547 4961 21575 4989
rect 21609 4961 21637 4989
rect 21671 4961 21699 4989
rect 21485 -588 21513 -560
rect 21547 -588 21575 -560
rect 21609 -588 21637 -560
rect 21671 -588 21699 -560
rect 21485 -650 21513 -622
rect 21547 -650 21575 -622
rect 21609 -650 21637 -622
rect 21671 -650 21699 -622
rect 21485 -712 21513 -684
rect 21547 -712 21575 -684
rect 21609 -712 21637 -684
rect 21671 -712 21699 -684
rect 21485 -774 21513 -746
rect 21547 -774 21575 -746
rect 21609 -774 21637 -746
rect 21671 -774 21699 -746
rect 28625 298578 28653 298606
rect 28687 298578 28715 298606
rect 28749 298578 28777 298606
rect 28811 298578 28839 298606
rect 28625 298516 28653 298544
rect 28687 298516 28715 298544
rect 28749 298516 28777 298544
rect 28811 298516 28839 298544
rect 28625 298454 28653 298482
rect 28687 298454 28715 298482
rect 28749 298454 28777 298482
rect 28811 298454 28839 298482
rect 28625 298392 28653 298420
rect 28687 298392 28715 298420
rect 28749 298392 28777 298420
rect 28811 298392 28839 298420
rect 28625 290147 28653 290175
rect 28687 290147 28715 290175
rect 28749 290147 28777 290175
rect 28811 290147 28839 290175
rect 28625 290085 28653 290113
rect 28687 290085 28715 290113
rect 28749 290085 28777 290113
rect 28811 290085 28839 290113
rect 28625 290023 28653 290051
rect 28687 290023 28715 290051
rect 28749 290023 28777 290051
rect 28811 290023 28839 290051
rect 28625 289961 28653 289989
rect 28687 289961 28715 289989
rect 28749 289961 28777 289989
rect 28811 289961 28839 289989
rect 28625 281147 28653 281175
rect 28687 281147 28715 281175
rect 28749 281147 28777 281175
rect 28811 281147 28839 281175
rect 28625 281085 28653 281113
rect 28687 281085 28715 281113
rect 28749 281085 28777 281113
rect 28811 281085 28839 281113
rect 28625 281023 28653 281051
rect 28687 281023 28715 281051
rect 28749 281023 28777 281051
rect 28811 281023 28839 281051
rect 28625 280961 28653 280989
rect 28687 280961 28715 280989
rect 28749 280961 28777 280989
rect 28811 280961 28839 280989
rect 28625 272147 28653 272175
rect 28687 272147 28715 272175
rect 28749 272147 28777 272175
rect 28811 272147 28839 272175
rect 28625 272085 28653 272113
rect 28687 272085 28715 272113
rect 28749 272085 28777 272113
rect 28811 272085 28839 272113
rect 28625 272023 28653 272051
rect 28687 272023 28715 272051
rect 28749 272023 28777 272051
rect 28811 272023 28839 272051
rect 28625 271961 28653 271989
rect 28687 271961 28715 271989
rect 28749 271961 28777 271989
rect 28811 271961 28839 271989
rect 28625 263147 28653 263175
rect 28687 263147 28715 263175
rect 28749 263147 28777 263175
rect 28811 263147 28839 263175
rect 28625 263085 28653 263113
rect 28687 263085 28715 263113
rect 28749 263085 28777 263113
rect 28811 263085 28839 263113
rect 28625 263023 28653 263051
rect 28687 263023 28715 263051
rect 28749 263023 28777 263051
rect 28811 263023 28839 263051
rect 28625 262961 28653 262989
rect 28687 262961 28715 262989
rect 28749 262961 28777 262989
rect 28811 262961 28839 262989
rect 28625 254147 28653 254175
rect 28687 254147 28715 254175
rect 28749 254147 28777 254175
rect 28811 254147 28839 254175
rect 28625 254085 28653 254113
rect 28687 254085 28715 254113
rect 28749 254085 28777 254113
rect 28811 254085 28839 254113
rect 28625 254023 28653 254051
rect 28687 254023 28715 254051
rect 28749 254023 28777 254051
rect 28811 254023 28839 254051
rect 28625 253961 28653 253989
rect 28687 253961 28715 253989
rect 28749 253961 28777 253989
rect 28811 253961 28839 253989
rect 28625 245147 28653 245175
rect 28687 245147 28715 245175
rect 28749 245147 28777 245175
rect 28811 245147 28839 245175
rect 28625 245085 28653 245113
rect 28687 245085 28715 245113
rect 28749 245085 28777 245113
rect 28811 245085 28839 245113
rect 28625 245023 28653 245051
rect 28687 245023 28715 245051
rect 28749 245023 28777 245051
rect 28811 245023 28839 245051
rect 28625 244961 28653 244989
rect 28687 244961 28715 244989
rect 28749 244961 28777 244989
rect 28811 244961 28839 244989
rect 28625 236147 28653 236175
rect 28687 236147 28715 236175
rect 28749 236147 28777 236175
rect 28811 236147 28839 236175
rect 28625 236085 28653 236113
rect 28687 236085 28715 236113
rect 28749 236085 28777 236113
rect 28811 236085 28839 236113
rect 28625 236023 28653 236051
rect 28687 236023 28715 236051
rect 28749 236023 28777 236051
rect 28811 236023 28839 236051
rect 28625 235961 28653 235989
rect 28687 235961 28715 235989
rect 28749 235961 28777 235989
rect 28811 235961 28839 235989
rect 28625 227147 28653 227175
rect 28687 227147 28715 227175
rect 28749 227147 28777 227175
rect 28811 227147 28839 227175
rect 28625 227085 28653 227113
rect 28687 227085 28715 227113
rect 28749 227085 28777 227113
rect 28811 227085 28839 227113
rect 28625 227023 28653 227051
rect 28687 227023 28715 227051
rect 28749 227023 28777 227051
rect 28811 227023 28839 227051
rect 28625 226961 28653 226989
rect 28687 226961 28715 226989
rect 28749 226961 28777 226989
rect 28811 226961 28839 226989
rect 28625 218147 28653 218175
rect 28687 218147 28715 218175
rect 28749 218147 28777 218175
rect 28811 218147 28839 218175
rect 28625 218085 28653 218113
rect 28687 218085 28715 218113
rect 28749 218085 28777 218113
rect 28811 218085 28839 218113
rect 28625 218023 28653 218051
rect 28687 218023 28715 218051
rect 28749 218023 28777 218051
rect 28811 218023 28839 218051
rect 28625 217961 28653 217989
rect 28687 217961 28715 217989
rect 28749 217961 28777 217989
rect 28811 217961 28839 217989
rect 28625 209147 28653 209175
rect 28687 209147 28715 209175
rect 28749 209147 28777 209175
rect 28811 209147 28839 209175
rect 28625 209085 28653 209113
rect 28687 209085 28715 209113
rect 28749 209085 28777 209113
rect 28811 209085 28839 209113
rect 28625 209023 28653 209051
rect 28687 209023 28715 209051
rect 28749 209023 28777 209051
rect 28811 209023 28839 209051
rect 28625 208961 28653 208989
rect 28687 208961 28715 208989
rect 28749 208961 28777 208989
rect 28811 208961 28839 208989
rect 28625 200147 28653 200175
rect 28687 200147 28715 200175
rect 28749 200147 28777 200175
rect 28811 200147 28839 200175
rect 28625 200085 28653 200113
rect 28687 200085 28715 200113
rect 28749 200085 28777 200113
rect 28811 200085 28839 200113
rect 28625 200023 28653 200051
rect 28687 200023 28715 200051
rect 28749 200023 28777 200051
rect 28811 200023 28839 200051
rect 28625 199961 28653 199989
rect 28687 199961 28715 199989
rect 28749 199961 28777 199989
rect 28811 199961 28839 199989
rect 28625 191147 28653 191175
rect 28687 191147 28715 191175
rect 28749 191147 28777 191175
rect 28811 191147 28839 191175
rect 28625 191085 28653 191113
rect 28687 191085 28715 191113
rect 28749 191085 28777 191113
rect 28811 191085 28839 191113
rect 28625 191023 28653 191051
rect 28687 191023 28715 191051
rect 28749 191023 28777 191051
rect 28811 191023 28839 191051
rect 28625 190961 28653 190989
rect 28687 190961 28715 190989
rect 28749 190961 28777 190989
rect 28811 190961 28839 190989
rect 28625 182147 28653 182175
rect 28687 182147 28715 182175
rect 28749 182147 28777 182175
rect 28811 182147 28839 182175
rect 28625 182085 28653 182113
rect 28687 182085 28715 182113
rect 28749 182085 28777 182113
rect 28811 182085 28839 182113
rect 28625 182023 28653 182051
rect 28687 182023 28715 182051
rect 28749 182023 28777 182051
rect 28811 182023 28839 182051
rect 28625 181961 28653 181989
rect 28687 181961 28715 181989
rect 28749 181961 28777 181989
rect 28811 181961 28839 181989
rect 28625 173147 28653 173175
rect 28687 173147 28715 173175
rect 28749 173147 28777 173175
rect 28811 173147 28839 173175
rect 28625 173085 28653 173113
rect 28687 173085 28715 173113
rect 28749 173085 28777 173113
rect 28811 173085 28839 173113
rect 28625 173023 28653 173051
rect 28687 173023 28715 173051
rect 28749 173023 28777 173051
rect 28811 173023 28839 173051
rect 28625 172961 28653 172989
rect 28687 172961 28715 172989
rect 28749 172961 28777 172989
rect 28811 172961 28839 172989
rect 28625 164147 28653 164175
rect 28687 164147 28715 164175
rect 28749 164147 28777 164175
rect 28811 164147 28839 164175
rect 28625 164085 28653 164113
rect 28687 164085 28715 164113
rect 28749 164085 28777 164113
rect 28811 164085 28839 164113
rect 28625 164023 28653 164051
rect 28687 164023 28715 164051
rect 28749 164023 28777 164051
rect 28811 164023 28839 164051
rect 28625 163961 28653 163989
rect 28687 163961 28715 163989
rect 28749 163961 28777 163989
rect 28811 163961 28839 163989
rect 28625 155147 28653 155175
rect 28687 155147 28715 155175
rect 28749 155147 28777 155175
rect 28811 155147 28839 155175
rect 28625 155085 28653 155113
rect 28687 155085 28715 155113
rect 28749 155085 28777 155113
rect 28811 155085 28839 155113
rect 28625 155023 28653 155051
rect 28687 155023 28715 155051
rect 28749 155023 28777 155051
rect 28811 155023 28839 155051
rect 28625 154961 28653 154989
rect 28687 154961 28715 154989
rect 28749 154961 28777 154989
rect 28811 154961 28839 154989
rect 28625 146147 28653 146175
rect 28687 146147 28715 146175
rect 28749 146147 28777 146175
rect 28811 146147 28839 146175
rect 28625 146085 28653 146113
rect 28687 146085 28715 146113
rect 28749 146085 28777 146113
rect 28811 146085 28839 146113
rect 28625 146023 28653 146051
rect 28687 146023 28715 146051
rect 28749 146023 28777 146051
rect 28811 146023 28839 146051
rect 28625 145961 28653 145989
rect 28687 145961 28715 145989
rect 28749 145961 28777 145989
rect 28811 145961 28839 145989
rect 28625 137147 28653 137175
rect 28687 137147 28715 137175
rect 28749 137147 28777 137175
rect 28811 137147 28839 137175
rect 28625 137085 28653 137113
rect 28687 137085 28715 137113
rect 28749 137085 28777 137113
rect 28811 137085 28839 137113
rect 28625 137023 28653 137051
rect 28687 137023 28715 137051
rect 28749 137023 28777 137051
rect 28811 137023 28839 137051
rect 28625 136961 28653 136989
rect 28687 136961 28715 136989
rect 28749 136961 28777 136989
rect 28811 136961 28839 136989
rect 28625 128147 28653 128175
rect 28687 128147 28715 128175
rect 28749 128147 28777 128175
rect 28811 128147 28839 128175
rect 28625 128085 28653 128113
rect 28687 128085 28715 128113
rect 28749 128085 28777 128113
rect 28811 128085 28839 128113
rect 28625 128023 28653 128051
rect 28687 128023 28715 128051
rect 28749 128023 28777 128051
rect 28811 128023 28839 128051
rect 28625 127961 28653 127989
rect 28687 127961 28715 127989
rect 28749 127961 28777 127989
rect 28811 127961 28839 127989
rect 28625 119147 28653 119175
rect 28687 119147 28715 119175
rect 28749 119147 28777 119175
rect 28811 119147 28839 119175
rect 28625 119085 28653 119113
rect 28687 119085 28715 119113
rect 28749 119085 28777 119113
rect 28811 119085 28839 119113
rect 28625 119023 28653 119051
rect 28687 119023 28715 119051
rect 28749 119023 28777 119051
rect 28811 119023 28839 119051
rect 28625 118961 28653 118989
rect 28687 118961 28715 118989
rect 28749 118961 28777 118989
rect 28811 118961 28839 118989
rect 28625 110147 28653 110175
rect 28687 110147 28715 110175
rect 28749 110147 28777 110175
rect 28811 110147 28839 110175
rect 28625 110085 28653 110113
rect 28687 110085 28715 110113
rect 28749 110085 28777 110113
rect 28811 110085 28839 110113
rect 28625 110023 28653 110051
rect 28687 110023 28715 110051
rect 28749 110023 28777 110051
rect 28811 110023 28839 110051
rect 28625 109961 28653 109989
rect 28687 109961 28715 109989
rect 28749 109961 28777 109989
rect 28811 109961 28839 109989
rect 28625 101147 28653 101175
rect 28687 101147 28715 101175
rect 28749 101147 28777 101175
rect 28811 101147 28839 101175
rect 28625 101085 28653 101113
rect 28687 101085 28715 101113
rect 28749 101085 28777 101113
rect 28811 101085 28839 101113
rect 28625 101023 28653 101051
rect 28687 101023 28715 101051
rect 28749 101023 28777 101051
rect 28811 101023 28839 101051
rect 28625 100961 28653 100989
rect 28687 100961 28715 100989
rect 28749 100961 28777 100989
rect 28811 100961 28839 100989
rect 28625 92147 28653 92175
rect 28687 92147 28715 92175
rect 28749 92147 28777 92175
rect 28811 92147 28839 92175
rect 28625 92085 28653 92113
rect 28687 92085 28715 92113
rect 28749 92085 28777 92113
rect 28811 92085 28839 92113
rect 28625 92023 28653 92051
rect 28687 92023 28715 92051
rect 28749 92023 28777 92051
rect 28811 92023 28839 92051
rect 28625 91961 28653 91989
rect 28687 91961 28715 91989
rect 28749 91961 28777 91989
rect 28811 91961 28839 91989
rect 28625 83147 28653 83175
rect 28687 83147 28715 83175
rect 28749 83147 28777 83175
rect 28811 83147 28839 83175
rect 28625 83085 28653 83113
rect 28687 83085 28715 83113
rect 28749 83085 28777 83113
rect 28811 83085 28839 83113
rect 28625 83023 28653 83051
rect 28687 83023 28715 83051
rect 28749 83023 28777 83051
rect 28811 83023 28839 83051
rect 28625 82961 28653 82989
rect 28687 82961 28715 82989
rect 28749 82961 28777 82989
rect 28811 82961 28839 82989
rect 28625 74147 28653 74175
rect 28687 74147 28715 74175
rect 28749 74147 28777 74175
rect 28811 74147 28839 74175
rect 28625 74085 28653 74113
rect 28687 74085 28715 74113
rect 28749 74085 28777 74113
rect 28811 74085 28839 74113
rect 28625 74023 28653 74051
rect 28687 74023 28715 74051
rect 28749 74023 28777 74051
rect 28811 74023 28839 74051
rect 28625 73961 28653 73989
rect 28687 73961 28715 73989
rect 28749 73961 28777 73989
rect 28811 73961 28839 73989
rect 28625 65147 28653 65175
rect 28687 65147 28715 65175
rect 28749 65147 28777 65175
rect 28811 65147 28839 65175
rect 28625 65085 28653 65113
rect 28687 65085 28715 65113
rect 28749 65085 28777 65113
rect 28811 65085 28839 65113
rect 28625 65023 28653 65051
rect 28687 65023 28715 65051
rect 28749 65023 28777 65051
rect 28811 65023 28839 65051
rect 28625 64961 28653 64989
rect 28687 64961 28715 64989
rect 28749 64961 28777 64989
rect 28811 64961 28839 64989
rect 28625 56147 28653 56175
rect 28687 56147 28715 56175
rect 28749 56147 28777 56175
rect 28811 56147 28839 56175
rect 28625 56085 28653 56113
rect 28687 56085 28715 56113
rect 28749 56085 28777 56113
rect 28811 56085 28839 56113
rect 28625 56023 28653 56051
rect 28687 56023 28715 56051
rect 28749 56023 28777 56051
rect 28811 56023 28839 56051
rect 28625 55961 28653 55989
rect 28687 55961 28715 55989
rect 28749 55961 28777 55989
rect 28811 55961 28839 55989
rect 28625 47147 28653 47175
rect 28687 47147 28715 47175
rect 28749 47147 28777 47175
rect 28811 47147 28839 47175
rect 28625 47085 28653 47113
rect 28687 47085 28715 47113
rect 28749 47085 28777 47113
rect 28811 47085 28839 47113
rect 28625 47023 28653 47051
rect 28687 47023 28715 47051
rect 28749 47023 28777 47051
rect 28811 47023 28839 47051
rect 28625 46961 28653 46989
rect 28687 46961 28715 46989
rect 28749 46961 28777 46989
rect 28811 46961 28839 46989
rect 28625 38147 28653 38175
rect 28687 38147 28715 38175
rect 28749 38147 28777 38175
rect 28811 38147 28839 38175
rect 28625 38085 28653 38113
rect 28687 38085 28715 38113
rect 28749 38085 28777 38113
rect 28811 38085 28839 38113
rect 28625 38023 28653 38051
rect 28687 38023 28715 38051
rect 28749 38023 28777 38051
rect 28811 38023 28839 38051
rect 28625 37961 28653 37989
rect 28687 37961 28715 37989
rect 28749 37961 28777 37989
rect 28811 37961 28839 37989
rect 28625 29147 28653 29175
rect 28687 29147 28715 29175
rect 28749 29147 28777 29175
rect 28811 29147 28839 29175
rect 28625 29085 28653 29113
rect 28687 29085 28715 29113
rect 28749 29085 28777 29113
rect 28811 29085 28839 29113
rect 28625 29023 28653 29051
rect 28687 29023 28715 29051
rect 28749 29023 28777 29051
rect 28811 29023 28839 29051
rect 28625 28961 28653 28989
rect 28687 28961 28715 28989
rect 28749 28961 28777 28989
rect 28811 28961 28839 28989
rect 28625 20147 28653 20175
rect 28687 20147 28715 20175
rect 28749 20147 28777 20175
rect 28811 20147 28839 20175
rect 28625 20085 28653 20113
rect 28687 20085 28715 20113
rect 28749 20085 28777 20113
rect 28811 20085 28839 20113
rect 28625 20023 28653 20051
rect 28687 20023 28715 20051
rect 28749 20023 28777 20051
rect 28811 20023 28839 20051
rect 28625 19961 28653 19989
rect 28687 19961 28715 19989
rect 28749 19961 28777 19989
rect 28811 19961 28839 19989
rect 28625 11147 28653 11175
rect 28687 11147 28715 11175
rect 28749 11147 28777 11175
rect 28811 11147 28839 11175
rect 28625 11085 28653 11113
rect 28687 11085 28715 11113
rect 28749 11085 28777 11113
rect 28811 11085 28839 11113
rect 28625 11023 28653 11051
rect 28687 11023 28715 11051
rect 28749 11023 28777 11051
rect 28811 11023 28839 11051
rect 28625 10961 28653 10989
rect 28687 10961 28715 10989
rect 28749 10961 28777 10989
rect 28811 10961 28839 10989
rect 28625 2147 28653 2175
rect 28687 2147 28715 2175
rect 28749 2147 28777 2175
rect 28811 2147 28839 2175
rect 28625 2085 28653 2113
rect 28687 2085 28715 2113
rect 28749 2085 28777 2113
rect 28811 2085 28839 2113
rect 28625 2023 28653 2051
rect 28687 2023 28715 2051
rect 28749 2023 28777 2051
rect 28811 2023 28839 2051
rect 28625 1961 28653 1989
rect 28687 1961 28715 1989
rect 28749 1961 28777 1989
rect 28811 1961 28839 1989
rect 28625 -108 28653 -80
rect 28687 -108 28715 -80
rect 28749 -108 28777 -80
rect 28811 -108 28839 -80
rect 28625 -170 28653 -142
rect 28687 -170 28715 -142
rect 28749 -170 28777 -142
rect 28811 -170 28839 -142
rect 28625 -232 28653 -204
rect 28687 -232 28715 -204
rect 28749 -232 28777 -204
rect 28811 -232 28839 -204
rect 28625 -294 28653 -266
rect 28687 -294 28715 -266
rect 28749 -294 28777 -266
rect 28811 -294 28839 -266
rect 30485 299058 30513 299086
rect 30547 299058 30575 299086
rect 30609 299058 30637 299086
rect 30671 299058 30699 299086
rect 30485 298996 30513 299024
rect 30547 298996 30575 299024
rect 30609 298996 30637 299024
rect 30671 298996 30699 299024
rect 30485 298934 30513 298962
rect 30547 298934 30575 298962
rect 30609 298934 30637 298962
rect 30671 298934 30699 298962
rect 30485 298872 30513 298900
rect 30547 298872 30575 298900
rect 30609 298872 30637 298900
rect 30671 298872 30699 298900
rect 30485 293147 30513 293175
rect 30547 293147 30575 293175
rect 30609 293147 30637 293175
rect 30671 293147 30699 293175
rect 30485 293085 30513 293113
rect 30547 293085 30575 293113
rect 30609 293085 30637 293113
rect 30671 293085 30699 293113
rect 30485 293023 30513 293051
rect 30547 293023 30575 293051
rect 30609 293023 30637 293051
rect 30671 293023 30699 293051
rect 30485 292961 30513 292989
rect 30547 292961 30575 292989
rect 30609 292961 30637 292989
rect 30671 292961 30699 292989
rect 30485 284147 30513 284175
rect 30547 284147 30575 284175
rect 30609 284147 30637 284175
rect 30671 284147 30699 284175
rect 30485 284085 30513 284113
rect 30547 284085 30575 284113
rect 30609 284085 30637 284113
rect 30671 284085 30699 284113
rect 30485 284023 30513 284051
rect 30547 284023 30575 284051
rect 30609 284023 30637 284051
rect 30671 284023 30699 284051
rect 30485 283961 30513 283989
rect 30547 283961 30575 283989
rect 30609 283961 30637 283989
rect 30671 283961 30699 283989
rect 30485 275147 30513 275175
rect 30547 275147 30575 275175
rect 30609 275147 30637 275175
rect 30671 275147 30699 275175
rect 30485 275085 30513 275113
rect 30547 275085 30575 275113
rect 30609 275085 30637 275113
rect 30671 275085 30699 275113
rect 30485 275023 30513 275051
rect 30547 275023 30575 275051
rect 30609 275023 30637 275051
rect 30671 275023 30699 275051
rect 30485 274961 30513 274989
rect 30547 274961 30575 274989
rect 30609 274961 30637 274989
rect 30671 274961 30699 274989
rect 30485 266147 30513 266175
rect 30547 266147 30575 266175
rect 30609 266147 30637 266175
rect 30671 266147 30699 266175
rect 30485 266085 30513 266113
rect 30547 266085 30575 266113
rect 30609 266085 30637 266113
rect 30671 266085 30699 266113
rect 30485 266023 30513 266051
rect 30547 266023 30575 266051
rect 30609 266023 30637 266051
rect 30671 266023 30699 266051
rect 30485 265961 30513 265989
rect 30547 265961 30575 265989
rect 30609 265961 30637 265989
rect 30671 265961 30699 265989
rect 30485 257147 30513 257175
rect 30547 257147 30575 257175
rect 30609 257147 30637 257175
rect 30671 257147 30699 257175
rect 30485 257085 30513 257113
rect 30547 257085 30575 257113
rect 30609 257085 30637 257113
rect 30671 257085 30699 257113
rect 30485 257023 30513 257051
rect 30547 257023 30575 257051
rect 30609 257023 30637 257051
rect 30671 257023 30699 257051
rect 30485 256961 30513 256989
rect 30547 256961 30575 256989
rect 30609 256961 30637 256989
rect 30671 256961 30699 256989
rect 30485 248147 30513 248175
rect 30547 248147 30575 248175
rect 30609 248147 30637 248175
rect 30671 248147 30699 248175
rect 30485 248085 30513 248113
rect 30547 248085 30575 248113
rect 30609 248085 30637 248113
rect 30671 248085 30699 248113
rect 30485 248023 30513 248051
rect 30547 248023 30575 248051
rect 30609 248023 30637 248051
rect 30671 248023 30699 248051
rect 30485 247961 30513 247989
rect 30547 247961 30575 247989
rect 30609 247961 30637 247989
rect 30671 247961 30699 247989
rect 30485 239147 30513 239175
rect 30547 239147 30575 239175
rect 30609 239147 30637 239175
rect 30671 239147 30699 239175
rect 30485 239085 30513 239113
rect 30547 239085 30575 239113
rect 30609 239085 30637 239113
rect 30671 239085 30699 239113
rect 30485 239023 30513 239051
rect 30547 239023 30575 239051
rect 30609 239023 30637 239051
rect 30671 239023 30699 239051
rect 30485 238961 30513 238989
rect 30547 238961 30575 238989
rect 30609 238961 30637 238989
rect 30671 238961 30699 238989
rect 30485 230147 30513 230175
rect 30547 230147 30575 230175
rect 30609 230147 30637 230175
rect 30671 230147 30699 230175
rect 30485 230085 30513 230113
rect 30547 230085 30575 230113
rect 30609 230085 30637 230113
rect 30671 230085 30699 230113
rect 30485 230023 30513 230051
rect 30547 230023 30575 230051
rect 30609 230023 30637 230051
rect 30671 230023 30699 230051
rect 30485 229961 30513 229989
rect 30547 229961 30575 229989
rect 30609 229961 30637 229989
rect 30671 229961 30699 229989
rect 30485 221147 30513 221175
rect 30547 221147 30575 221175
rect 30609 221147 30637 221175
rect 30671 221147 30699 221175
rect 30485 221085 30513 221113
rect 30547 221085 30575 221113
rect 30609 221085 30637 221113
rect 30671 221085 30699 221113
rect 30485 221023 30513 221051
rect 30547 221023 30575 221051
rect 30609 221023 30637 221051
rect 30671 221023 30699 221051
rect 30485 220961 30513 220989
rect 30547 220961 30575 220989
rect 30609 220961 30637 220989
rect 30671 220961 30699 220989
rect 30485 212147 30513 212175
rect 30547 212147 30575 212175
rect 30609 212147 30637 212175
rect 30671 212147 30699 212175
rect 30485 212085 30513 212113
rect 30547 212085 30575 212113
rect 30609 212085 30637 212113
rect 30671 212085 30699 212113
rect 30485 212023 30513 212051
rect 30547 212023 30575 212051
rect 30609 212023 30637 212051
rect 30671 212023 30699 212051
rect 30485 211961 30513 211989
rect 30547 211961 30575 211989
rect 30609 211961 30637 211989
rect 30671 211961 30699 211989
rect 30485 203147 30513 203175
rect 30547 203147 30575 203175
rect 30609 203147 30637 203175
rect 30671 203147 30699 203175
rect 30485 203085 30513 203113
rect 30547 203085 30575 203113
rect 30609 203085 30637 203113
rect 30671 203085 30699 203113
rect 30485 203023 30513 203051
rect 30547 203023 30575 203051
rect 30609 203023 30637 203051
rect 30671 203023 30699 203051
rect 30485 202961 30513 202989
rect 30547 202961 30575 202989
rect 30609 202961 30637 202989
rect 30671 202961 30699 202989
rect 30485 194147 30513 194175
rect 30547 194147 30575 194175
rect 30609 194147 30637 194175
rect 30671 194147 30699 194175
rect 30485 194085 30513 194113
rect 30547 194085 30575 194113
rect 30609 194085 30637 194113
rect 30671 194085 30699 194113
rect 30485 194023 30513 194051
rect 30547 194023 30575 194051
rect 30609 194023 30637 194051
rect 30671 194023 30699 194051
rect 30485 193961 30513 193989
rect 30547 193961 30575 193989
rect 30609 193961 30637 193989
rect 30671 193961 30699 193989
rect 30485 185147 30513 185175
rect 30547 185147 30575 185175
rect 30609 185147 30637 185175
rect 30671 185147 30699 185175
rect 30485 185085 30513 185113
rect 30547 185085 30575 185113
rect 30609 185085 30637 185113
rect 30671 185085 30699 185113
rect 30485 185023 30513 185051
rect 30547 185023 30575 185051
rect 30609 185023 30637 185051
rect 30671 185023 30699 185051
rect 30485 184961 30513 184989
rect 30547 184961 30575 184989
rect 30609 184961 30637 184989
rect 30671 184961 30699 184989
rect 30485 176147 30513 176175
rect 30547 176147 30575 176175
rect 30609 176147 30637 176175
rect 30671 176147 30699 176175
rect 30485 176085 30513 176113
rect 30547 176085 30575 176113
rect 30609 176085 30637 176113
rect 30671 176085 30699 176113
rect 30485 176023 30513 176051
rect 30547 176023 30575 176051
rect 30609 176023 30637 176051
rect 30671 176023 30699 176051
rect 30485 175961 30513 175989
rect 30547 175961 30575 175989
rect 30609 175961 30637 175989
rect 30671 175961 30699 175989
rect 30485 167147 30513 167175
rect 30547 167147 30575 167175
rect 30609 167147 30637 167175
rect 30671 167147 30699 167175
rect 30485 167085 30513 167113
rect 30547 167085 30575 167113
rect 30609 167085 30637 167113
rect 30671 167085 30699 167113
rect 30485 167023 30513 167051
rect 30547 167023 30575 167051
rect 30609 167023 30637 167051
rect 30671 167023 30699 167051
rect 30485 166961 30513 166989
rect 30547 166961 30575 166989
rect 30609 166961 30637 166989
rect 30671 166961 30699 166989
rect 30485 158147 30513 158175
rect 30547 158147 30575 158175
rect 30609 158147 30637 158175
rect 30671 158147 30699 158175
rect 30485 158085 30513 158113
rect 30547 158085 30575 158113
rect 30609 158085 30637 158113
rect 30671 158085 30699 158113
rect 30485 158023 30513 158051
rect 30547 158023 30575 158051
rect 30609 158023 30637 158051
rect 30671 158023 30699 158051
rect 30485 157961 30513 157989
rect 30547 157961 30575 157989
rect 30609 157961 30637 157989
rect 30671 157961 30699 157989
rect 30485 149147 30513 149175
rect 30547 149147 30575 149175
rect 30609 149147 30637 149175
rect 30671 149147 30699 149175
rect 30485 149085 30513 149113
rect 30547 149085 30575 149113
rect 30609 149085 30637 149113
rect 30671 149085 30699 149113
rect 30485 149023 30513 149051
rect 30547 149023 30575 149051
rect 30609 149023 30637 149051
rect 30671 149023 30699 149051
rect 30485 148961 30513 148989
rect 30547 148961 30575 148989
rect 30609 148961 30637 148989
rect 30671 148961 30699 148989
rect 30485 140147 30513 140175
rect 30547 140147 30575 140175
rect 30609 140147 30637 140175
rect 30671 140147 30699 140175
rect 30485 140085 30513 140113
rect 30547 140085 30575 140113
rect 30609 140085 30637 140113
rect 30671 140085 30699 140113
rect 30485 140023 30513 140051
rect 30547 140023 30575 140051
rect 30609 140023 30637 140051
rect 30671 140023 30699 140051
rect 30485 139961 30513 139989
rect 30547 139961 30575 139989
rect 30609 139961 30637 139989
rect 30671 139961 30699 139989
rect 30485 131147 30513 131175
rect 30547 131147 30575 131175
rect 30609 131147 30637 131175
rect 30671 131147 30699 131175
rect 30485 131085 30513 131113
rect 30547 131085 30575 131113
rect 30609 131085 30637 131113
rect 30671 131085 30699 131113
rect 30485 131023 30513 131051
rect 30547 131023 30575 131051
rect 30609 131023 30637 131051
rect 30671 131023 30699 131051
rect 30485 130961 30513 130989
rect 30547 130961 30575 130989
rect 30609 130961 30637 130989
rect 30671 130961 30699 130989
rect 30485 122147 30513 122175
rect 30547 122147 30575 122175
rect 30609 122147 30637 122175
rect 30671 122147 30699 122175
rect 30485 122085 30513 122113
rect 30547 122085 30575 122113
rect 30609 122085 30637 122113
rect 30671 122085 30699 122113
rect 30485 122023 30513 122051
rect 30547 122023 30575 122051
rect 30609 122023 30637 122051
rect 30671 122023 30699 122051
rect 30485 121961 30513 121989
rect 30547 121961 30575 121989
rect 30609 121961 30637 121989
rect 30671 121961 30699 121989
rect 30485 113147 30513 113175
rect 30547 113147 30575 113175
rect 30609 113147 30637 113175
rect 30671 113147 30699 113175
rect 30485 113085 30513 113113
rect 30547 113085 30575 113113
rect 30609 113085 30637 113113
rect 30671 113085 30699 113113
rect 30485 113023 30513 113051
rect 30547 113023 30575 113051
rect 30609 113023 30637 113051
rect 30671 113023 30699 113051
rect 30485 112961 30513 112989
rect 30547 112961 30575 112989
rect 30609 112961 30637 112989
rect 30671 112961 30699 112989
rect 30485 104147 30513 104175
rect 30547 104147 30575 104175
rect 30609 104147 30637 104175
rect 30671 104147 30699 104175
rect 30485 104085 30513 104113
rect 30547 104085 30575 104113
rect 30609 104085 30637 104113
rect 30671 104085 30699 104113
rect 30485 104023 30513 104051
rect 30547 104023 30575 104051
rect 30609 104023 30637 104051
rect 30671 104023 30699 104051
rect 30485 103961 30513 103989
rect 30547 103961 30575 103989
rect 30609 103961 30637 103989
rect 30671 103961 30699 103989
rect 30485 95147 30513 95175
rect 30547 95147 30575 95175
rect 30609 95147 30637 95175
rect 30671 95147 30699 95175
rect 30485 95085 30513 95113
rect 30547 95085 30575 95113
rect 30609 95085 30637 95113
rect 30671 95085 30699 95113
rect 30485 95023 30513 95051
rect 30547 95023 30575 95051
rect 30609 95023 30637 95051
rect 30671 95023 30699 95051
rect 30485 94961 30513 94989
rect 30547 94961 30575 94989
rect 30609 94961 30637 94989
rect 30671 94961 30699 94989
rect 30485 86147 30513 86175
rect 30547 86147 30575 86175
rect 30609 86147 30637 86175
rect 30671 86147 30699 86175
rect 30485 86085 30513 86113
rect 30547 86085 30575 86113
rect 30609 86085 30637 86113
rect 30671 86085 30699 86113
rect 30485 86023 30513 86051
rect 30547 86023 30575 86051
rect 30609 86023 30637 86051
rect 30671 86023 30699 86051
rect 30485 85961 30513 85989
rect 30547 85961 30575 85989
rect 30609 85961 30637 85989
rect 30671 85961 30699 85989
rect 30485 77147 30513 77175
rect 30547 77147 30575 77175
rect 30609 77147 30637 77175
rect 30671 77147 30699 77175
rect 30485 77085 30513 77113
rect 30547 77085 30575 77113
rect 30609 77085 30637 77113
rect 30671 77085 30699 77113
rect 30485 77023 30513 77051
rect 30547 77023 30575 77051
rect 30609 77023 30637 77051
rect 30671 77023 30699 77051
rect 30485 76961 30513 76989
rect 30547 76961 30575 76989
rect 30609 76961 30637 76989
rect 30671 76961 30699 76989
rect 30485 68147 30513 68175
rect 30547 68147 30575 68175
rect 30609 68147 30637 68175
rect 30671 68147 30699 68175
rect 30485 68085 30513 68113
rect 30547 68085 30575 68113
rect 30609 68085 30637 68113
rect 30671 68085 30699 68113
rect 30485 68023 30513 68051
rect 30547 68023 30575 68051
rect 30609 68023 30637 68051
rect 30671 68023 30699 68051
rect 30485 67961 30513 67989
rect 30547 67961 30575 67989
rect 30609 67961 30637 67989
rect 30671 67961 30699 67989
rect 30485 59147 30513 59175
rect 30547 59147 30575 59175
rect 30609 59147 30637 59175
rect 30671 59147 30699 59175
rect 30485 59085 30513 59113
rect 30547 59085 30575 59113
rect 30609 59085 30637 59113
rect 30671 59085 30699 59113
rect 30485 59023 30513 59051
rect 30547 59023 30575 59051
rect 30609 59023 30637 59051
rect 30671 59023 30699 59051
rect 30485 58961 30513 58989
rect 30547 58961 30575 58989
rect 30609 58961 30637 58989
rect 30671 58961 30699 58989
rect 30485 50147 30513 50175
rect 30547 50147 30575 50175
rect 30609 50147 30637 50175
rect 30671 50147 30699 50175
rect 30485 50085 30513 50113
rect 30547 50085 30575 50113
rect 30609 50085 30637 50113
rect 30671 50085 30699 50113
rect 30485 50023 30513 50051
rect 30547 50023 30575 50051
rect 30609 50023 30637 50051
rect 30671 50023 30699 50051
rect 30485 49961 30513 49989
rect 30547 49961 30575 49989
rect 30609 49961 30637 49989
rect 30671 49961 30699 49989
rect 30485 41147 30513 41175
rect 30547 41147 30575 41175
rect 30609 41147 30637 41175
rect 30671 41147 30699 41175
rect 30485 41085 30513 41113
rect 30547 41085 30575 41113
rect 30609 41085 30637 41113
rect 30671 41085 30699 41113
rect 30485 41023 30513 41051
rect 30547 41023 30575 41051
rect 30609 41023 30637 41051
rect 30671 41023 30699 41051
rect 30485 40961 30513 40989
rect 30547 40961 30575 40989
rect 30609 40961 30637 40989
rect 30671 40961 30699 40989
rect 30485 32147 30513 32175
rect 30547 32147 30575 32175
rect 30609 32147 30637 32175
rect 30671 32147 30699 32175
rect 30485 32085 30513 32113
rect 30547 32085 30575 32113
rect 30609 32085 30637 32113
rect 30671 32085 30699 32113
rect 30485 32023 30513 32051
rect 30547 32023 30575 32051
rect 30609 32023 30637 32051
rect 30671 32023 30699 32051
rect 30485 31961 30513 31989
rect 30547 31961 30575 31989
rect 30609 31961 30637 31989
rect 30671 31961 30699 31989
rect 30485 23147 30513 23175
rect 30547 23147 30575 23175
rect 30609 23147 30637 23175
rect 30671 23147 30699 23175
rect 30485 23085 30513 23113
rect 30547 23085 30575 23113
rect 30609 23085 30637 23113
rect 30671 23085 30699 23113
rect 30485 23023 30513 23051
rect 30547 23023 30575 23051
rect 30609 23023 30637 23051
rect 30671 23023 30699 23051
rect 30485 22961 30513 22989
rect 30547 22961 30575 22989
rect 30609 22961 30637 22989
rect 30671 22961 30699 22989
rect 30485 14147 30513 14175
rect 30547 14147 30575 14175
rect 30609 14147 30637 14175
rect 30671 14147 30699 14175
rect 30485 14085 30513 14113
rect 30547 14085 30575 14113
rect 30609 14085 30637 14113
rect 30671 14085 30699 14113
rect 30485 14023 30513 14051
rect 30547 14023 30575 14051
rect 30609 14023 30637 14051
rect 30671 14023 30699 14051
rect 30485 13961 30513 13989
rect 30547 13961 30575 13989
rect 30609 13961 30637 13989
rect 30671 13961 30699 13989
rect 30485 5147 30513 5175
rect 30547 5147 30575 5175
rect 30609 5147 30637 5175
rect 30671 5147 30699 5175
rect 30485 5085 30513 5113
rect 30547 5085 30575 5113
rect 30609 5085 30637 5113
rect 30671 5085 30699 5113
rect 30485 5023 30513 5051
rect 30547 5023 30575 5051
rect 30609 5023 30637 5051
rect 30671 5023 30699 5051
rect 30485 4961 30513 4989
rect 30547 4961 30575 4989
rect 30609 4961 30637 4989
rect 30671 4961 30699 4989
rect 30485 -588 30513 -560
rect 30547 -588 30575 -560
rect 30609 -588 30637 -560
rect 30671 -588 30699 -560
rect 30485 -650 30513 -622
rect 30547 -650 30575 -622
rect 30609 -650 30637 -622
rect 30671 -650 30699 -622
rect 30485 -712 30513 -684
rect 30547 -712 30575 -684
rect 30609 -712 30637 -684
rect 30671 -712 30699 -684
rect 30485 -774 30513 -746
rect 30547 -774 30575 -746
rect 30609 -774 30637 -746
rect 30671 -774 30699 -746
rect 37625 298578 37653 298606
rect 37687 298578 37715 298606
rect 37749 298578 37777 298606
rect 37811 298578 37839 298606
rect 37625 298516 37653 298544
rect 37687 298516 37715 298544
rect 37749 298516 37777 298544
rect 37811 298516 37839 298544
rect 37625 298454 37653 298482
rect 37687 298454 37715 298482
rect 37749 298454 37777 298482
rect 37811 298454 37839 298482
rect 37625 298392 37653 298420
rect 37687 298392 37715 298420
rect 37749 298392 37777 298420
rect 37811 298392 37839 298420
rect 37625 290147 37653 290175
rect 37687 290147 37715 290175
rect 37749 290147 37777 290175
rect 37811 290147 37839 290175
rect 37625 290085 37653 290113
rect 37687 290085 37715 290113
rect 37749 290085 37777 290113
rect 37811 290085 37839 290113
rect 37625 290023 37653 290051
rect 37687 290023 37715 290051
rect 37749 290023 37777 290051
rect 37811 290023 37839 290051
rect 37625 289961 37653 289989
rect 37687 289961 37715 289989
rect 37749 289961 37777 289989
rect 37811 289961 37839 289989
rect 37625 281147 37653 281175
rect 37687 281147 37715 281175
rect 37749 281147 37777 281175
rect 37811 281147 37839 281175
rect 37625 281085 37653 281113
rect 37687 281085 37715 281113
rect 37749 281085 37777 281113
rect 37811 281085 37839 281113
rect 37625 281023 37653 281051
rect 37687 281023 37715 281051
rect 37749 281023 37777 281051
rect 37811 281023 37839 281051
rect 37625 280961 37653 280989
rect 37687 280961 37715 280989
rect 37749 280961 37777 280989
rect 37811 280961 37839 280989
rect 37625 272147 37653 272175
rect 37687 272147 37715 272175
rect 37749 272147 37777 272175
rect 37811 272147 37839 272175
rect 37625 272085 37653 272113
rect 37687 272085 37715 272113
rect 37749 272085 37777 272113
rect 37811 272085 37839 272113
rect 37625 272023 37653 272051
rect 37687 272023 37715 272051
rect 37749 272023 37777 272051
rect 37811 272023 37839 272051
rect 37625 271961 37653 271989
rect 37687 271961 37715 271989
rect 37749 271961 37777 271989
rect 37811 271961 37839 271989
rect 37625 263147 37653 263175
rect 37687 263147 37715 263175
rect 37749 263147 37777 263175
rect 37811 263147 37839 263175
rect 37625 263085 37653 263113
rect 37687 263085 37715 263113
rect 37749 263085 37777 263113
rect 37811 263085 37839 263113
rect 37625 263023 37653 263051
rect 37687 263023 37715 263051
rect 37749 263023 37777 263051
rect 37811 263023 37839 263051
rect 37625 262961 37653 262989
rect 37687 262961 37715 262989
rect 37749 262961 37777 262989
rect 37811 262961 37839 262989
rect 37625 254147 37653 254175
rect 37687 254147 37715 254175
rect 37749 254147 37777 254175
rect 37811 254147 37839 254175
rect 37625 254085 37653 254113
rect 37687 254085 37715 254113
rect 37749 254085 37777 254113
rect 37811 254085 37839 254113
rect 37625 254023 37653 254051
rect 37687 254023 37715 254051
rect 37749 254023 37777 254051
rect 37811 254023 37839 254051
rect 37625 253961 37653 253989
rect 37687 253961 37715 253989
rect 37749 253961 37777 253989
rect 37811 253961 37839 253989
rect 37625 245147 37653 245175
rect 37687 245147 37715 245175
rect 37749 245147 37777 245175
rect 37811 245147 37839 245175
rect 37625 245085 37653 245113
rect 37687 245085 37715 245113
rect 37749 245085 37777 245113
rect 37811 245085 37839 245113
rect 37625 245023 37653 245051
rect 37687 245023 37715 245051
rect 37749 245023 37777 245051
rect 37811 245023 37839 245051
rect 37625 244961 37653 244989
rect 37687 244961 37715 244989
rect 37749 244961 37777 244989
rect 37811 244961 37839 244989
rect 37625 236147 37653 236175
rect 37687 236147 37715 236175
rect 37749 236147 37777 236175
rect 37811 236147 37839 236175
rect 37625 236085 37653 236113
rect 37687 236085 37715 236113
rect 37749 236085 37777 236113
rect 37811 236085 37839 236113
rect 37625 236023 37653 236051
rect 37687 236023 37715 236051
rect 37749 236023 37777 236051
rect 37811 236023 37839 236051
rect 37625 235961 37653 235989
rect 37687 235961 37715 235989
rect 37749 235961 37777 235989
rect 37811 235961 37839 235989
rect 37625 227147 37653 227175
rect 37687 227147 37715 227175
rect 37749 227147 37777 227175
rect 37811 227147 37839 227175
rect 37625 227085 37653 227113
rect 37687 227085 37715 227113
rect 37749 227085 37777 227113
rect 37811 227085 37839 227113
rect 37625 227023 37653 227051
rect 37687 227023 37715 227051
rect 37749 227023 37777 227051
rect 37811 227023 37839 227051
rect 37625 226961 37653 226989
rect 37687 226961 37715 226989
rect 37749 226961 37777 226989
rect 37811 226961 37839 226989
rect 37625 218147 37653 218175
rect 37687 218147 37715 218175
rect 37749 218147 37777 218175
rect 37811 218147 37839 218175
rect 37625 218085 37653 218113
rect 37687 218085 37715 218113
rect 37749 218085 37777 218113
rect 37811 218085 37839 218113
rect 37625 218023 37653 218051
rect 37687 218023 37715 218051
rect 37749 218023 37777 218051
rect 37811 218023 37839 218051
rect 37625 217961 37653 217989
rect 37687 217961 37715 217989
rect 37749 217961 37777 217989
rect 37811 217961 37839 217989
rect 37625 209147 37653 209175
rect 37687 209147 37715 209175
rect 37749 209147 37777 209175
rect 37811 209147 37839 209175
rect 37625 209085 37653 209113
rect 37687 209085 37715 209113
rect 37749 209085 37777 209113
rect 37811 209085 37839 209113
rect 37625 209023 37653 209051
rect 37687 209023 37715 209051
rect 37749 209023 37777 209051
rect 37811 209023 37839 209051
rect 37625 208961 37653 208989
rect 37687 208961 37715 208989
rect 37749 208961 37777 208989
rect 37811 208961 37839 208989
rect 37625 200147 37653 200175
rect 37687 200147 37715 200175
rect 37749 200147 37777 200175
rect 37811 200147 37839 200175
rect 37625 200085 37653 200113
rect 37687 200085 37715 200113
rect 37749 200085 37777 200113
rect 37811 200085 37839 200113
rect 37625 200023 37653 200051
rect 37687 200023 37715 200051
rect 37749 200023 37777 200051
rect 37811 200023 37839 200051
rect 37625 199961 37653 199989
rect 37687 199961 37715 199989
rect 37749 199961 37777 199989
rect 37811 199961 37839 199989
rect 37625 191147 37653 191175
rect 37687 191147 37715 191175
rect 37749 191147 37777 191175
rect 37811 191147 37839 191175
rect 37625 191085 37653 191113
rect 37687 191085 37715 191113
rect 37749 191085 37777 191113
rect 37811 191085 37839 191113
rect 37625 191023 37653 191051
rect 37687 191023 37715 191051
rect 37749 191023 37777 191051
rect 37811 191023 37839 191051
rect 37625 190961 37653 190989
rect 37687 190961 37715 190989
rect 37749 190961 37777 190989
rect 37811 190961 37839 190989
rect 37625 182147 37653 182175
rect 37687 182147 37715 182175
rect 37749 182147 37777 182175
rect 37811 182147 37839 182175
rect 37625 182085 37653 182113
rect 37687 182085 37715 182113
rect 37749 182085 37777 182113
rect 37811 182085 37839 182113
rect 37625 182023 37653 182051
rect 37687 182023 37715 182051
rect 37749 182023 37777 182051
rect 37811 182023 37839 182051
rect 37625 181961 37653 181989
rect 37687 181961 37715 181989
rect 37749 181961 37777 181989
rect 37811 181961 37839 181989
rect 37625 173147 37653 173175
rect 37687 173147 37715 173175
rect 37749 173147 37777 173175
rect 37811 173147 37839 173175
rect 37625 173085 37653 173113
rect 37687 173085 37715 173113
rect 37749 173085 37777 173113
rect 37811 173085 37839 173113
rect 37625 173023 37653 173051
rect 37687 173023 37715 173051
rect 37749 173023 37777 173051
rect 37811 173023 37839 173051
rect 37625 172961 37653 172989
rect 37687 172961 37715 172989
rect 37749 172961 37777 172989
rect 37811 172961 37839 172989
rect 37625 164147 37653 164175
rect 37687 164147 37715 164175
rect 37749 164147 37777 164175
rect 37811 164147 37839 164175
rect 37625 164085 37653 164113
rect 37687 164085 37715 164113
rect 37749 164085 37777 164113
rect 37811 164085 37839 164113
rect 37625 164023 37653 164051
rect 37687 164023 37715 164051
rect 37749 164023 37777 164051
rect 37811 164023 37839 164051
rect 37625 163961 37653 163989
rect 37687 163961 37715 163989
rect 37749 163961 37777 163989
rect 37811 163961 37839 163989
rect 37625 155147 37653 155175
rect 37687 155147 37715 155175
rect 37749 155147 37777 155175
rect 37811 155147 37839 155175
rect 37625 155085 37653 155113
rect 37687 155085 37715 155113
rect 37749 155085 37777 155113
rect 37811 155085 37839 155113
rect 37625 155023 37653 155051
rect 37687 155023 37715 155051
rect 37749 155023 37777 155051
rect 37811 155023 37839 155051
rect 37625 154961 37653 154989
rect 37687 154961 37715 154989
rect 37749 154961 37777 154989
rect 37811 154961 37839 154989
rect 37625 146147 37653 146175
rect 37687 146147 37715 146175
rect 37749 146147 37777 146175
rect 37811 146147 37839 146175
rect 37625 146085 37653 146113
rect 37687 146085 37715 146113
rect 37749 146085 37777 146113
rect 37811 146085 37839 146113
rect 37625 146023 37653 146051
rect 37687 146023 37715 146051
rect 37749 146023 37777 146051
rect 37811 146023 37839 146051
rect 37625 145961 37653 145989
rect 37687 145961 37715 145989
rect 37749 145961 37777 145989
rect 37811 145961 37839 145989
rect 37625 137147 37653 137175
rect 37687 137147 37715 137175
rect 37749 137147 37777 137175
rect 37811 137147 37839 137175
rect 37625 137085 37653 137113
rect 37687 137085 37715 137113
rect 37749 137085 37777 137113
rect 37811 137085 37839 137113
rect 37625 137023 37653 137051
rect 37687 137023 37715 137051
rect 37749 137023 37777 137051
rect 37811 137023 37839 137051
rect 37625 136961 37653 136989
rect 37687 136961 37715 136989
rect 37749 136961 37777 136989
rect 37811 136961 37839 136989
rect 37625 128147 37653 128175
rect 37687 128147 37715 128175
rect 37749 128147 37777 128175
rect 37811 128147 37839 128175
rect 37625 128085 37653 128113
rect 37687 128085 37715 128113
rect 37749 128085 37777 128113
rect 37811 128085 37839 128113
rect 37625 128023 37653 128051
rect 37687 128023 37715 128051
rect 37749 128023 37777 128051
rect 37811 128023 37839 128051
rect 37625 127961 37653 127989
rect 37687 127961 37715 127989
rect 37749 127961 37777 127989
rect 37811 127961 37839 127989
rect 37625 119147 37653 119175
rect 37687 119147 37715 119175
rect 37749 119147 37777 119175
rect 37811 119147 37839 119175
rect 37625 119085 37653 119113
rect 37687 119085 37715 119113
rect 37749 119085 37777 119113
rect 37811 119085 37839 119113
rect 37625 119023 37653 119051
rect 37687 119023 37715 119051
rect 37749 119023 37777 119051
rect 37811 119023 37839 119051
rect 37625 118961 37653 118989
rect 37687 118961 37715 118989
rect 37749 118961 37777 118989
rect 37811 118961 37839 118989
rect 37625 110147 37653 110175
rect 37687 110147 37715 110175
rect 37749 110147 37777 110175
rect 37811 110147 37839 110175
rect 37625 110085 37653 110113
rect 37687 110085 37715 110113
rect 37749 110085 37777 110113
rect 37811 110085 37839 110113
rect 37625 110023 37653 110051
rect 37687 110023 37715 110051
rect 37749 110023 37777 110051
rect 37811 110023 37839 110051
rect 37625 109961 37653 109989
rect 37687 109961 37715 109989
rect 37749 109961 37777 109989
rect 37811 109961 37839 109989
rect 37625 101147 37653 101175
rect 37687 101147 37715 101175
rect 37749 101147 37777 101175
rect 37811 101147 37839 101175
rect 37625 101085 37653 101113
rect 37687 101085 37715 101113
rect 37749 101085 37777 101113
rect 37811 101085 37839 101113
rect 37625 101023 37653 101051
rect 37687 101023 37715 101051
rect 37749 101023 37777 101051
rect 37811 101023 37839 101051
rect 37625 100961 37653 100989
rect 37687 100961 37715 100989
rect 37749 100961 37777 100989
rect 37811 100961 37839 100989
rect 37625 92147 37653 92175
rect 37687 92147 37715 92175
rect 37749 92147 37777 92175
rect 37811 92147 37839 92175
rect 37625 92085 37653 92113
rect 37687 92085 37715 92113
rect 37749 92085 37777 92113
rect 37811 92085 37839 92113
rect 37625 92023 37653 92051
rect 37687 92023 37715 92051
rect 37749 92023 37777 92051
rect 37811 92023 37839 92051
rect 37625 91961 37653 91989
rect 37687 91961 37715 91989
rect 37749 91961 37777 91989
rect 37811 91961 37839 91989
rect 37625 83147 37653 83175
rect 37687 83147 37715 83175
rect 37749 83147 37777 83175
rect 37811 83147 37839 83175
rect 37625 83085 37653 83113
rect 37687 83085 37715 83113
rect 37749 83085 37777 83113
rect 37811 83085 37839 83113
rect 37625 83023 37653 83051
rect 37687 83023 37715 83051
rect 37749 83023 37777 83051
rect 37811 83023 37839 83051
rect 37625 82961 37653 82989
rect 37687 82961 37715 82989
rect 37749 82961 37777 82989
rect 37811 82961 37839 82989
rect 37625 74147 37653 74175
rect 37687 74147 37715 74175
rect 37749 74147 37777 74175
rect 37811 74147 37839 74175
rect 37625 74085 37653 74113
rect 37687 74085 37715 74113
rect 37749 74085 37777 74113
rect 37811 74085 37839 74113
rect 37625 74023 37653 74051
rect 37687 74023 37715 74051
rect 37749 74023 37777 74051
rect 37811 74023 37839 74051
rect 37625 73961 37653 73989
rect 37687 73961 37715 73989
rect 37749 73961 37777 73989
rect 37811 73961 37839 73989
rect 37625 65147 37653 65175
rect 37687 65147 37715 65175
rect 37749 65147 37777 65175
rect 37811 65147 37839 65175
rect 37625 65085 37653 65113
rect 37687 65085 37715 65113
rect 37749 65085 37777 65113
rect 37811 65085 37839 65113
rect 37625 65023 37653 65051
rect 37687 65023 37715 65051
rect 37749 65023 37777 65051
rect 37811 65023 37839 65051
rect 37625 64961 37653 64989
rect 37687 64961 37715 64989
rect 37749 64961 37777 64989
rect 37811 64961 37839 64989
rect 37625 56147 37653 56175
rect 37687 56147 37715 56175
rect 37749 56147 37777 56175
rect 37811 56147 37839 56175
rect 37625 56085 37653 56113
rect 37687 56085 37715 56113
rect 37749 56085 37777 56113
rect 37811 56085 37839 56113
rect 37625 56023 37653 56051
rect 37687 56023 37715 56051
rect 37749 56023 37777 56051
rect 37811 56023 37839 56051
rect 37625 55961 37653 55989
rect 37687 55961 37715 55989
rect 37749 55961 37777 55989
rect 37811 55961 37839 55989
rect 37625 47147 37653 47175
rect 37687 47147 37715 47175
rect 37749 47147 37777 47175
rect 37811 47147 37839 47175
rect 37625 47085 37653 47113
rect 37687 47085 37715 47113
rect 37749 47085 37777 47113
rect 37811 47085 37839 47113
rect 37625 47023 37653 47051
rect 37687 47023 37715 47051
rect 37749 47023 37777 47051
rect 37811 47023 37839 47051
rect 37625 46961 37653 46989
rect 37687 46961 37715 46989
rect 37749 46961 37777 46989
rect 37811 46961 37839 46989
rect 37625 38147 37653 38175
rect 37687 38147 37715 38175
rect 37749 38147 37777 38175
rect 37811 38147 37839 38175
rect 37625 38085 37653 38113
rect 37687 38085 37715 38113
rect 37749 38085 37777 38113
rect 37811 38085 37839 38113
rect 37625 38023 37653 38051
rect 37687 38023 37715 38051
rect 37749 38023 37777 38051
rect 37811 38023 37839 38051
rect 37625 37961 37653 37989
rect 37687 37961 37715 37989
rect 37749 37961 37777 37989
rect 37811 37961 37839 37989
rect 37625 29147 37653 29175
rect 37687 29147 37715 29175
rect 37749 29147 37777 29175
rect 37811 29147 37839 29175
rect 37625 29085 37653 29113
rect 37687 29085 37715 29113
rect 37749 29085 37777 29113
rect 37811 29085 37839 29113
rect 37625 29023 37653 29051
rect 37687 29023 37715 29051
rect 37749 29023 37777 29051
rect 37811 29023 37839 29051
rect 37625 28961 37653 28989
rect 37687 28961 37715 28989
rect 37749 28961 37777 28989
rect 37811 28961 37839 28989
rect 37625 20147 37653 20175
rect 37687 20147 37715 20175
rect 37749 20147 37777 20175
rect 37811 20147 37839 20175
rect 37625 20085 37653 20113
rect 37687 20085 37715 20113
rect 37749 20085 37777 20113
rect 37811 20085 37839 20113
rect 37625 20023 37653 20051
rect 37687 20023 37715 20051
rect 37749 20023 37777 20051
rect 37811 20023 37839 20051
rect 37625 19961 37653 19989
rect 37687 19961 37715 19989
rect 37749 19961 37777 19989
rect 37811 19961 37839 19989
rect 37625 11147 37653 11175
rect 37687 11147 37715 11175
rect 37749 11147 37777 11175
rect 37811 11147 37839 11175
rect 37625 11085 37653 11113
rect 37687 11085 37715 11113
rect 37749 11085 37777 11113
rect 37811 11085 37839 11113
rect 37625 11023 37653 11051
rect 37687 11023 37715 11051
rect 37749 11023 37777 11051
rect 37811 11023 37839 11051
rect 37625 10961 37653 10989
rect 37687 10961 37715 10989
rect 37749 10961 37777 10989
rect 37811 10961 37839 10989
rect 37625 2147 37653 2175
rect 37687 2147 37715 2175
rect 37749 2147 37777 2175
rect 37811 2147 37839 2175
rect 37625 2085 37653 2113
rect 37687 2085 37715 2113
rect 37749 2085 37777 2113
rect 37811 2085 37839 2113
rect 37625 2023 37653 2051
rect 37687 2023 37715 2051
rect 37749 2023 37777 2051
rect 37811 2023 37839 2051
rect 37625 1961 37653 1989
rect 37687 1961 37715 1989
rect 37749 1961 37777 1989
rect 37811 1961 37839 1989
rect 37625 -108 37653 -80
rect 37687 -108 37715 -80
rect 37749 -108 37777 -80
rect 37811 -108 37839 -80
rect 37625 -170 37653 -142
rect 37687 -170 37715 -142
rect 37749 -170 37777 -142
rect 37811 -170 37839 -142
rect 37625 -232 37653 -204
rect 37687 -232 37715 -204
rect 37749 -232 37777 -204
rect 37811 -232 37839 -204
rect 37625 -294 37653 -266
rect 37687 -294 37715 -266
rect 37749 -294 37777 -266
rect 37811 -294 37839 -266
rect 39485 299058 39513 299086
rect 39547 299058 39575 299086
rect 39609 299058 39637 299086
rect 39671 299058 39699 299086
rect 39485 298996 39513 299024
rect 39547 298996 39575 299024
rect 39609 298996 39637 299024
rect 39671 298996 39699 299024
rect 39485 298934 39513 298962
rect 39547 298934 39575 298962
rect 39609 298934 39637 298962
rect 39671 298934 39699 298962
rect 39485 298872 39513 298900
rect 39547 298872 39575 298900
rect 39609 298872 39637 298900
rect 39671 298872 39699 298900
rect 39485 293147 39513 293175
rect 39547 293147 39575 293175
rect 39609 293147 39637 293175
rect 39671 293147 39699 293175
rect 39485 293085 39513 293113
rect 39547 293085 39575 293113
rect 39609 293085 39637 293113
rect 39671 293085 39699 293113
rect 39485 293023 39513 293051
rect 39547 293023 39575 293051
rect 39609 293023 39637 293051
rect 39671 293023 39699 293051
rect 39485 292961 39513 292989
rect 39547 292961 39575 292989
rect 39609 292961 39637 292989
rect 39671 292961 39699 292989
rect 39485 284147 39513 284175
rect 39547 284147 39575 284175
rect 39609 284147 39637 284175
rect 39671 284147 39699 284175
rect 39485 284085 39513 284113
rect 39547 284085 39575 284113
rect 39609 284085 39637 284113
rect 39671 284085 39699 284113
rect 39485 284023 39513 284051
rect 39547 284023 39575 284051
rect 39609 284023 39637 284051
rect 39671 284023 39699 284051
rect 39485 283961 39513 283989
rect 39547 283961 39575 283989
rect 39609 283961 39637 283989
rect 39671 283961 39699 283989
rect 39485 275147 39513 275175
rect 39547 275147 39575 275175
rect 39609 275147 39637 275175
rect 39671 275147 39699 275175
rect 39485 275085 39513 275113
rect 39547 275085 39575 275113
rect 39609 275085 39637 275113
rect 39671 275085 39699 275113
rect 39485 275023 39513 275051
rect 39547 275023 39575 275051
rect 39609 275023 39637 275051
rect 39671 275023 39699 275051
rect 39485 274961 39513 274989
rect 39547 274961 39575 274989
rect 39609 274961 39637 274989
rect 39671 274961 39699 274989
rect 39485 266147 39513 266175
rect 39547 266147 39575 266175
rect 39609 266147 39637 266175
rect 39671 266147 39699 266175
rect 39485 266085 39513 266113
rect 39547 266085 39575 266113
rect 39609 266085 39637 266113
rect 39671 266085 39699 266113
rect 39485 266023 39513 266051
rect 39547 266023 39575 266051
rect 39609 266023 39637 266051
rect 39671 266023 39699 266051
rect 39485 265961 39513 265989
rect 39547 265961 39575 265989
rect 39609 265961 39637 265989
rect 39671 265961 39699 265989
rect 39485 257147 39513 257175
rect 39547 257147 39575 257175
rect 39609 257147 39637 257175
rect 39671 257147 39699 257175
rect 39485 257085 39513 257113
rect 39547 257085 39575 257113
rect 39609 257085 39637 257113
rect 39671 257085 39699 257113
rect 39485 257023 39513 257051
rect 39547 257023 39575 257051
rect 39609 257023 39637 257051
rect 39671 257023 39699 257051
rect 39485 256961 39513 256989
rect 39547 256961 39575 256989
rect 39609 256961 39637 256989
rect 39671 256961 39699 256989
rect 39485 248147 39513 248175
rect 39547 248147 39575 248175
rect 39609 248147 39637 248175
rect 39671 248147 39699 248175
rect 39485 248085 39513 248113
rect 39547 248085 39575 248113
rect 39609 248085 39637 248113
rect 39671 248085 39699 248113
rect 39485 248023 39513 248051
rect 39547 248023 39575 248051
rect 39609 248023 39637 248051
rect 39671 248023 39699 248051
rect 39485 247961 39513 247989
rect 39547 247961 39575 247989
rect 39609 247961 39637 247989
rect 39671 247961 39699 247989
rect 39485 239147 39513 239175
rect 39547 239147 39575 239175
rect 39609 239147 39637 239175
rect 39671 239147 39699 239175
rect 39485 239085 39513 239113
rect 39547 239085 39575 239113
rect 39609 239085 39637 239113
rect 39671 239085 39699 239113
rect 39485 239023 39513 239051
rect 39547 239023 39575 239051
rect 39609 239023 39637 239051
rect 39671 239023 39699 239051
rect 39485 238961 39513 238989
rect 39547 238961 39575 238989
rect 39609 238961 39637 238989
rect 39671 238961 39699 238989
rect 39485 230147 39513 230175
rect 39547 230147 39575 230175
rect 39609 230147 39637 230175
rect 39671 230147 39699 230175
rect 39485 230085 39513 230113
rect 39547 230085 39575 230113
rect 39609 230085 39637 230113
rect 39671 230085 39699 230113
rect 39485 230023 39513 230051
rect 39547 230023 39575 230051
rect 39609 230023 39637 230051
rect 39671 230023 39699 230051
rect 39485 229961 39513 229989
rect 39547 229961 39575 229989
rect 39609 229961 39637 229989
rect 39671 229961 39699 229989
rect 39485 221147 39513 221175
rect 39547 221147 39575 221175
rect 39609 221147 39637 221175
rect 39671 221147 39699 221175
rect 39485 221085 39513 221113
rect 39547 221085 39575 221113
rect 39609 221085 39637 221113
rect 39671 221085 39699 221113
rect 39485 221023 39513 221051
rect 39547 221023 39575 221051
rect 39609 221023 39637 221051
rect 39671 221023 39699 221051
rect 39485 220961 39513 220989
rect 39547 220961 39575 220989
rect 39609 220961 39637 220989
rect 39671 220961 39699 220989
rect 39485 212147 39513 212175
rect 39547 212147 39575 212175
rect 39609 212147 39637 212175
rect 39671 212147 39699 212175
rect 39485 212085 39513 212113
rect 39547 212085 39575 212113
rect 39609 212085 39637 212113
rect 39671 212085 39699 212113
rect 39485 212023 39513 212051
rect 39547 212023 39575 212051
rect 39609 212023 39637 212051
rect 39671 212023 39699 212051
rect 39485 211961 39513 211989
rect 39547 211961 39575 211989
rect 39609 211961 39637 211989
rect 39671 211961 39699 211989
rect 39485 203147 39513 203175
rect 39547 203147 39575 203175
rect 39609 203147 39637 203175
rect 39671 203147 39699 203175
rect 39485 203085 39513 203113
rect 39547 203085 39575 203113
rect 39609 203085 39637 203113
rect 39671 203085 39699 203113
rect 39485 203023 39513 203051
rect 39547 203023 39575 203051
rect 39609 203023 39637 203051
rect 39671 203023 39699 203051
rect 39485 202961 39513 202989
rect 39547 202961 39575 202989
rect 39609 202961 39637 202989
rect 39671 202961 39699 202989
rect 39485 194147 39513 194175
rect 39547 194147 39575 194175
rect 39609 194147 39637 194175
rect 39671 194147 39699 194175
rect 39485 194085 39513 194113
rect 39547 194085 39575 194113
rect 39609 194085 39637 194113
rect 39671 194085 39699 194113
rect 39485 194023 39513 194051
rect 39547 194023 39575 194051
rect 39609 194023 39637 194051
rect 39671 194023 39699 194051
rect 39485 193961 39513 193989
rect 39547 193961 39575 193989
rect 39609 193961 39637 193989
rect 39671 193961 39699 193989
rect 39485 185147 39513 185175
rect 39547 185147 39575 185175
rect 39609 185147 39637 185175
rect 39671 185147 39699 185175
rect 39485 185085 39513 185113
rect 39547 185085 39575 185113
rect 39609 185085 39637 185113
rect 39671 185085 39699 185113
rect 39485 185023 39513 185051
rect 39547 185023 39575 185051
rect 39609 185023 39637 185051
rect 39671 185023 39699 185051
rect 39485 184961 39513 184989
rect 39547 184961 39575 184989
rect 39609 184961 39637 184989
rect 39671 184961 39699 184989
rect 39485 176147 39513 176175
rect 39547 176147 39575 176175
rect 39609 176147 39637 176175
rect 39671 176147 39699 176175
rect 39485 176085 39513 176113
rect 39547 176085 39575 176113
rect 39609 176085 39637 176113
rect 39671 176085 39699 176113
rect 39485 176023 39513 176051
rect 39547 176023 39575 176051
rect 39609 176023 39637 176051
rect 39671 176023 39699 176051
rect 39485 175961 39513 175989
rect 39547 175961 39575 175989
rect 39609 175961 39637 175989
rect 39671 175961 39699 175989
rect 39485 167147 39513 167175
rect 39547 167147 39575 167175
rect 39609 167147 39637 167175
rect 39671 167147 39699 167175
rect 39485 167085 39513 167113
rect 39547 167085 39575 167113
rect 39609 167085 39637 167113
rect 39671 167085 39699 167113
rect 39485 167023 39513 167051
rect 39547 167023 39575 167051
rect 39609 167023 39637 167051
rect 39671 167023 39699 167051
rect 39485 166961 39513 166989
rect 39547 166961 39575 166989
rect 39609 166961 39637 166989
rect 39671 166961 39699 166989
rect 39485 158147 39513 158175
rect 39547 158147 39575 158175
rect 39609 158147 39637 158175
rect 39671 158147 39699 158175
rect 39485 158085 39513 158113
rect 39547 158085 39575 158113
rect 39609 158085 39637 158113
rect 39671 158085 39699 158113
rect 39485 158023 39513 158051
rect 39547 158023 39575 158051
rect 39609 158023 39637 158051
rect 39671 158023 39699 158051
rect 39485 157961 39513 157989
rect 39547 157961 39575 157989
rect 39609 157961 39637 157989
rect 39671 157961 39699 157989
rect 39485 149147 39513 149175
rect 39547 149147 39575 149175
rect 39609 149147 39637 149175
rect 39671 149147 39699 149175
rect 39485 149085 39513 149113
rect 39547 149085 39575 149113
rect 39609 149085 39637 149113
rect 39671 149085 39699 149113
rect 39485 149023 39513 149051
rect 39547 149023 39575 149051
rect 39609 149023 39637 149051
rect 39671 149023 39699 149051
rect 39485 148961 39513 148989
rect 39547 148961 39575 148989
rect 39609 148961 39637 148989
rect 39671 148961 39699 148989
rect 39485 140147 39513 140175
rect 39547 140147 39575 140175
rect 39609 140147 39637 140175
rect 39671 140147 39699 140175
rect 39485 140085 39513 140113
rect 39547 140085 39575 140113
rect 39609 140085 39637 140113
rect 39671 140085 39699 140113
rect 39485 140023 39513 140051
rect 39547 140023 39575 140051
rect 39609 140023 39637 140051
rect 39671 140023 39699 140051
rect 39485 139961 39513 139989
rect 39547 139961 39575 139989
rect 39609 139961 39637 139989
rect 39671 139961 39699 139989
rect 39485 131147 39513 131175
rect 39547 131147 39575 131175
rect 39609 131147 39637 131175
rect 39671 131147 39699 131175
rect 39485 131085 39513 131113
rect 39547 131085 39575 131113
rect 39609 131085 39637 131113
rect 39671 131085 39699 131113
rect 39485 131023 39513 131051
rect 39547 131023 39575 131051
rect 39609 131023 39637 131051
rect 39671 131023 39699 131051
rect 39485 130961 39513 130989
rect 39547 130961 39575 130989
rect 39609 130961 39637 130989
rect 39671 130961 39699 130989
rect 39485 122147 39513 122175
rect 39547 122147 39575 122175
rect 39609 122147 39637 122175
rect 39671 122147 39699 122175
rect 39485 122085 39513 122113
rect 39547 122085 39575 122113
rect 39609 122085 39637 122113
rect 39671 122085 39699 122113
rect 39485 122023 39513 122051
rect 39547 122023 39575 122051
rect 39609 122023 39637 122051
rect 39671 122023 39699 122051
rect 39485 121961 39513 121989
rect 39547 121961 39575 121989
rect 39609 121961 39637 121989
rect 39671 121961 39699 121989
rect 39485 113147 39513 113175
rect 39547 113147 39575 113175
rect 39609 113147 39637 113175
rect 39671 113147 39699 113175
rect 39485 113085 39513 113113
rect 39547 113085 39575 113113
rect 39609 113085 39637 113113
rect 39671 113085 39699 113113
rect 39485 113023 39513 113051
rect 39547 113023 39575 113051
rect 39609 113023 39637 113051
rect 39671 113023 39699 113051
rect 39485 112961 39513 112989
rect 39547 112961 39575 112989
rect 39609 112961 39637 112989
rect 39671 112961 39699 112989
rect 39485 104147 39513 104175
rect 39547 104147 39575 104175
rect 39609 104147 39637 104175
rect 39671 104147 39699 104175
rect 39485 104085 39513 104113
rect 39547 104085 39575 104113
rect 39609 104085 39637 104113
rect 39671 104085 39699 104113
rect 39485 104023 39513 104051
rect 39547 104023 39575 104051
rect 39609 104023 39637 104051
rect 39671 104023 39699 104051
rect 39485 103961 39513 103989
rect 39547 103961 39575 103989
rect 39609 103961 39637 103989
rect 39671 103961 39699 103989
rect 39485 95147 39513 95175
rect 39547 95147 39575 95175
rect 39609 95147 39637 95175
rect 39671 95147 39699 95175
rect 39485 95085 39513 95113
rect 39547 95085 39575 95113
rect 39609 95085 39637 95113
rect 39671 95085 39699 95113
rect 39485 95023 39513 95051
rect 39547 95023 39575 95051
rect 39609 95023 39637 95051
rect 39671 95023 39699 95051
rect 39485 94961 39513 94989
rect 39547 94961 39575 94989
rect 39609 94961 39637 94989
rect 39671 94961 39699 94989
rect 39485 86147 39513 86175
rect 39547 86147 39575 86175
rect 39609 86147 39637 86175
rect 39671 86147 39699 86175
rect 39485 86085 39513 86113
rect 39547 86085 39575 86113
rect 39609 86085 39637 86113
rect 39671 86085 39699 86113
rect 39485 86023 39513 86051
rect 39547 86023 39575 86051
rect 39609 86023 39637 86051
rect 39671 86023 39699 86051
rect 39485 85961 39513 85989
rect 39547 85961 39575 85989
rect 39609 85961 39637 85989
rect 39671 85961 39699 85989
rect 39485 77147 39513 77175
rect 39547 77147 39575 77175
rect 39609 77147 39637 77175
rect 39671 77147 39699 77175
rect 39485 77085 39513 77113
rect 39547 77085 39575 77113
rect 39609 77085 39637 77113
rect 39671 77085 39699 77113
rect 39485 77023 39513 77051
rect 39547 77023 39575 77051
rect 39609 77023 39637 77051
rect 39671 77023 39699 77051
rect 39485 76961 39513 76989
rect 39547 76961 39575 76989
rect 39609 76961 39637 76989
rect 39671 76961 39699 76989
rect 39485 68147 39513 68175
rect 39547 68147 39575 68175
rect 39609 68147 39637 68175
rect 39671 68147 39699 68175
rect 39485 68085 39513 68113
rect 39547 68085 39575 68113
rect 39609 68085 39637 68113
rect 39671 68085 39699 68113
rect 39485 68023 39513 68051
rect 39547 68023 39575 68051
rect 39609 68023 39637 68051
rect 39671 68023 39699 68051
rect 39485 67961 39513 67989
rect 39547 67961 39575 67989
rect 39609 67961 39637 67989
rect 39671 67961 39699 67989
rect 39485 59147 39513 59175
rect 39547 59147 39575 59175
rect 39609 59147 39637 59175
rect 39671 59147 39699 59175
rect 39485 59085 39513 59113
rect 39547 59085 39575 59113
rect 39609 59085 39637 59113
rect 39671 59085 39699 59113
rect 39485 59023 39513 59051
rect 39547 59023 39575 59051
rect 39609 59023 39637 59051
rect 39671 59023 39699 59051
rect 39485 58961 39513 58989
rect 39547 58961 39575 58989
rect 39609 58961 39637 58989
rect 39671 58961 39699 58989
rect 39485 50147 39513 50175
rect 39547 50147 39575 50175
rect 39609 50147 39637 50175
rect 39671 50147 39699 50175
rect 39485 50085 39513 50113
rect 39547 50085 39575 50113
rect 39609 50085 39637 50113
rect 39671 50085 39699 50113
rect 39485 50023 39513 50051
rect 39547 50023 39575 50051
rect 39609 50023 39637 50051
rect 39671 50023 39699 50051
rect 39485 49961 39513 49989
rect 39547 49961 39575 49989
rect 39609 49961 39637 49989
rect 39671 49961 39699 49989
rect 39485 41147 39513 41175
rect 39547 41147 39575 41175
rect 39609 41147 39637 41175
rect 39671 41147 39699 41175
rect 39485 41085 39513 41113
rect 39547 41085 39575 41113
rect 39609 41085 39637 41113
rect 39671 41085 39699 41113
rect 39485 41023 39513 41051
rect 39547 41023 39575 41051
rect 39609 41023 39637 41051
rect 39671 41023 39699 41051
rect 39485 40961 39513 40989
rect 39547 40961 39575 40989
rect 39609 40961 39637 40989
rect 39671 40961 39699 40989
rect 39485 32147 39513 32175
rect 39547 32147 39575 32175
rect 39609 32147 39637 32175
rect 39671 32147 39699 32175
rect 39485 32085 39513 32113
rect 39547 32085 39575 32113
rect 39609 32085 39637 32113
rect 39671 32085 39699 32113
rect 39485 32023 39513 32051
rect 39547 32023 39575 32051
rect 39609 32023 39637 32051
rect 39671 32023 39699 32051
rect 39485 31961 39513 31989
rect 39547 31961 39575 31989
rect 39609 31961 39637 31989
rect 39671 31961 39699 31989
rect 39485 23147 39513 23175
rect 39547 23147 39575 23175
rect 39609 23147 39637 23175
rect 39671 23147 39699 23175
rect 39485 23085 39513 23113
rect 39547 23085 39575 23113
rect 39609 23085 39637 23113
rect 39671 23085 39699 23113
rect 39485 23023 39513 23051
rect 39547 23023 39575 23051
rect 39609 23023 39637 23051
rect 39671 23023 39699 23051
rect 39485 22961 39513 22989
rect 39547 22961 39575 22989
rect 39609 22961 39637 22989
rect 39671 22961 39699 22989
rect 39485 14147 39513 14175
rect 39547 14147 39575 14175
rect 39609 14147 39637 14175
rect 39671 14147 39699 14175
rect 39485 14085 39513 14113
rect 39547 14085 39575 14113
rect 39609 14085 39637 14113
rect 39671 14085 39699 14113
rect 39485 14023 39513 14051
rect 39547 14023 39575 14051
rect 39609 14023 39637 14051
rect 39671 14023 39699 14051
rect 39485 13961 39513 13989
rect 39547 13961 39575 13989
rect 39609 13961 39637 13989
rect 39671 13961 39699 13989
rect 39485 5147 39513 5175
rect 39547 5147 39575 5175
rect 39609 5147 39637 5175
rect 39671 5147 39699 5175
rect 39485 5085 39513 5113
rect 39547 5085 39575 5113
rect 39609 5085 39637 5113
rect 39671 5085 39699 5113
rect 39485 5023 39513 5051
rect 39547 5023 39575 5051
rect 39609 5023 39637 5051
rect 39671 5023 39699 5051
rect 39485 4961 39513 4989
rect 39547 4961 39575 4989
rect 39609 4961 39637 4989
rect 39671 4961 39699 4989
rect 39485 -588 39513 -560
rect 39547 -588 39575 -560
rect 39609 -588 39637 -560
rect 39671 -588 39699 -560
rect 39485 -650 39513 -622
rect 39547 -650 39575 -622
rect 39609 -650 39637 -622
rect 39671 -650 39699 -622
rect 39485 -712 39513 -684
rect 39547 -712 39575 -684
rect 39609 -712 39637 -684
rect 39671 -712 39699 -684
rect 39485 -774 39513 -746
rect 39547 -774 39575 -746
rect 39609 -774 39637 -746
rect 39671 -774 39699 -746
rect 46625 298578 46653 298606
rect 46687 298578 46715 298606
rect 46749 298578 46777 298606
rect 46811 298578 46839 298606
rect 46625 298516 46653 298544
rect 46687 298516 46715 298544
rect 46749 298516 46777 298544
rect 46811 298516 46839 298544
rect 46625 298454 46653 298482
rect 46687 298454 46715 298482
rect 46749 298454 46777 298482
rect 46811 298454 46839 298482
rect 46625 298392 46653 298420
rect 46687 298392 46715 298420
rect 46749 298392 46777 298420
rect 46811 298392 46839 298420
rect 46625 290147 46653 290175
rect 46687 290147 46715 290175
rect 46749 290147 46777 290175
rect 46811 290147 46839 290175
rect 46625 290085 46653 290113
rect 46687 290085 46715 290113
rect 46749 290085 46777 290113
rect 46811 290085 46839 290113
rect 46625 290023 46653 290051
rect 46687 290023 46715 290051
rect 46749 290023 46777 290051
rect 46811 290023 46839 290051
rect 46625 289961 46653 289989
rect 46687 289961 46715 289989
rect 46749 289961 46777 289989
rect 46811 289961 46839 289989
rect 46625 281147 46653 281175
rect 46687 281147 46715 281175
rect 46749 281147 46777 281175
rect 46811 281147 46839 281175
rect 46625 281085 46653 281113
rect 46687 281085 46715 281113
rect 46749 281085 46777 281113
rect 46811 281085 46839 281113
rect 46625 281023 46653 281051
rect 46687 281023 46715 281051
rect 46749 281023 46777 281051
rect 46811 281023 46839 281051
rect 46625 280961 46653 280989
rect 46687 280961 46715 280989
rect 46749 280961 46777 280989
rect 46811 280961 46839 280989
rect 46625 272147 46653 272175
rect 46687 272147 46715 272175
rect 46749 272147 46777 272175
rect 46811 272147 46839 272175
rect 46625 272085 46653 272113
rect 46687 272085 46715 272113
rect 46749 272085 46777 272113
rect 46811 272085 46839 272113
rect 46625 272023 46653 272051
rect 46687 272023 46715 272051
rect 46749 272023 46777 272051
rect 46811 272023 46839 272051
rect 46625 271961 46653 271989
rect 46687 271961 46715 271989
rect 46749 271961 46777 271989
rect 46811 271961 46839 271989
rect 46625 263147 46653 263175
rect 46687 263147 46715 263175
rect 46749 263147 46777 263175
rect 46811 263147 46839 263175
rect 46625 263085 46653 263113
rect 46687 263085 46715 263113
rect 46749 263085 46777 263113
rect 46811 263085 46839 263113
rect 46625 263023 46653 263051
rect 46687 263023 46715 263051
rect 46749 263023 46777 263051
rect 46811 263023 46839 263051
rect 46625 262961 46653 262989
rect 46687 262961 46715 262989
rect 46749 262961 46777 262989
rect 46811 262961 46839 262989
rect 46625 254147 46653 254175
rect 46687 254147 46715 254175
rect 46749 254147 46777 254175
rect 46811 254147 46839 254175
rect 46625 254085 46653 254113
rect 46687 254085 46715 254113
rect 46749 254085 46777 254113
rect 46811 254085 46839 254113
rect 46625 254023 46653 254051
rect 46687 254023 46715 254051
rect 46749 254023 46777 254051
rect 46811 254023 46839 254051
rect 46625 253961 46653 253989
rect 46687 253961 46715 253989
rect 46749 253961 46777 253989
rect 46811 253961 46839 253989
rect 46625 245147 46653 245175
rect 46687 245147 46715 245175
rect 46749 245147 46777 245175
rect 46811 245147 46839 245175
rect 46625 245085 46653 245113
rect 46687 245085 46715 245113
rect 46749 245085 46777 245113
rect 46811 245085 46839 245113
rect 46625 245023 46653 245051
rect 46687 245023 46715 245051
rect 46749 245023 46777 245051
rect 46811 245023 46839 245051
rect 46625 244961 46653 244989
rect 46687 244961 46715 244989
rect 46749 244961 46777 244989
rect 46811 244961 46839 244989
rect 46625 236147 46653 236175
rect 46687 236147 46715 236175
rect 46749 236147 46777 236175
rect 46811 236147 46839 236175
rect 46625 236085 46653 236113
rect 46687 236085 46715 236113
rect 46749 236085 46777 236113
rect 46811 236085 46839 236113
rect 46625 236023 46653 236051
rect 46687 236023 46715 236051
rect 46749 236023 46777 236051
rect 46811 236023 46839 236051
rect 46625 235961 46653 235989
rect 46687 235961 46715 235989
rect 46749 235961 46777 235989
rect 46811 235961 46839 235989
rect 46625 227147 46653 227175
rect 46687 227147 46715 227175
rect 46749 227147 46777 227175
rect 46811 227147 46839 227175
rect 46625 227085 46653 227113
rect 46687 227085 46715 227113
rect 46749 227085 46777 227113
rect 46811 227085 46839 227113
rect 46625 227023 46653 227051
rect 46687 227023 46715 227051
rect 46749 227023 46777 227051
rect 46811 227023 46839 227051
rect 46625 226961 46653 226989
rect 46687 226961 46715 226989
rect 46749 226961 46777 226989
rect 46811 226961 46839 226989
rect 46625 218147 46653 218175
rect 46687 218147 46715 218175
rect 46749 218147 46777 218175
rect 46811 218147 46839 218175
rect 46625 218085 46653 218113
rect 46687 218085 46715 218113
rect 46749 218085 46777 218113
rect 46811 218085 46839 218113
rect 46625 218023 46653 218051
rect 46687 218023 46715 218051
rect 46749 218023 46777 218051
rect 46811 218023 46839 218051
rect 46625 217961 46653 217989
rect 46687 217961 46715 217989
rect 46749 217961 46777 217989
rect 46811 217961 46839 217989
rect 46625 209147 46653 209175
rect 46687 209147 46715 209175
rect 46749 209147 46777 209175
rect 46811 209147 46839 209175
rect 46625 209085 46653 209113
rect 46687 209085 46715 209113
rect 46749 209085 46777 209113
rect 46811 209085 46839 209113
rect 46625 209023 46653 209051
rect 46687 209023 46715 209051
rect 46749 209023 46777 209051
rect 46811 209023 46839 209051
rect 46625 208961 46653 208989
rect 46687 208961 46715 208989
rect 46749 208961 46777 208989
rect 46811 208961 46839 208989
rect 46625 200147 46653 200175
rect 46687 200147 46715 200175
rect 46749 200147 46777 200175
rect 46811 200147 46839 200175
rect 46625 200085 46653 200113
rect 46687 200085 46715 200113
rect 46749 200085 46777 200113
rect 46811 200085 46839 200113
rect 46625 200023 46653 200051
rect 46687 200023 46715 200051
rect 46749 200023 46777 200051
rect 46811 200023 46839 200051
rect 46625 199961 46653 199989
rect 46687 199961 46715 199989
rect 46749 199961 46777 199989
rect 46811 199961 46839 199989
rect 46625 191147 46653 191175
rect 46687 191147 46715 191175
rect 46749 191147 46777 191175
rect 46811 191147 46839 191175
rect 46625 191085 46653 191113
rect 46687 191085 46715 191113
rect 46749 191085 46777 191113
rect 46811 191085 46839 191113
rect 46625 191023 46653 191051
rect 46687 191023 46715 191051
rect 46749 191023 46777 191051
rect 46811 191023 46839 191051
rect 46625 190961 46653 190989
rect 46687 190961 46715 190989
rect 46749 190961 46777 190989
rect 46811 190961 46839 190989
rect 46625 182147 46653 182175
rect 46687 182147 46715 182175
rect 46749 182147 46777 182175
rect 46811 182147 46839 182175
rect 46625 182085 46653 182113
rect 46687 182085 46715 182113
rect 46749 182085 46777 182113
rect 46811 182085 46839 182113
rect 46625 182023 46653 182051
rect 46687 182023 46715 182051
rect 46749 182023 46777 182051
rect 46811 182023 46839 182051
rect 46625 181961 46653 181989
rect 46687 181961 46715 181989
rect 46749 181961 46777 181989
rect 46811 181961 46839 181989
rect 46625 173147 46653 173175
rect 46687 173147 46715 173175
rect 46749 173147 46777 173175
rect 46811 173147 46839 173175
rect 46625 173085 46653 173113
rect 46687 173085 46715 173113
rect 46749 173085 46777 173113
rect 46811 173085 46839 173113
rect 46625 173023 46653 173051
rect 46687 173023 46715 173051
rect 46749 173023 46777 173051
rect 46811 173023 46839 173051
rect 46625 172961 46653 172989
rect 46687 172961 46715 172989
rect 46749 172961 46777 172989
rect 46811 172961 46839 172989
rect 46625 164147 46653 164175
rect 46687 164147 46715 164175
rect 46749 164147 46777 164175
rect 46811 164147 46839 164175
rect 46625 164085 46653 164113
rect 46687 164085 46715 164113
rect 46749 164085 46777 164113
rect 46811 164085 46839 164113
rect 46625 164023 46653 164051
rect 46687 164023 46715 164051
rect 46749 164023 46777 164051
rect 46811 164023 46839 164051
rect 46625 163961 46653 163989
rect 46687 163961 46715 163989
rect 46749 163961 46777 163989
rect 46811 163961 46839 163989
rect 46625 155147 46653 155175
rect 46687 155147 46715 155175
rect 46749 155147 46777 155175
rect 46811 155147 46839 155175
rect 46625 155085 46653 155113
rect 46687 155085 46715 155113
rect 46749 155085 46777 155113
rect 46811 155085 46839 155113
rect 46625 155023 46653 155051
rect 46687 155023 46715 155051
rect 46749 155023 46777 155051
rect 46811 155023 46839 155051
rect 46625 154961 46653 154989
rect 46687 154961 46715 154989
rect 46749 154961 46777 154989
rect 46811 154961 46839 154989
rect 46625 146147 46653 146175
rect 46687 146147 46715 146175
rect 46749 146147 46777 146175
rect 46811 146147 46839 146175
rect 46625 146085 46653 146113
rect 46687 146085 46715 146113
rect 46749 146085 46777 146113
rect 46811 146085 46839 146113
rect 46625 146023 46653 146051
rect 46687 146023 46715 146051
rect 46749 146023 46777 146051
rect 46811 146023 46839 146051
rect 46625 145961 46653 145989
rect 46687 145961 46715 145989
rect 46749 145961 46777 145989
rect 46811 145961 46839 145989
rect 46625 137147 46653 137175
rect 46687 137147 46715 137175
rect 46749 137147 46777 137175
rect 46811 137147 46839 137175
rect 46625 137085 46653 137113
rect 46687 137085 46715 137113
rect 46749 137085 46777 137113
rect 46811 137085 46839 137113
rect 46625 137023 46653 137051
rect 46687 137023 46715 137051
rect 46749 137023 46777 137051
rect 46811 137023 46839 137051
rect 46625 136961 46653 136989
rect 46687 136961 46715 136989
rect 46749 136961 46777 136989
rect 46811 136961 46839 136989
rect 46625 128147 46653 128175
rect 46687 128147 46715 128175
rect 46749 128147 46777 128175
rect 46811 128147 46839 128175
rect 46625 128085 46653 128113
rect 46687 128085 46715 128113
rect 46749 128085 46777 128113
rect 46811 128085 46839 128113
rect 46625 128023 46653 128051
rect 46687 128023 46715 128051
rect 46749 128023 46777 128051
rect 46811 128023 46839 128051
rect 46625 127961 46653 127989
rect 46687 127961 46715 127989
rect 46749 127961 46777 127989
rect 46811 127961 46839 127989
rect 46625 119147 46653 119175
rect 46687 119147 46715 119175
rect 46749 119147 46777 119175
rect 46811 119147 46839 119175
rect 46625 119085 46653 119113
rect 46687 119085 46715 119113
rect 46749 119085 46777 119113
rect 46811 119085 46839 119113
rect 46625 119023 46653 119051
rect 46687 119023 46715 119051
rect 46749 119023 46777 119051
rect 46811 119023 46839 119051
rect 46625 118961 46653 118989
rect 46687 118961 46715 118989
rect 46749 118961 46777 118989
rect 46811 118961 46839 118989
rect 46625 110147 46653 110175
rect 46687 110147 46715 110175
rect 46749 110147 46777 110175
rect 46811 110147 46839 110175
rect 46625 110085 46653 110113
rect 46687 110085 46715 110113
rect 46749 110085 46777 110113
rect 46811 110085 46839 110113
rect 46625 110023 46653 110051
rect 46687 110023 46715 110051
rect 46749 110023 46777 110051
rect 46811 110023 46839 110051
rect 46625 109961 46653 109989
rect 46687 109961 46715 109989
rect 46749 109961 46777 109989
rect 46811 109961 46839 109989
rect 46625 101147 46653 101175
rect 46687 101147 46715 101175
rect 46749 101147 46777 101175
rect 46811 101147 46839 101175
rect 46625 101085 46653 101113
rect 46687 101085 46715 101113
rect 46749 101085 46777 101113
rect 46811 101085 46839 101113
rect 46625 101023 46653 101051
rect 46687 101023 46715 101051
rect 46749 101023 46777 101051
rect 46811 101023 46839 101051
rect 46625 100961 46653 100989
rect 46687 100961 46715 100989
rect 46749 100961 46777 100989
rect 46811 100961 46839 100989
rect 46625 92147 46653 92175
rect 46687 92147 46715 92175
rect 46749 92147 46777 92175
rect 46811 92147 46839 92175
rect 46625 92085 46653 92113
rect 46687 92085 46715 92113
rect 46749 92085 46777 92113
rect 46811 92085 46839 92113
rect 46625 92023 46653 92051
rect 46687 92023 46715 92051
rect 46749 92023 46777 92051
rect 46811 92023 46839 92051
rect 46625 91961 46653 91989
rect 46687 91961 46715 91989
rect 46749 91961 46777 91989
rect 46811 91961 46839 91989
rect 46625 83147 46653 83175
rect 46687 83147 46715 83175
rect 46749 83147 46777 83175
rect 46811 83147 46839 83175
rect 46625 83085 46653 83113
rect 46687 83085 46715 83113
rect 46749 83085 46777 83113
rect 46811 83085 46839 83113
rect 46625 83023 46653 83051
rect 46687 83023 46715 83051
rect 46749 83023 46777 83051
rect 46811 83023 46839 83051
rect 46625 82961 46653 82989
rect 46687 82961 46715 82989
rect 46749 82961 46777 82989
rect 46811 82961 46839 82989
rect 46625 74147 46653 74175
rect 46687 74147 46715 74175
rect 46749 74147 46777 74175
rect 46811 74147 46839 74175
rect 46625 74085 46653 74113
rect 46687 74085 46715 74113
rect 46749 74085 46777 74113
rect 46811 74085 46839 74113
rect 46625 74023 46653 74051
rect 46687 74023 46715 74051
rect 46749 74023 46777 74051
rect 46811 74023 46839 74051
rect 46625 73961 46653 73989
rect 46687 73961 46715 73989
rect 46749 73961 46777 73989
rect 46811 73961 46839 73989
rect 46625 65147 46653 65175
rect 46687 65147 46715 65175
rect 46749 65147 46777 65175
rect 46811 65147 46839 65175
rect 46625 65085 46653 65113
rect 46687 65085 46715 65113
rect 46749 65085 46777 65113
rect 46811 65085 46839 65113
rect 46625 65023 46653 65051
rect 46687 65023 46715 65051
rect 46749 65023 46777 65051
rect 46811 65023 46839 65051
rect 46625 64961 46653 64989
rect 46687 64961 46715 64989
rect 46749 64961 46777 64989
rect 46811 64961 46839 64989
rect 46625 56147 46653 56175
rect 46687 56147 46715 56175
rect 46749 56147 46777 56175
rect 46811 56147 46839 56175
rect 46625 56085 46653 56113
rect 46687 56085 46715 56113
rect 46749 56085 46777 56113
rect 46811 56085 46839 56113
rect 46625 56023 46653 56051
rect 46687 56023 46715 56051
rect 46749 56023 46777 56051
rect 46811 56023 46839 56051
rect 46625 55961 46653 55989
rect 46687 55961 46715 55989
rect 46749 55961 46777 55989
rect 46811 55961 46839 55989
rect 46625 47147 46653 47175
rect 46687 47147 46715 47175
rect 46749 47147 46777 47175
rect 46811 47147 46839 47175
rect 46625 47085 46653 47113
rect 46687 47085 46715 47113
rect 46749 47085 46777 47113
rect 46811 47085 46839 47113
rect 46625 47023 46653 47051
rect 46687 47023 46715 47051
rect 46749 47023 46777 47051
rect 46811 47023 46839 47051
rect 46625 46961 46653 46989
rect 46687 46961 46715 46989
rect 46749 46961 46777 46989
rect 46811 46961 46839 46989
rect 46625 38147 46653 38175
rect 46687 38147 46715 38175
rect 46749 38147 46777 38175
rect 46811 38147 46839 38175
rect 46625 38085 46653 38113
rect 46687 38085 46715 38113
rect 46749 38085 46777 38113
rect 46811 38085 46839 38113
rect 46625 38023 46653 38051
rect 46687 38023 46715 38051
rect 46749 38023 46777 38051
rect 46811 38023 46839 38051
rect 46625 37961 46653 37989
rect 46687 37961 46715 37989
rect 46749 37961 46777 37989
rect 46811 37961 46839 37989
rect 46625 29147 46653 29175
rect 46687 29147 46715 29175
rect 46749 29147 46777 29175
rect 46811 29147 46839 29175
rect 46625 29085 46653 29113
rect 46687 29085 46715 29113
rect 46749 29085 46777 29113
rect 46811 29085 46839 29113
rect 46625 29023 46653 29051
rect 46687 29023 46715 29051
rect 46749 29023 46777 29051
rect 46811 29023 46839 29051
rect 46625 28961 46653 28989
rect 46687 28961 46715 28989
rect 46749 28961 46777 28989
rect 46811 28961 46839 28989
rect 46625 20147 46653 20175
rect 46687 20147 46715 20175
rect 46749 20147 46777 20175
rect 46811 20147 46839 20175
rect 46625 20085 46653 20113
rect 46687 20085 46715 20113
rect 46749 20085 46777 20113
rect 46811 20085 46839 20113
rect 46625 20023 46653 20051
rect 46687 20023 46715 20051
rect 46749 20023 46777 20051
rect 46811 20023 46839 20051
rect 46625 19961 46653 19989
rect 46687 19961 46715 19989
rect 46749 19961 46777 19989
rect 46811 19961 46839 19989
rect 46625 11147 46653 11175
rect 46687 11147 46715 11175
rect 46749 11147 46777 11175
rect 46811 11147 46839 11175
rect 46625 11085 46653 11113
rect 46687 11085 46715 11113
rect 46749 11085 46777 11113
rect 46811 11085 46839 11113
rect 46625 11023 46653 11051
rect 46687 11023 46715 11051
rect 46749 11023 46777 11051
rect 46811 11023 46839 11051
rect 46625 10961 46653 10989
rect 46687 10961 46715 10989
rect 46749 10961 46777 10989
rect 46811 10961 46839 10989
rect 46625 2147 46653 2175
rect 46687 2147 46715 2175
rect 46749 2147 46777 2175
rect 46811 2147 46839 2175
rect 46625 2085 46653 2113
rect 46687 2085 46715 2113
rect 46749 2085 46777 2113
rect 46811 2085 46839 2113
rect 46625 2023 46653 2051
rect 46687 2023 46715 2051
rect 46749 2023 46777 2051
rect 46811 2023 46839 2051
rect 46625 1961 46653 1989
rect 46687 1961 46715 1989
rect 46749 1961 46777 1989
rect 46811 1961 46839 1989
rect 46625 -108 46653 -80
rect 46687 -108 46715 -80
rect 46749 -108 46777 -80
rect 46811 -108 46839 -80
rect 46625 -170 46653 -142
rect 46687 -170 46715 -142
rect 46749 -170 46777 -142
rect 46811 -170 46839 -142
rect 46625 -232 46653 -204
rect 46687 -232 46715 -204
rect 46749 -232 46777 -204
rect 46811 -232 46839 -204
rect 46625 -294 46653 -266
rect 46687 -294 46715 -266
rect 46749 -294 46777 -266
rect 46811 -294 46839 -266
rect 48485 299058 48513 299086
rect 48547 299058 48575 299086
rect 48609 299058 48637 299086
rect 48671 299058 48699 299086
rect 48485 298996 48513 299024
rect 48547 298996 48575 299024
rect 48609 298996 48637 299024
rect 48671 298996 48699 299024
rect 48485 298934 48513 298962
rect 48547 298934 48575 298962
rect 48609 298934 48637 298962
rect 48671 298934 48699 298962
rect 48485 298872 48513 298900
rect 48547 298872 48575 298900
rect 48609 298872 48637 298900
rect 48671 298872 48699 298900
rect 48485 293147 48513 293175
rect 48547 293147 48575 293175
rect 48609 293147 48637 293175
rect 48671 293147 48699 293175
rect 48485 293085 48513 293113
rect 48547 293085 48575 293113
rect 48609 293085 48637 293113
rect 48671 293085 48699 293113
rect 48485 293023 48513 293051
rect 48547 293023 48575 293051
rect 48609 293023 48637 293051
rect 48671 293023 48699 293051
rect 48485 292961 48513 292989
rect 48547 292961 48575 292989
rect 48609 292961 48637 292989
rect 48671 292961 48699 292989
rect 48485 284147 48513 284175
rect 48547 284147 48575 284175
rect 48609 284147 48637 284175
rect 48671 284147 48699 284175
rect 48485 284085 48513 284113
rect 48547 284085 48575 284113
rect 48609 284085 48637 284113
rect 48671 284085 48699 284113
rect 48485 284023 48513 284051
rect 48547 284023 48575 284051
rect 48609 284023 48637 284051
rect 48671 284023 48699 284051
rect 48485 283961 48513 283989
rect 48547 283961 48575 283989
rect 48609 283961 48637 283989
rect 48671 283961 48699 283989
rect 48485 275147 48513 275175
rect 48547 275147 48575 275175
rect 48609 275147 48637 275175
rect 48671 275147 48699 275175
rect 48485 275085 48513 275113
rect 48547 275085 48575 275113
rect 48609 275085 48637 275113
rect 48671 275085 48699 275113
rect 48485 275023 48513 275051
rect 48547 275023 48575 275051
rect 48609 275023 48637 275051
rect 48671 275023 48699 275051
rect 48485 274961 48513 274989
rect 48547 274961 48575 274989
rect 48609 274961 48637 274989
rect 48671 274961 48699 274989
rect 48485 266147 48513 266175
rect 48547 266147 48575 266175
rect 48609 266147 48637 266175
rect 48671 266147 48699 266175
rect 48485 266085 48513 266113
rect 48547 266085 48575 266113
rect 48609 266085 48637 266113
rect 48671 266085 48699 266113
rect 48485 266023 48513 266051
rect 48547 266023 48575 266051
rect 48609 266023 48637 266051
rect 48671 266023 48699 266051
rect 48485 265961 48513 265989
rect 48547 265961 48575 265989
rect 48609 265961 48637 265989
rect 48671 265961 48699 265989
rect 55625 298578 55653 298606
rect 55687 298578 55715 298606
rect 55749 298578 55777 298606
rect 55811 298578 55839 298606
rect 55625 298516 55653 298544
rect 55687 298516 55715 298544
rect 55749 298516 55777 298544
rect 55811 298516 55839 298544
rect 55625 298454 55653 298482
rect 55687 298454 55715 298482
rect 55749 298454 55777 298482
rect 55811 298454 55839 298482
rect 55625 298392 55653 298420
rect 55687 298392 55715 298420
rect 55749 298392 55777 298420
rect 55811 298392 55839 298420
rect 55625 290147 55653 290175
rect 55687 290147 55715 290175
rect 55749 290147 55777 290175
rect 55811 290147 55839 290175
rect 55625 290085 55653 290113
rect 55687 290085 55715 290113
rect 55749 290085 55777 290113
rect 55811 290085 55839 290113
rect 55625 290023 55653 290051
rect 55687 290023 55715 290051
rect 55749 290023 55777 290051
rect 55811 290023 55839 290051
rect 55625 289961 55653 289989
rect 55687 289961 55715 289989
rect 55749 289961 55777 289989
rect 55811 289961 55839 289989
rect 55625 281147 55653 281175
rect 55687 281147 55715 281175
rect 55749 281147 55777 281175
rect 55811 281147 55839 281175
rect 55625 281085 55653 281113
rect 55687 281085 55715 281113
rect 55749 281085 55777 281113
rect 55811 281085 55839 281113
rect 55625 281023 55653 281051
rect 55687 281023 55715 281051
rect 55749 281023 55777 281051
rect 55811 281023 55839 281051
rect 55625 280961 55653 280989
rect 55687 280961 55715 280989
rect 55749 280961 55777 280989
rect 55811 280961 55839 280989
rect 55625 272147 55653 272175
rect 55687 272147 55715 272175
rect 55749 272147 55777 272175
rect 55811 272147 55839 272175
rect 55625 272085 55653 272113
rect 55687 272085 55715 272113
rect 55749 272085 55777 272113
rect 55811 272085 55839 272113
rect 55625 272023 55653 272051
rect 55687 272023 55715 272051
rect 55749 272023 55777 272051
rect 55811 272023 55839 272051
rect 55625 271961 55653 271989
rect 55687 271961 55715 271989
rect 55749 271961 55777 271989
rect 55811 271961 55839 271989
rect 55625 263147 55653 263175
rect 55687 263147 55715 263175
rect 55749 263147 55777 263175
rect 55811 263147 55839 263175
rect 55625 263085 55653 263113
rect 55687 263085 55715 263113
rect 55749 263085 55777 263113
rect 55811 263085 55839 263113
rect 55625 263023 55653 263051
rect 55687 263023 55715 263051
rect 55749 263023 55777 263051
rect 55811 263023 55839 263051
rect 55625 262961 55653 262989
rect 55687 262961 55715 262989
rect 55749 262961 55777 262989
rect 55811 262961 55839 262989
rect 57485 299058 57513 299086
rect 57547 299058 57575 299086
rect 57609 299058 57637 299086
rect 57671 299058 57699 299086
rect 57485 298996 57513 299024
rect 57547 298996 57575 299024
rect 57609 298996 57637 299024
rect 57671 298996 57699 299024
rect 57485 298934 57513 298962
rect 57547 298934 57575 298962
rect 57609 298934 57637 298962
rect 57671 298934 57699 298962
rect 57485 298872 57513 298900
rect 57547 298872 57575 298900
rect 57609 298872 57637 298900
rect 57671 298872 57699 298900
rect 57485 293147 57513 293175
rect 57547 293147 57575 293175
rect 57609 293147 57637 293175
rect 57671 293147 57699 293175
rect 57485 293085 57513 293113
rect 57547 293085 57575 293113
rect 57609 293085 57637 293113
rect 57671 293085 57699 293113
rect 57485 293023 57513 293051
rect 57547 293023 57575 293051
rect 57609 293023 57637 293051
rect 57671 293023 57699 293051
rect 57485 292961 57513 292989
rect 57547 292961 57575 292989
rect 57609 292961 57637 292989
rect 57671 292961 57699 292989
rect 57485 284147 57513 284175
rect 57547 284147 57575 284175
rect 57609 284147 57637 284175
rect 57671 284147 57699 284175
rect 57485 284085 57513 284113
rect 57547 284085 57575 284113
rect 57609 284085 57637 284113
rect 57671 284085 57699 284113
rect 57485 284023 57513 284051
rect 57547 284023 57575 284051
rect 57609 284023 57637 284051
rect 57671 284023 57699 284051
rect 57485 283961 57513 283989
rect 57547 283961 57575 283989
rect 57609 283961 57637 283989
rect 57671 283961 57699 283989
rect 57485 275147 57513 275175
rect 57547 275147 57575 275175
rect 57609 275147 57637 275175
rect 57671 275147 57699 275175
rect 57485 275085 57513 275113
rect 57547 275085 57575 275113
rect 57609 275085 57637 275113
rect 57671 275085 57699 275113
rect 57485 275023 57513 275051
rect 57547 275023 57575 275051
rect 57609 275023 57637 275051
rect 57671 275023 57699 275051
rect 57485 274961 57513 274989
rect 57547 274961 57575 274989
rect 57609 274961 57637 274989
rect 57671 274961 57699 274989
rect 57485 266147 57513 266175
rect 57547 266147 57575 266175
rect 57609 266147 57637 266175
rect 57671 266147 57699 266175
rect 57485 266085 57513 266113
rect 57547 266085 57575 266113
rect 57609 266085 57637 266113
rect 57671 266085 57699 266113
rect 57485 266023 57513 266051
rect 57547 266023 57575 266051
rect 57609 266023 57637 266051
rect 57671 266023 57699 266051
rect 57485 265961 57513 265989
rect 57547 265961 57575 265989
rect 57609 265961 57637 265989
rect 57671 265961 57699 265989
rect 64625 298578 64653 298606
rect 64687 298578 64715 298606
rect 64749 298578 64777 298606
rect 64811 298578 64839 298606
rect 64625 298516 64653 298544
rect 64687 298516 64715 298544
rect 64749 298516 64777 298544
rect 64811 298516 64839 298544
rect 64625 298454 64653 298482
rect 64687 298454 64715 298482
rect 64749 298454 64777 298482
rect 64811 298454 64839 298482
rect 64625 298392 64653 298420
rect 64687 298392 64715 298420
rect 64749 298392 64777 298420
rect 64811 298392 64839 298420
rect 64625 290147 64653 290175
rect 64687 290147 64715 290175
rect 64749 290147 64777 290175
rect 64811 290147 64839 290175
rect 64625 290085 64653 290113
rect 64687 290085 64715 290113
rect 64749 290085 64777 290113
rect 64811 290085 64839 290113
rect 64625 290023 64653 290051
rect 64687 290023 64715 290051
rect 64749 290023 64777 290051
rect 64811 290023 64839 290051
rect 64625 289961 64653 289989
rect 64687 289961 64715 289989
rect 64749 289961 64777 289989
rect 64811 289961 64839 289989
rect 64625 281147 64653 281175
rect 64687 281147 64715 281175
rect 64749 281147 64777 281175
rect 64811 281147 64839 281175
rect 64625 281085 64653 281113
rect 64687 281085 64715 281113
rect 64749 281085 64777 281113
rect 64811 281085 64839 281113
rect 64625 281023 64653 281051
rect 64687 281023 64715 281051
rect 64749 281023 64777 281051
rect 64811 281023 64839 281051
rect 64625 280961 64653 280989
rect 64687 280961 64715 280989
rect 64749 280961 64777 280989
rect 64811 280961 64839 280989
rect 64625 272147 64653 272175
rect 64687 272147 64715 272175
rect 64749 272147 64777 272175
rect 64811 272147 64839 272175
rect 64625 272085 64653 272113
rect 64687 272085 64715 272113
rect 64749 272085 64777 272113
rect 64811 272085 64839 272113
rect 64625 272023 64653 272051
rect 64687 272023 64715 272051
rect 64749 272023 64777 272051
rect 64811 272023 64839 272051
rect 64625 271961 64653 271989
rect 64687 271961 64715 271989
rect 64749 271961 64777 271989
rect 64811 271961 64839 271989
rect 64625 263147 64653 263175
rect 64687 263147 64715 263175
rect 64749 263147 64777 263175
rect 64811 263147 64839 263175
rect 64625 263085 64653 263113
rect 64687 263085 64715 263113
rect 64749 263085 64777 263113
rect 64811 263085 64839 263113
rect 64625 263023 64653 263051
rect 64687 263023 64715 263051
rect 64749 263023 64777 263051
rect 64811 263023 64839 263051
rect 64625 262961 64653 262989
rect 64687 262961 64715 262989
rect 64749 262961 64777 262989
rect 64811 262961 64839 262989
rect 66485 299058 66513 299086
rect 66547 299058 66575 299086
rect 66609 299058 66637 299086
rect 66671 299058 66699 299086
rect 66485 298996 66513 299024
rect 66547 298996 66575 299024
rect 66609 298996 66637 299024
rect 66671 298996 66699 299024
rect 66485 298934 66513 298962
rect 66547 298934 66575 298962
rect 66609 298934 66637 298962
rect 66671 298934 66699 298962
rect 66485 298872 66513 298900
rect 66547 298872 66575 298900
rect 66609 298872 66637 298900
rect 66671 298872 66699 298900
rect 66485 293147 66513 293175
rect 66547 293147 66575 293175
rect 66609 293147 66637 293175
rect 66671 293147 66699 293175
rect 66485 293085 66513 293113
rect 66547 293085 66575 293113
rect 66609 293085 66637 293113
rect 66671 293085 66699 293113
rect 66485 293023 66513 293051
rect 66547 293023 66575 293051
rect 66609 293023 66637 293051
rect 66671 293023 66699 293051
rect 66485 292961 66513 292989
rect 66547 292961 66575 292989
rect 66609 292961 66637 292989
rect 66671 292961 66699 292989
rect 66485 284147 66513 284175
rect 66547 284147 66575 284175
rect 66609 284147 66637 284175
rect 66671 284147 66699 284175
rect 66485 284085 66513 284113
rect 66547 284085 66575 284113
rect 66609 284085 66637 284113
rect 66671 284085 66699 284113
rect 66485 284023 66513 284051
rect 66547 284023 66575 284051
rect 66609 284023 66637 284051
rect 66671 284023 66699 284051
rect 66485 283961 66513 283989
rect 66547 283961 66575 283989
rect 66609 283961 66637 283989
rect 66671 283961 66699 283989
rect 66485 275147 66513 275175
rect 66547 275147 66575 275175
rect 66609 275147 66637 275175
rect 66671 275147 66699 275175
rect 66485 275085 66513 275113
rect 66547 275085 66575 275113
rect 66609 275085 66637 275113
rect 66671 275085 66699 275113
rect 66485 275023 66513 275051
rect 66547 275023 66575 275051
rect 66609 275023 66637 275051
rect 66671 275023 66699 275051
rect 66485 274961 66513 274989
rect 66547 274961 66575 274989
rect 66609 274961 66637 274989
rect 66671 274961 66699 274989
rect 66485 266147 66513 266175
rect 66547 266147 66575 266175
rect 66609 266147 66637 266175
rect 66671 266147 66699 266175
rect 66485 266085 66513 266113
rect 66547 266085 66575 266113
rect 66609 266085 66637 266113
rect 66671 266085 66699 266113
rect 66485 266023 66513 266051
rect 66547 266023 66575 266051
rect 66609 266023 66637 266051
rect 66671 266023 66699 266051
rect 66485 265961 66513 265989
rect 66547 265961 66575 265989
rect 66609 265961 66637 265989
rect 66671 265961 66699 265989
rect 73625 298578 73653 298606
rect 73687 298578 73715 298606
rect 73749 298578 73777 298606
rect 73811 298578 73839 298606
rect 73625 298516 73653 298544
rect 73687 298516 73715 298544
rect 73749 298516 73777 298544
rect 73811 298516 73839 298544
rect 73625 298454 73653 298482
rect 73687 298454 73715 298482
rect 73749 298454 73777 298482
rect 73811 298454 73839 298482
rect 73625 298392 73653 298420
rect 73687 298392 73715 298420
rect 73749 298392 73777 298420
rect 73811 298392 73839 298420
rect 73625 290147 73653 290175
rect 73687 290147 73715 290175
rect 73749 290147 73777 290175
rect 73811 290147 73839 290175
rect 73625 290085 73653 290113
rect 73687 290085 73715 290113
rect 73749 290085 73777 290113
rect 73811 290085 73839 290113
rect 73625 290023 73653 290051
rect 73687 290023 73715 290051
rect 73749 290023 73777 290051
rect 73811 290023 73839 290051
rect 73625 289961 73653 289989
rect 73687 289961 73715 289989
rect 73749 289961 73777 289989
rect 73811 289961 73839 289989
rect 73625 281147 73653 281175
rect 73687 281147 73715 281175
rect 73749 281147 73777 281175
rect 73811 281147 73839 281175
rect 73625 281085 73653 281113
rect 73687 281085 73715 281113
rect 73749 281085 73777 281113
rect 73811 281085 73839 281113
rect 73625 281023 73653 281051
rect 73687 281023 73715 281051
rect 73749 281023 73777 281051
rect 73811 281023 73839 281051
rect 73625 280961 73653 280989
rect 73687 280961 73715 280989
rect 73749 280961 73777 280989
rect 73811 280961 73839 280989
rect 73625 272147 73653 272175
rect 73687 272147 73715 272175
rect 73749 272147 73777 272175
rect 73811 272147 73839 272175
rect 73625 272085 73653 272113
rect 73687 272085 73715 272113
rect 73749 272085 73777 272113
rect 73811 272085 73839 272113
rect 73625 272023 73653 272051
rect 73687 272023 73715 272051
rect 73749 272023 73777 272051
rect 73811 272023 73839 272051
rect 73625 271961 73653 271989
rect 73687 271961 73715 271989
rect 73749 271961 73777 271989
rect 73811 271961 73839 271989
rect 73625 263147 73653 263175
rect 73687 263147 73715 263175
rect 73749 263147 73777 263175
rect 73811 263147 73839 263175
rect 73625 263085 73653 263113
rect 73687 263085 73715 263113
rect 73749 263085 73777 263113
rect 73811 263085 73839 263113
rect 73625 263023 73653 263051
rect 73687 263023 73715 263051
rect 73749 263023 73777 263051
rect 73811 263023 73839 263051
rect 73625 262961 73653 262989
rect 73687 262961 73715 262989
rect 73749 262961 73777 262989
rect 73811 262961 73839 262989
rect 75485 299058 75513 299086
rect 75547 299058 75575 299086
rect 75609 299058 75637 299086
rect 75671 299058 75699 299086
rect 75485 298996 75513 299024
rect 75547 298996 75575 299024
rect 75609 298996 75637 299024
rect 75671 298996 75699 299024
rect 75485 298934 75513 298962
rect 75547 298934 75575 298962
rect 75609 298934 75637 298962
rect 75671 298934 75699 298962
rect 75485 298872 75513 298900
rect 75547 298872 75575 298900
rect 75609 298872 75637 298900
rect 75671 298872 75699 298900
rect 75485 293147 75513 293175
rect 75547 293147 75575 293175
rect 75609 293147 75637 293175
rect 75671 293147 75699 293175
rect 75485 293085 75513 293113
rect 75547 293085 75575 293113
rect 75609 293085 75637 293113
rect 75671 293085 75699 293113
rect 75485 293023 75513 293051
rect 75547 293023 75575 293051
rect 75609 293023 75637 293051
rect 75671 293023 75699 293051
rect 75485 292961 75513 292989
rect 75547 292961 75575 292989
rect 75609 292961 75637 292989
rect 75671 292961 75699 292989
rect 75485 284147 75513 284175
rect 75547 284147 75575 284175
rect 75609 284147 75637 284175
rect 75671 284147 75699 284175
rect 75485 284085 75513 284113
rect 75547 284085 75575 284113
rect 75609 284085 75637 284113
rect 75671 284085 75699 284113
rect 75485 284023 75513 284051
rect 75547 284023 75575 284051
rect 75609 284023 75637 284051
rect 75671 284023 75699 284051
rect 75485 283961 75513 283989
rect 75547 283961 75575 283989
rect 75609 283961 75637 283989
rect 75671 283961 75699 283989
rect 75485 275147 75513 275175
rect 75547 275147 75575 275175
rect 75609 275147 75637 275175
rect 75671 275147 75699 275175
rect 75485 275085 75513 275113
rect 75547 275085 75575 275113
rect 75609 275085 75637 275113
rect 75671 275085 75699 275113
rect 75485 275023 75513 275051
rect 75547 275023 75575 275051
rect 75609 275023 75637 275051
rect 75671 275023 75699 275051
rect 75485 274961 75513 274989
rect 75547 274961 75575 274989
rect 75609 274961 75637 274989
rect 75671 274961 75699 274989
rect 75485 266147 75513 266175
rect 75547 266147 75575 266175
rect 75609 266147 75637 266175
rect 75671 266147 75699 266175
rect 75485 266085 75513 266113
rect 75547 266085 75575 266113
rect 75609 266085 75637 266113
rect 75671 266085 75699 266113
rect 75485 266023 75513 266051
rect 75547 266023 75575 266051
rect 75609 266023 75637 266051
rect 75671 266023 75699 266051
rect 75485 265961 75513 265989
rect 75547 265961 75575 265989
rect 75609 265961 75637 265989
rect 75671 265961 75699 265989
rect 82625 298578 82653 298606
rect 82687 298578 82715 298606
rect 82749 298578 82777 298606
rect 82811 298578 82839 298606
rect 82625 298516 82653 298544
rect 82687 298516 82715 298544
rect 82749 298516 82777 298544
rect 82811 298516 82839 298544
rect 82625 298454 82653 298482
rect 82687 298454 82715 298482
rect 82749 298454 82777 298482
rect 82811 298454 82839 298482
rect 82625 298392 82653 298420
rect 82687 298392 82715 298420
rect 82749 298392 82777 298420
rect 82811 298392 82839 298420
rect 82625 290147 82653 290175
rect 82687 290147 82715 290175
rect 82749 290147 82777 290175
rect 82811 290147 82839 290175
rect 82625 290085 82653 290113
rect 82687 290085 82715 290113
rect 82749 290085 82777 290113
rect 82811 290085 82839 290113
rect 82625 290023 82653 290051
rect 82687 290023 82715 290051
rect 82749 290023 82777 290051
rect 82811 290023 82839 290051
rect 82625 289961 82653 289989
rect 82687 289961 82715 289989
rect 82749 289961 82777 289989
rect 82811 289961 82839 289989
rect 82625 281147 82653 281175
rect 82687 281147 82715 281175
rect 82749 281147 82777 281175
rect 82811 281147 82839 281175
rect 82625 281085 82653 281113
rect 82687 281085 82715 281113
rect 82749 281085 82777 281113
rect 82811 281085 82839 281113
rect 82625 281023 82653 281051
rect 82687 281023 82715 281051
rect 82749 281023 82777 281051
rect 82811 281023 82839 281051
rect 82625 280961 82653 280989
rect 82687 280961 82715 280989
rect 82749 280961 82777 280989
rect 82811 280961 82839 280989
rect 82625 272147 82653 272175
rect 82687 272147 82715 272175
rect 82749 272147 82777 272175
rect 82811 272147 82839 272175
rect 82625 272085 82653 272113
rect 82687 272085 82715 272113
rect 82749 272085 82777 272113
rect 82811 272085 82839 272113
rect 82625 272023 82653 272051
rect 82687 272023 82715 272051
rect 82749 272023 82777 272051
rect 82811 272023 82839 272051
rect 82625 271961 82653 271989
rect 82687 271961 82715 271989
rect 82749 271961 82777 271989
rect 82811 271961 82839 271989
rect 82625 263147 82653 263175
rect 82687 263147 82715 263175
rect 82749 263147 82777 263175
rect 82811 263147 82839 263175
rect 82625 263085 82653 263113
rect 82687 263085 82715 263113
rect 82749 263085 82777 263113
rect 82811 263085 82839 263113
rect 82625 263023 82653 263051
rect 82687 263023 82715 263051
rect 82749 263023 82777 263051
rect 82811 263023 82839 263051
rect 82625 262961 82653 262989
rect 82687 262961 82715 262989
rect 82749 262961 82777 262989
rect 82811 262961 82839 262989
rect 84485 299058 84513 299086
rect 84547 299058 84575 299086
rect 84609 299058 84637 299086
rect 84671 299058 84699 299086
rect 84485 298996 84513 299024
rect 84547 298996 84575 299024
rect 84609 298996 84637 299024
rect 84671 298996 84699 299024
rect 84485 298934 84513 298962
rect 84547 298934 84575 298962
rect 84609 298934 84637 298962
rect 84671 298934 84699 298962
rect 84485 298872 84513 298900
rect 84547 298872 84575 298900
rect 84609 298872 84637 298900
rect 84671 298872 84699 298900
rect 84485 293147 84513 293175
rect 84547 293147 84575 293175
rect 84609 293147 84637 293175
rect 84671 293147 84699 293175
rect 84485 293085 84513 293113
rect 84547 293085 84575 293113
rect 84609 293085 84637 293113
rect 84671 293085 84699 293113
rect 84485 293023 84513 293051
rect 84547 293023 84575 293051
rect 84609 293023 84637 293051
rect 84671 293023 84699 293051
rect 84485 292961 84513 292989
rect 84547 292961 84575 292989
rect 84609 292961 84637 292989
rect 84671 292961 84699 292989
rect 84485 284147 84513 284175
rect 84547 284147 84575 284175
rect 84609 284147 84637 284175
rect 84671 284147 84699 284175
rect 84485 284085 84513 284113
rect 84547 284085 84575 284113
rect 84609 284085 84637 284113
rect 84671 284085 84699 284113
rect 84485 284023 84513 284051
rect 84547 284023 84575 284051
rect 84609 284023 84637 284051
rect 84671 284023 84699 284051
rect 84485 283961 84513 283989
rect 84547 283961 84575 283989
rect 84609 283961 84637 283989
rect 84671 283961 84699 283989
rect 84485 275147 84513 275175
rect 84547 275147 84575 275175
rect 84609 275147 84637 275175
rect 84671 275147 84699 275175
rect 84485 275085 84513 275113
rect 84547 275085 84575 275113
rect 84609 275085 84637 275113
rect 84671 275085 84699 275113
rect 84485 275023 84513 275051
rect 84547 275023 84575 275051
rect 84609 275023 84637 275051
rect 84671 275023 84699 275051
rect 84485 274961 84513 274989
rect 84547 274961 84575 274989
rect 84609 274961 84637 274989
rect 84671 274961 84699 274989
rect 84485 266147 84513 266175
rect 84547 266147 84575 266175
rect 84609 266147 84637 266175
rect 84671 266147 84699 266175
rect 84485 266085 84513 266113
rect 84547 266085 84575 266113
rect 84609 266085 84637 266113
rect 84671 266085 84699 266113
rect 84485 266023 84513 266051
rect 84547 266023 84575 266051
rect 84609 266023 84637 266051
rect 84671 266023 84699 266051
rect 84485 265961 84513 265989
rect 84547 265961 84575 265989
rect 84609 265961 84637 265989
rect 84671 265961 84699 265989
rect 91625 298578 91653 298606
rect 91687 298578 91715 298606
rect 91749 298578 91777 298606
rect 91811 298578 91839 298606
rect 91625 298516 91653 298544
rect 91687 298516 91715 298544
rect 91749 298516 91777 298544
rect 91811 298516 91839 298544
rect 91625 298454 91653 298482
rect 91687 298454 91715 298482
rect 91749 298454 91777 298482
rect 91811 298454 91839 298482
rect 91625 298392 91653 298420
rect 91687 298392 91715 298420
rect 91749 298392 91777 298420
rect 91811 298392 91839 298420
rect 91625 290147 91653 290175
rect 91687 290147 91715 290175
rect 91749 290147 91777 290175
rect 91811 290147 91839 290175
rect 91625 290085 91653 290113
rect 91687 290085 91715 290113
rect 91749 290085 91777 290113
rect 91811 290085 91839 290113
rect 91625 290023 91653 290051
rect 91687 290023 91715 290051
rect 91749 290023 91777 290051
rect 91811 290023 91839 290051
rect 91625 289961 91653 289989
rect 91687 289961 91715 289989
rect 91749 289961 91777 289989
rect 91811 289961 91839 289989
rect 91625 281147 91653 281175
rect 91687 281147 91715 281175
rect 91749 281147 91777 281175
rect 91811 281147 91839 281175
rect 91625 281085 91653 281113
rect 91687 281085 91715 281113
rect 91749 281085 91777 281113
rect 91811 281085 91839 281113
rect 91625 281023 91653 281051
rect 91687 281023 91715 281051
rect 91749 281023 91777 281051
rect 91811 281023 91839 281051
rect 91625 280961 91653 280989
rect 91687 280961 91715 280989
rect 91749 280961 91777 280989
rect 91811 280961 91839 280989
rect 91625 272147 91653 272175
rect 91687 272147 91715 272175
rect 91749 272147 91777 272175
rect 91811 272147 91839 272175
rect 91625 272085 91653 272113
rect 91687 272085 91715 272113
rect 91749 272085 91777 272113
rect 91811 272085 91839 272113
rect 91625 272023 91653 272051
rect 91687 272023 91715 272051
rect 91749 272023 91777 272051
rect 91811 272023 91839 272051
rect 91625 271961 91653 271989
rect 91687 271961 91715 271989
rect 91749 271961 91777 271989
rect 91811 271961 91839 271989
rect 91625 263147 91653 263175
rect 91687 263147 91715 263175
rect 91749 263147 91777 263175
rect 91811 263147 91839 263175
rect 91625 263085 91653 263113
rect 91687 263085 91715 263113
rect 91749 263085 91777 263113
rect 91811 263085 91839 263113
rect 91625 263023 91653 263051
rect 91687 263023 91715 263051
rect 91749 263023 91777 263051
rect 91811 263023 91839 263051
rect 91625 262961 91653 262989
rect 91687 262961 91715 262989
rect 91749 262961 91777 262989
rect 91811 262961 91839 262989
rect 93485 299058 93513 299086
rect 93547 299058 93575 299086
rect 93609 299058 93637 299086
rect 93671 299058 93699 299086
rect 93485 298996 93513 299024
rect 93547 298996 93575 299024
rect 93609 298996 93637 299024
rect 93671 298996 93699 299024
rect 93485 298934 93513 298962
rect 93547 298934 93575 298962
rect 93609 298934 93637 298962
rect 93671 298934 93699 298962
rect 93485 298872 93513 298900
rect 93547 298872 93575 298900
rect 93609 298872 93637 298900
rect 93671 298872 93699 298900
rect 93485 293147 93513 293175
rect 93547 293147 93575 293175
rect 93609 293147 93637 293175
rect 93671 293147 93699 293175
rect 93485 293085 93513 293113
rect 93547 293085 93575 293113
rect 93609 293085 93637 293113
rect 93671 293085 93699 293113
rect 93485 293023 93513 293051
rect 93547 293023 93575 293051
rect 93609 293023 93637 293051
rect 93671 293023 93699 293051
rect 93485 292961 93513 292989
rect 93547 292961 93575 292989
rect 93609 292961 93637 292989
rect 93671 292961 93699 292989
rect 93485 284147 93513 284175
rect 93547 284147 93575 284175
rect 93609 284147 93637 284175
rect 93671 284147 93699 284175
rect 93485 284085 93513 284113
rect 93547 284085 93575 284113
rect 93609 284085 93637 284113
rect 93671 284085 93699 284113
rect 93485 284023 93513 284051
rect 93547 284023 93575 284051
rect 93609 284023 93637 284051
rect 93671 284023 93699 284051
rect 93485 283961 93513 283989
rect 93547 283961 93575 283989
rect 93609 283961 93637 283989
rect 93671 283961 93699 283989
rect 93485 275147 93513 275175
rect 93547 275147 93575 275175
rect 93609 275147 93637 275175
rect 93671 275147 93699 275175
rect 93485 275085 93513 275113
rect 93547 275085 93575 275113
rect 93609 275085 93637 275113
rect 93671 275085 93699 275113
rect 93485 275023 93513 275051
rect 93547 275023 93575 275051
rect 93609 275023 93637 275051
rect 93671 275023 93699 275051
rect 93485 274961 93513 274989
rect 93547 274961 93575 274989
rect 93609 274961 93637 274989
rect 93671 274961 93699 274989
rect 93485 266147 93513 266175
rect 93547 266147 93575 266175
rect 93609 266147 93637 266175
rect 93671 266147 93699 266175
rect 93485 266085 93513 266113
rect 93547 266085 93575 266113
rect 93609 266085 93637 266113
rect 93671 266085 93699 266113
rect 93485 266023 93513 266051
rect 93547 266023 93575 266051
rect 93609 266023 93637 266051
rect 93671 266023 93699 266051
rect 93485 265961 93513 265989
rect 93547 265961 93575 265989
rect 93609 265961 93637 265989
rect 93671 265961 93699 265989
rect 100625 298578 100653 298606
rect 100687 298578 100715 298606
rect 100749 298578 100777 298606
rect 100811 298578 100839 298606
rect 100625 298516 100653 298544
rect 100687 298516 100715 298544
rect 100749 298516 100777 298544
rect 100811 298516 100839 298544
rect 100625 298454 100653 298482
rect 100687 298454 100715 298482
rect 100749 298454 100777 298482
rect 100811 298454 100839 298482
rect 100625 298392 100653 298420
rect 100687 298392 100715 298420
rect 100749 298392 100777 298420
rect 100811 298392 100839 298420
rect 100625 290147 100653 290175
rect 100687 290147 100715 290175
rect 100749 290147 100777 290175
rect 100811 290147 100839 290175
rect 100625 290085 100653 290113
rect 100687 290085 100715 290113
rect 100749 290085 100777 290113
rect 100811 290085 100839 290113
rect 100625 290023 100653 290051
rect 100687 290023 100715 290051
rect 100749 290023 100777 290051
rect 100811 290023 100839 290051
rect 100625 289961 100653 289989
rect 100687 289961 100715 289989
rect 100749 289961 100777 289989
rect 100811 289961 100839 289989
rect 100625 281147 100653 281175
rect 100687 281147 100715 281175
rect 100749 281147 100777 281175
rect 100811 281147 100839 281175
rect 100625 281085 100653 281113
rect 100687 281085 100715 281113
rect 100749 281085 100777 281113
rect 100811 281085 100839 281113
rect 100625 281023 100653 281051
rect 100687 281023 100715 281051
rect 100749 281023 100777 281051
rect 100811 281023 100839 281051
rect 100625 280961 100653 280989
rect 100687 280961 100715 280989
rect 100749 280961 100777 280989
rect 100811 280961 100839 280989
rect 100625 272147 100653 272175
rect 100687 272147 100715 272175
rect 100749 272147 100777 272175
rect 100811 272147 100839 272175
rect 100625 272085 100653 272113
rect 100687 272085 100715 272113
rect 100749 272085 100777 272113
rect 100811 272085 100839 272113
rect 100625 272023 100653 272051
rect 100687 272023 100715 272051
rect 100749 272023 100777 272051
rect 100811 272023 100839 272051
rect 100625 271961 100653 271989
rect 100687 271961 100715 271989
rect 100749 271961 100777 271989
rect 100811 271961 100839 271989
rect 100625 263147 100653 263175
rect 100687 263147 100715 263175
rect 100749 263147 100777 263175
rect 100811 263147 100839 263175
rect 100625 263085 100653 263113
rect 100687 263085 100715 263113
rect 100749 263085 100777 263113
rect 100811 263085 100839 263113
rect 100625 263023 100653 263051
rect 100687 263023 100715 263051
rect 100749 263023 100777 263051
rect 100811 263023 100839 263051
rect 100625 262961 100653 262989
rect 100687 262961 100715 262989
rect 100749 262961 100777 262989
rect 100811 262961 100839 262989
rect 102485 299058 102513 299086
rect 102547 299058 102575 299086
rect 102609 299058 102637 299086
rect 102671 299058 102699 299086
rect 102485 298996 102513 299024
rect 102547 298996 102575 299024
rect 102609 298996 102637 299024
rect 102671 298996 102699 299024
rect 102485 298934 102513 298962
rect 102547 298934 102575 298962
rect 102609 298934 102637 298962
rect 102671 298934 102699 298962
rect 102485 298872 102513 298900
rect 102547 298872 102575 298900
rect 102609 298872 102637 298900
rect 102671 298872 102699 298900
rect 102485 293147 102513 293175
rect 102547 293147 102575 293175
rect 102609 293147 102637 293175
rect 102671 293147 102699 293175
rect 102485 293085 102513 293113
rect 102547 293085 102575 293113
rect 102609 293085 102637 293113
rect 102671 293085 102699 293113
rect 102485 293023 102513 293051
rect 102547 293023 102575 293051
rect 102609 293023 102637 293051
rect 102671 293023 102699 293051
rect 102485 292961 102513 292989
rect 102547 292961 102575 292989
rect 102609 292961 102637 292989
rect 102671 292961 102699 292989
rect 102485 284147 102513 284175
rect 102547 284147 102575 284175
rect 102609 284147 102637 284175
rect 102671 284147 102699 284175
rect 102485 284085 102513 284113
rect 102547 284085 102575 284113
rect 102609 284085 102637 284113
rect 102671 284085 102699 284113
rect 102485 284023 102513 284051
rect 102547 284023 102575 284051
rect 102609 284023 102637 284051
rect 102671 284023 102699 284051
rect 102485 283961 102513 283989
rect 102547 283961 102575 283989
rect 102609 283961 102637 283989
rect 102671 283961 102699 283989
rect 102485 275147 102513 275175
rect 102547 275147 102575 275175
rect 102609 275147 102637 275175
rect 102671 275147 102699 275175
rect 102485 275085 102513 275113
rect 102547 275085 102575 275113
rect 102609 275085 102637 275113
rect 102671 275085 102699 275113
rect 102485 275023 102513 275051
rect 102547 275023 102575 275051
rect 102609 275023 102637 275051
rect 102671 275023 102699 275051
rect 102485 274961 102513 274989
rect 102547 274961 102575 274989
rect 102609 274961 102637 274989
rect 102671 274961 102699 274989
rect 102485 266147 102513 266175
rect 102547 266147 102575 266175
rect 102609 266147 102637 266175
rect 102671 266147 102699 266175
rect 102485 266085 102513 266113
rect 102547 266085 102575 266113
rect 102609 266085 102637 266113
rect 102671 266085 102699 266113
rect 102485 266023 102513 266051
rect 102547 266023 102575 266051
rect 102609 266023 102637 266051
rect 102671 266023 102699 266051
rect 102485 265961 102513 265989
rect 102547 265961 102575 265989
rect 102609 265961 102637 265989
rect 102671 265961 102699 265989
rect 109625 298578 109653 298606
rect 109687 298578 109715 298606
rect 109749 298578 109777 298606
rect 109811 298578 109839 298606
rect 109625 298516 109653 298544
rect 109687 298516 109715 298544
rect 109749 298516 109777 298544
rect 109811 298516 109839 298544
rect 109625 298454 109653 298482
rect 109687 298454 109715 298482
rect 109749 298454 109777 298482
rect 109811 298454 109839 298482
rect 109625 298392 109653 298420
rect 109687 298392 109715 298420
rect 109749 298392 109777 298420
rect 109811 298392 109839 298420
rect 109625 290147 109653 290175
rect 109687 290147 109715 290175
rect 109749 290147 109777 290175
rect 109811 290147 109839 290175
rect 109625 290085 109653 290113
rect 109687 290085 109715 290113
rect 109749 290085 109777 290113
rect 109811 290085 109839 290113
rect 109625 290023 109653 290051
rect 109687 290023 109715 290051
rect 109749 290023 109777 290051
rect 109811 290023 109839 290051
rect 109625 289961 109653 289989
rect 109687 289961 109715 289989
rect 109749 289961 109777 289989
rect 109811 289961 109839 289989
rect 109625 281147 109653 281175
rect 109687 281147 109715 281175
rect 109749 281147 109777 281175
rect 109811 281147 109839 281175
rect 109625 281085 109653 281113
rect 109687 281085 109715 281113
rect 109749 281085 109777 281113
rect 109811 281085 109839 281113
rect 109625 281023 109653 281051
rect 109687 281023 109715 281051
rect 109749 281023 109777 281051
rect 109811 281023 109839 281051
rect 109625 280961 109653 280989
rect 109687 280961 109715 280989
rect 109749 280961 109777 280989
rect 109811 280961 109839 280989
rect 109625 272147 109653 272175
rect 109687 272147 109715 272175
rect 109749 272147 109777 272175
rect 109811 272147 109839 272175
rect 109625 272085 109653 272113
rect 109687 272085 109715 272113
rect 109749 272085 109777 272113
rect 109811 272085 109839 272113
rect 109625 272023 109653 272051
rect 109687 272023 109715 272051
rect 109749 272023 109777 272051
rect 109811 272023 109839 272051
rect 109625 271961 109653 271989
rect 109687 271961 109715 271989
rect 109749 271961 109777 271989
rect 109811 271961 109839 271989
rect 109625 263147 109653 263175
rect 109687 263147 109715 263175
rect 109749 263147 109777 263175
rect 109811 263147 109839 263175
rect 109625 263085 109653 263113
rect 109687 263085 109715 263113
rect 109749 263085 109777 263113
rect 109811 263085 109839 263113
rect 109625 263023 109653 263051
rect 109687 263023 109715 263051
rect 109749 263023 109777 263051
rect 109811 263023 109839 263051
rect 109625 262961 109653 262989
rect 109687 262961 109715 262989
rect 109749 262961 109777 262989
rect 109811 262961 109839 262989
rect 111485 299058 111513 299086
rect 111547 299058 111575 299086
rect 111609 299058 111637 299086
rect 111671 299058 111699 299086
rect 111485 298996 111513 299024
rect 111547 298996 111575 299024
rect 111609 298996 111637 299024
rect 111671 298996 111699 299024
rect 111485 298934 111513 298962
rect 111547 298934 111575 298962
rect 111609 298934 111637 298962
rect 111671 298934 111699 298962
rect 111485 298872 111513 298900
rect 111547 298872 111575 298900
rect 111609 298872 111637 298900
rect 111671 298872 111699 298900
rect 111485 293147 111513 293175
rect 111547 293147 111575 293175
rect 111609 293147 111637 293175
rect 111671 293147 111699 293175
rect 111485 293085 111513 293113
rect 111547 293085 111575 293113
rect 111609 293085 111637 293113
rect 111671 293085 111699 293113
rect 111485 293023 111513 293051
rect 111547 293023 111575 293051
rect 111609 293023 111637 293051
rect 111671 293023 111699 293051
rect 111485 292961 111513 292989
rect 111547 292961 111575 292989
rect 111609 292961 111637 292989
rect 111671 292961 111699 292989
rect 111485 284147 111513 284175
rect 111547 284147 111575 284175
rect 111609 284147 111637 284175
rect 111671 284147 111699 284175
rect 111485 284085 111513 284113
rect 111547 284085 111575 284113
rect 111609 284085 111637 284113
rect 111671 284085 111699 284113
rect 111485 284023 111513 284051
rect 111547 284023 111575 284051
rect 111609 284023 111637 284051
rect 111671 284023 111699 284051
rect 111485 283961 111513 283989
rect 111547 283961 111575 283989
rect 111609 283961 111637 283989
rect 111671 283961 111699 283989
rect 111485 275147 111513 275175
rect 111547 275147 111575 275175
rect 111609 275147 111637 275175
rect 111671 275147 111699 275175
rect 111485 275085 111513 275113
rect 111547 275085 111575 275113
rect 111609 275085 111637 275113
rect 111671 275085 111699 275113
rect 111485 275023 111513 275051
rect 111547 275023 111575 275051
rect 111609 275023 111637 275051
rect 111671 275023 111699 275051
rect 111485 274961 111513 274989
rect 111547 274961 111575 274989
rect 111609 274961 111637 274989
rect 111671 274961 111699 274989
rect 111485 266147 111513 266175
rect 111547 266147 111575 266175
rect 111609 266147 111637 266175
rect 111671 266147 111699 266175
rect 111485 266085 111513 266113
rect 111547 266085 111575 266113
rect 111609 266085 111637 266113
rect 111671 266085 111699 266113
rect 111485 266023 111513 266051
rect 111547 266023 111575 266051
rect 111609 266023 111637 266051
rect 111671 266023 111699 266051
rect 111485 265961 111513 265989
rect 111547 265961 111575 265989
rect 111609 265961 111637 265989
rect 111671 265961 111699 265989
rect 118625 298578 118653 298606
rect 118687 298578 118715 298606
rect 118749 298578 118777 298606
rect 118811 298578 118839 298606
rect 118625 298516 118653 298544
rect 118687 298516 118715 298544
rect 118749 298516 118777 298544
rect 118811 298516 118839 298544
rect 118625 298454 118653 298482
rect 118687 298454 118715 298482
rect 118749 298454 118777 298482
rect 118811 298454 118839 298482
rect 118625 298392 118653 298420
rect 118687 298392 118715 298420
rect 118749 298392 118777 298420
rect 118811 298392 118839 298420
rect 118625 290147 118653 290175
rect 118687 290147 118715 290175
rect 118749 290147 118777 290175
rect 118811 290147 118839 290175
rect 118625 290085 118653 290113
rect 118687 290085 118715 290113
rect 118749 290085 118777 290113
rect 118811 290085 118839 290113
rect 118625 290023 118653 290051
rect 118687 290023 118715 290051
rect 118749 290023 118777 290051
rect 118811 290023 118839 290051
rect 118625 289961 118653 289989
rect 118687 289961 118715 289989
rect 118749 289961 118777 289989
rect 118811 289961 118839 289989
rect 118625 281147 118653 281175
rect 118687 281147 118715 281175
rect 118749 281147 118777 281175
rect 118811 281147 118839 281175
rect 118625 281085 118653 281113
rect 118687 281085 118715 281113
rect 118749 281085 118777 281113
rect 118811 281085 118839 281113
rect 118625 281023 118653 281051
rect 118687 281023 118715 281051
rect 118749 281023 118777 281051
rect 118811 281023 118839 281051
rect 118625 280961 118653 280989
rect 118687 280961 118715 280989
rect 118749 280961 118777 280989
rect 118811 280961 118839 280989
rect 118625 272147 118653 272175
rect 118687 272147 118715 272175
rect 118749 272147 118777 272175
rect 118811 272147 118839 272175
rect 118625 272085 118653 272113
rect 118687 272085 118715 272113
rect 118749 272085 118777 272113
rect 118811 272085 118839 272113
rect 118625 272023 118653 272051
rect 118687 272023 118715 272051
rect 118749 272023 118777 272051
rect 118811 272023 118839 272051
rect 118625 271961 118653 271989
rect 118687 271961 118715 271989
rect 118749 271961 118777 271989
rect 118811 271961 118839 271989
rect 118625 263147 118653 263175
rect 118687 263147 118715 263175
rect 118749 263147 118777 263175
rect 118811 263147 118839 263175
rect 118625 263085 118653 263113
rect 118687 263085 118715 263113
rect 118749 263085 118777 263113
rect 118811 263085 118839 263113
rect 118625 263023 118653 263051
rect 118687 263023 118715 263051
rect 118749 263023 118777 263051
rect 118811 263023 118839 263051
rect 118625 262961 118653 262989
rect 118687 262961 118715 262989
rect 118749 262961 118777 262989
rect 118811 262961 118839 262989
rect 120485 299058 120513 299086
rect 120547 299058 120575 299086
rect 120609 299058 120637 299086
rect 120671 299058 120699 299086
rect 120485 298996 120513 299024
rect 120547 298996 120575 299024
rect 120609 298996 120637 299024
rect 120671 298996 120699 299024
rect 120485 298934 120513 298962
rect 120547 298934 120575 298962
rect 120609 298934 120637 298962
rect 120671 298934 120699 298962
rect 120485 298872 120513 298900
rect 120547 298872 120575 298900
rect 120609 298872 120637 298900
rect 120671 298872 120699 298900
rect 120485 293147 120513 293175
rect 120547 293147 120575 293175
rect 120609 293147 120637 293175
rect 120671 293147 120699 293175
rect 120485 293085 120513 293113
rect 120547 293085 120575 293113
rect 120609 293085 120637 293113
rect 120671 293085 120699 293113
rect 120485 293023 120513 293051
rect 120547 293023 120575 293051
rect 120609 293023 120637 293051
rect 120671 293023 120699 293051
rect 120485 292961 120513 292989
rect 120547 292961 120575 292989
rect 120609 292961 120637 292989
rect 120671 292961 120699 292989
rect 120485 284147 120513 284175
rect 120547 284147 120575 284175
rect 120609 284147 120637 284175
rect 120671 284147 120699 284175
rect 120485 284085 120513 284113
rect 120547 284085 120575 284113
rect 120609 284085 120637 284113
rect 120671 284085 120699 284113
rect 120485 284023 120513 284051
rect 120547 284023 120575 284051
rect 120609 284023 120637 284051
rect 120671 284023 120699 284051
rect 120485 283961 120513 283989
rect 120547 283961 120575 283989
rect 120609 283961 120637 283989
rect 120671 283961 120699 283989
rect 120485 275147 120513 275175
rect 120547 275147 120575 275175
rect 120609 275147 120637 275175
rect 120671 275147 120699 275175
rect 120485 275085 120513 275113
rect 120547 275085 120575 275113
rect 120609 275085 120637 275113
rect 120671 275085 120699 275113
rect 120485 275023 120513 275051
rect 120547 275023 120575 275051
rect 120609 275023 120637 275051
rect 120671 275023 120699 275051
rect 120485 274961 120513 274989
rect 120547 274961 120575 274989
rect 120609 274961 120637 274989
rect 120671 274961 120699 274989
rect 120485 266147 120513 266175
rect 120547 266147 120575 266175
rect 120609 266147 120637 266175
rect 120671 266147 120699 266175
rect 120485 266085 120513 266113
rect 120547 266085 120575 266113
rect 120609 266085 120637 266113
rect 120671 266085 120699 266113
rect 120485 266023 120513 266051
rect 120547 266023 120575 266051
rect 120609 266023 120637 266051
rect 120671 266023 120699 266051
rect 120485 265961 120513 265989
rect 120547 265961 120575 265989
rect 120609 265961 120637 265989
rect 120671 265961 120699 265989
rect 127625 298578 127653 298606
rect 127687 298578 127715 298606
rect 127749 298578 127777 298606
rect 127811 298578 127839 298606
rect 127625 298516 127653 298544
rect 127687 298516 127715 298544
rect 127749 298516 127777 298544
rect 127811 298516 127839 298544
rect 127625 298454 127653 298482
rect 127687 298454 127715 298482
rect 127749 298454 127777 298482
rect 127811 298454 127839 298482
rect 127625 298392 127653 298420
rect 127687 298392 127715 298420
rect 127749 298392 127777 298420
rect 127811 298392 127839 298420
rect 127625 290147 127653 290175
rect 127687 290147 127715 290175
rect 127749 290147 127777 290175
rect 127811 290147 127839 290175
rect 127625 290085 127653 290113
rect 127687 290085 127715 290113
rect 127749 290085 127777 290113
rect 127811 290085 127839 290113
rect 127625 290023 127653 290051
rect 127687 290023 127715 290051
rect 127749 290023 127777 290051
rect 127811 290023 127839 290051
rect 127625 289961 127653 289989
rect 127687 289961 127715 289989
rect 127749 289961 127777 289989
rect 127811 289961 127839 289989
rect 127625 281147 127653 281175
rect 127687 281147 127715 281175
rect 127749 281147 127777 281175
rect 127811 281147 127839 281175
rect 127625 281085 127653 281113
rect 127687 281085 127715 281113
rect 127749 281085 127777 281113
rect 127811 281085 127839 281113
rect 127625 281023 127653 281051
rect 127687 281023 127715 281051
rect 127749 281023 127777 281051
rect 127811 281023 127839 281051
rect 127625 280961 127653 280989
rect 127687 280961 127715 280989
rect 127749 280961 127777 280989
rect 127811 280961 127839 280989
rect 127625 272147 127653 272175
rect 127687 272147 127715 272175
rect 127749 272147 127777 272175
rect 127811 272147 127839 272175
rect 127625 272085 127653 272113
rect 127687 272085 127715 272113
rect 127749 272085 127777 272113
rect 127811 272085 127839 272113
rect 127625 272023 127653 272051
rect 127687 272023 127715 272051
rect 127749 272023 127777 272051
rect 127811 272023 127839 272051
rect 127625 271961 127653 271989
rect 127687 271961 127715 271989
rect 127749 271961 127777 271989
rect 127811 271961 127839 271989
rect 127625 263147 127653 263175
rect 127687 263147 127715 263175
rect 127749 263147 127777 263175
rect 127811 263147 127839 263175
rect 127625 263085 127653 263113
rect 127687 263085 127715 263113
rect 127749 263085 127777 263113
rect 127811 263085 127839 263113
rect 127625 263023 127653 263051
rect 127687 263023 127715 263051
rect 127749 263023 127777 263051
rect 127811 263023 127839 263051
rect 127625 262961 127653 262989
rect 127687 262961 127715 262989
rect 127749 262961 127777 262989
rect 127811 262961 127839 262989
rect 129485 299058 129513 299086
rect 129547 299058 129575 299086
rect 129609 299058 129637 299086
rect 129671 299058 129699 299086
rect 129485 298996 129513 299024
rect 129547 298996 129575 299024
rect 129609 298996 129637 299024
rect 129671 298996 129699 299024
rect 129485 298934 129513 298962
rect 129547 298934 129575 298962
rect 129609 298934 129637 298962
rect 129671 298934 129699 298962
rect 129485 298872 129513 298900
rect 129547 298872 129575 298900
rect 129609 298872 129637 298900
rect 129671 298872 129699 298900
rect 129485 293147 129513 293175
rect 129547 293147 129575 293175
rect 129609 293147 129637 293175
rect 129671 293147 129699 293175
rect 129485 293085 129513 293113
rect 129547 293085 129575 293113
rect 129609 293085 129637 293113
rect 129671 293085 129699 293113
rect 129485 293023 129513 293051
rect 129547 293023 129575 293051
rect 129609 293023 129637 293051
rect 129671 293023 129699 293051
rect 129485 292961 129513 292989
rect 129547 292961 129575 292989
rect 129609 292961 129637 292989
rect 129671 292961 129699 292989
rect 129485 284147 129513 284175
rect 129547 284147 129575 284175
rect 129609 284147 129637 284175
rect 129671 284147 129699 284175
rect 129485 284085 129513 284113
rect 129547 284085 129575 284113
rect 129609 284085 129637 284113
rect 129671 284085 129699 284113
rect 129485 284023 129513 284051
rect 129547 284023 129575 284051
rect 129609 284023 129637 284051
rect 129671 284023 129699 284051
rect 129485 283961 129513 283989
rect 129547 283961 129575 283989
rect 129609 283961 129637 283989
rect 129671 283961 129699 283989
rect 129485 275147 129513 275175
rect 129547 275147 129575 275175
rect 129609 275147 129637 275175
rect 129671 275147 129699 275175
rect 129485 275085 129513 275113
rect 129547 275085 129575 275113
rect 129609 275085 129637 275113
rect 129671 275085 129699 275113
rect 129485 275023 129513 275051
rect 129547 275023 129575 275051
rect 129609 275023 129637 275051
rect 129671 275023 129699 275051
rect 129485 274961 129513 274989
rect 129547 274961 129575 274989
rect 129609 274961 129637 274989
rect 129671 274961 129699 274989
rect 129485 266147 129513 266175
rect 129547 266147 129575 266175
rect 129609 266147 129637 266175
rect 129671 266147 129699 266175
rect 129485 266085 129513 266113
rect 129547 266085 129575 266113
rect 129609 266085 129637 266113
rect 129671 266085 129699 266113
rect 129485 266023 129513 266051
rect 129547 266023 129575 266051
rect 129609 266023 129637 266051
rect 129671 266023 129699 266051
rect 129485 265961 129513 265989
rect 129547 265961 129575 265989
rect 129609 265961 129637 265989
rect 129671 265961 129699 265989
rect 136625 298578 136653 298606
rect 136687 298578 136715 298606
rect 136749 298578 136777 298606
rect 136811 298578 136839 298606
rect 136625 298516 136653 298544
rect 136687 298516 136715 298544
rect 136749 298516 136777 298544
rect 136811 298516 136839 298544
rect 136625 298454 136653 298482
rect 136687 298454 136715 298482
rect 136749 298454 136777 298482
rect 136811 298454 136839 298482
rect 136625 298392 136653 298420
rect 136687 298392 136715 298420
rect 136749 298392 136777 298420
rect 136811 298392 136839 298420
rect 136625 290147 136653 290175
rect 136687 290147 136715 290175
rect 136749 290147 136777 290175
rect 136811 290147 136839 290175
rect 136625 290085 136653 290113
rect 136687 290085 136715 290113
rect 136749 290085 136777 290113
rect 136811 290085 136839 290113
rect 136625 290023 136653 290051
rect 136687 290023 136715 290051
rect 136749 290023 136777 290051
rect 136811 290023 136839 290051
rect 136625 289961 136653 289989
rect 136687 289961 136715 289989
rect 136749 289961 136777 289989
rect 136811 289961 136839 289989
rect 136625 281147 136653 281175
rect 136687 281147 136715 281175
rect 136749 281147 136777 281175
rect 136811 281147 136839 281175
rect 136625 281085 136653 281113
rect 136687 281085 136715 281113
rect 136749 281085 136777 281113
rect 136811 281085 136839 281113
rect 136625 281023 136653 281051
rect 136687 281023 136715 281051
rect 136749 281023 136777 281051
rect 136811 281023 136839 281051
rect 136625 280961 136653 280989
rect 136687 280961 136715 280989
rect 136749 280961 136777 280989
rect 136811 280961 136839 280989
rect 136625 272147 136653 272175
rect 136687 272147 136715 272175
rect 136749 272147 136777 272175
rect 136811 272147 136839 272175
rect 136625 272085 136653 272113
rect 136687 272085 136715 272113
rect 136749 272085 136777 272113
rect 136811 272085 136839 272113
rect 136625 272023 136653 272051
rect 136687 272023 136715 272051
rect 136749 272023 136777 272051
rect 136811 272023 136839 272051
rect 136625 271961 136653 271989
rect 136687 271961 136715 271989
rect 136749 271961 136777 271989
rect 136811 271961 136839 271989
rect 136625 263147 136653 263175
rect 136687 263147 136715 263175
rect 136749 263147 136777 263175
rect 136811 263147 136839 263175
rect 136625 263085 136653 263113
rect 136687 263085 136715 263113
rect 136749 263085 136777 263113
rect 136811 263085 136839 263113
rect 136625 263023 136653 263051
rect 136687 263023 136715 263051
rect 136749 263023 136777 263051
rect 136811 263023 136839 263051
rect 136625 262961 136653 262989
rect 136687 262961 136715 262989
rect 136749 262961 136777 262989
rect 136811 262961 136839 262989
rect 138485 299058 138513 299086
rect 138547 299058 138575 299086
rect 138609 299058 138637 299086
rect 138671 299058 138699 299086
rect 138485 298996 138513 299024
rect 138547 298996 138575 299024
rect 138609 298996 138637 299024
rect 138671 298996 138699 299024
rect 138485 298934 138513 298962
rect 138547 298934 138575 298962
rect 138609 298934 138637 298962
rect 138671 298934 138699 298962
rect 138485 298872 138513 298900
rect 138547 298872 138575 298900
rect 138609 298872 138637 298900
rect 138671 298872 138699 298900
rect 138485 293147 138513 293175
rect 138547 293147 138575 293175
rect 138609 293147 138637 293175
rect 138671 293147 138699 293175
rect 138485 293085 138513 293113
rect 138547 293085 138575 293113
rect 138609 293085 138637 293113
rect 138671 293085 138699 293113
rect 138485 293023 138513 293051
rect 138547 293023 138575 293051
rect 138609 293023 138637 293051
rect 138671 293023 138699 293051
rect 138485 292961 138513 292989
rect 138547 292961 138575 292989
rect 138609 292961 138637 292989
rect 138671 292961 138699 292989
rect 138485 284147 138513 284175
rect 138547 284147 138575 284175
rect 138609 284147 138637 284175
rect 138671 284147 138699 284175
rect 138485 284085 138513 284113
rect 138547 284085 138575 284113
rect 138609 284085 138637 284113
rect 138671 284085 138699 284113
rect 138485 284023 138513 284051
rect 138547 284023 138575 284051
rect 138609 284023 138637 284051
rect 138671 284023 138699 284051
rect 138485 283961 138513 283989
rect 138547 283961 138575 283989
rect 138609 283961 138637 283989
rect 138671 283961 138699 283989
rect 138485 275147 138513 275175
rect 138547 275147 138575 275175
rect 138609 275147 138637 275175
rect 138671 275147 138699 275175
rect 138485 275085 138513 275113
rect 138547 275085 138575 275113
rect 138609 275085 138637 275113
rect 138671 275085 138699 275113
rect 138485 275023 138513 275051
rect 138547 275023 138575 275051
rect 138609 275023 138637 275051
rect 138671 275023 138699 275051
rect 138485 274961 138513 274989
rect 138547 274961 138575 274989
rect 138609 274961 138637 274989
rect 138671 274961 138699 274989
rect 138485 266147 138513 266175
rect 138547 266147 138575 266175
rect 138609 266147 138637 266175
rect 138671 266147 138699 266175
rect 138485 266085 138513 266113
rect 138547 266085 138575 266113
rect 138609 266085 138637 266113
rect 138671 266085 138699 266113
rect 138485 266023 138513 266051
rect 138547 266023 138575 266051
rect 138609 266023 138637 266051
rect 138671 266023 138699 266051
rect 138485 265961 138513 265989
rect 138547 265961 138575 265989
rect 138609 265961 138637 265989
rect 138671 265961 138699 265989
rect 145625 298578 145653 298606
rect 145687 298578 145715 298606
rect 145749 298578 145777 298606
rect 145811 298578 145839 298606
rect 145625 298516 145653 298544
rect 145687 298516 145715 298544
rect 145749 298516 145777 298544
rect 145811 298516 145839 298544
rect 145625 298454 145653 298482
rect 145687 298454 145715 298482
rect 145749 298454 145777 298482
rect 145811 298454 145839 298482
rect 145625 298392 145653 298420
rect 145687 298392 145715 298420
rect 145749 298392 145777 298420
rect 145811 298392 145839 298420
rect 145625 290147 145653 290175
rect 145687 290147 145715 290175
rect 145749 290147 145777 290175
rect 145811 290147 145839 290175
rect 145625 290085 145653 290113
rect 145687 290085 145715 290113
rect 145749 290085 145777 290113
rect 145811 290085 145839 290113
rect 145625 290023 145653 290051
rect 145687 290023 145715 290051
rect 145749 290023 145777 290051
rect 145811 290023 145839 290051
rect 145625 289961 145653 289989
rect 145687 289961 145715 289989
rect 145749 289961 145777 289989
rect 145811 289961 145839 289989
rect 145625 281147 145653 281175
rect 145687 281147 145715 281175
rect 145749 281147 145777 281175
rect 145811 281147 145839 281175
rect 145625 281085 145653 281113
rect 145687 281085 145715 281113
rect 145749 281085 145777 281113
rect 145811 281085 145839 281113
rect 145625 281023 145653 281051
rect 145687 281023 145715 281051
rect 145749 281023 145777 281051
rect 145811 281023 145839 281051
rect 145625 280961 145653 280989
rect 145687 280961 145715 280989
rect 145749 280961 145777 280989
rect 145811 280961 145839 280989
rect 145625 272147 145653 272175
rect 145687 272147 145715 272175
rect 145749 272147 145777 272175
rect 145811 272147 145839 272175
rect 145625 272085 145653 272113
rect 145687 272085 145715 272113
rect 145749 272085 145777 272113
rect 145811 272085 145839 272113
rect 145625 272023 145653 272051
rect 145687 272023 145715 272051
rect 145749 272023 145777 272051
rect 145811 272023 145839 272051
rect 145625 271961 145653 271989
rect 145687 271961 145715 271989
rect 145749 271961 145777 271989
rect 145811 271961 145839 271989
rect 145625 263147 145653 263175
rect 145687 263147 145715 263175
rect 145749 263147 145777 263175
rect 145811 263147 145839 263175
rect 145625 263085 145653 263113
rect 145687 263085 145715 263113
rect 145749 263085 145777 263113
rect 145811 263085 145839 263113
rect 145625 263023 145653 263051
rect 145687 263023 145715 263051
rect 145749 263023 145777 263051
rect 145811 263023 145839 263051
rect 145625 262961 145653 262989
rect 145687 262961 145715 262989
rect 145749 262961 145777 262989
rect 145811 262961 145839 262989
rect 147485 299058 147513 299086
rect 147547 299058 147575 299086
rect 147609 299058 147637 299086
rect 147671 299058 147699 299086
rect 147485 298996 147513 299024
rect 147547 298996 147575 299024
rect 147609 298996 147637 299024
rect 147671 298996 147699 299024
rect 147485 298934 147513 298962
rect 147547 298934 147575 298962
rect 147609 298934 147637 298962
rect 147671 298934 147699 298962
rect 147485 298872 147513 298900
rect 147547 298872 147575 298900
rect 147609 298872 147637 298900
rect 147671 298872 147699 298900
rect 147485 293147 147513 293175
rect 147547 293147 147575 293175
rect 147609 293147 147637 293175
rect 147671 293147 147699 293175
rect 147485 293085 147513 293113
rect 147547 293085 147575 293113
rect 147609 293085 147637 293113
rect 147671 293085 147699 293113
rect 147485 293023 147513 293051
rect 147547 293023 147575 293051
rect 147609 293023 147637 293051
rect 147671 293023 147699 293051
rect 147485 292961 147513 292989
rect 147547 292961 147575 292989
rect 147609 292961 147637 292989
rect 147671 292961 147699 292989
rect 147485 284147 147513 284175
rect 147547 284147 147575 284175
rect 147609 284147 147637 284175
rect 147671 284147 147699 284175
rect 147485 284085 147513 284113
rect 147547 284085 147575 284113
rect 147609 284085 147637 284113
rect 147671 284085 147699 284113
rect 147485 284023 147513 284051
rect 147547 284023 147575 284051
rect 147609 284023 147637 284051
rect 147671 284023 147699 284051
rect 147485 283961 147513 283989
rect 147547 283961 147575 283989
rect 147609 283961 147637 283989
rect 147671 283961 147699 283989
rect 147485 275147 147513 275175
rect 147547 275147 147575 275175
rect 147609 275147 147637 275175
rect 147671 275147 147699 275175
rect 147485 275085 147513 275113
rect 147547 275085 147575 275113
rect 147609 275085 147637 275113
rect 147671 275085 147699 275113
rect 147485 275023 147513 275051
rect 147547 275023 147575 275051
rect 147609 275023 147637 275051
rect 147671 275023 147699 275051
rect 147485 274961 147513 274989
rect 147547 274961 147575 274989
rect 147609 274961 147637 274989
rect 147671 274961 147699 274989
rect 147485 266147 147513 266175
rect 147547 266147 147575 266175
rect 147609 266147 147637 266175
rect 147671 266147 147699 266175
rect 147485 266085 147513 266113
rect 147547 266085 147575 266113
rect 147609 266085 147637 266113
rect 147671 266085 147699 266113
rect 147485 266023 147513 266051
rect 147547 266023 147575 266051
rect 147609 266023 147637 266051
rect 147671 266023 147699 266051
rect 147485 265961 147513 265989
rect 147547 265961 147575 265989
rect 147609 265961 147637 265989
rect 147671 265961 147699 265989
rect 154625 298578 154653 298606
rect 154687 298578 154715 298606
rect 154749 298578 154777 298606
rect 154811 298578 154839 298606
rect 154625 298516 154653 298544
rect 154687 298516 154715 298544
rect 154749 298516 154777 298544
rect 154811 298516 154839 298544
rect 154625 298454 154653 298482
rect 154687 298454 154715 298482
rect 154749 298454 154777 298482
rect 154811 298454 154839 298482
rect 154625 298392 154653 298420
rect 154687 298392 154715 298420
rect 154749 298392 154777 298420
rect 154811 298392 154839 298420
rect 154625 290147 154653 290175
rect 154687 290147 154715 290175
rect 154749 290147 154777 290175
rect 154811 290147 154839 290175
rect 154625 290085 154653 290113
rect 154687 290085 154715 290113
rect 154749 290085 154777 290113
rect 154811 290085 154839 290113
rect 154625 290023 154653 290051
rect 154687 290023 154715 290051
rect 154749 290023 154777 290051
rect 154811 290023 154839 290051
rect 154625 289961 154653 289989
rect 154687 289961 154715 289989
rect 154749 289961 154777 289989
rect 154811 289961 154839 289989
rect 154625 281147 154653 281175
rect 154687 281147 154715 281175
rect 154749 281147 154777 281175
rect 154811 281147 154839 281175
rect 154625 281085 154653 281113
rect 154687 281085 154715 281113
rect 154749 281085 154777 281113
rect 154811 281085 154839 281113
rect 154625 281023 154653 281051
rect 154687 281023 154715 281051
rect 154749 281023 154777 281051
rect 154811 281023 154839 281051
rect 154625 280961 154653 280989
rect 154687 280961 154715 280989
rect 154749 280961 154777 280989
rect 154811 280961 154839 280989
rect 154625 272147 154653 272175
rect 154687 272147 154715 272175
rect 154749 272147 154777 272175
rect 154811 272147 154839 272175
rect 154625 272085 154653 272113
rect 154687 272085 154715 272113
rect 154749 272085 154777 272113
rect 154811 272085 154839 272113
rect 154625 272023 154653 272051
rect 154687 272023 154715 272051
rect 154749 272023 154777 272051
rect 154811 272023 154839 272051
rect 154625 271961 154653 271989
rect 154687 271961 154715 271989
rect 154749 271961 154777 271989
rect 154811 271961 154839 271989
rect 154625 263147 154653 263175
rect 154687 263147 154715 263175
rect 154749 263147 154777 263175
rect 154811 263147 154839 263175
rect 154625 263085 154653 263113
rect 154687 263085 154715 263113
rect 154749 263085 154777 263113
rect 154811 263085 154839 263113
rect 154625 263023 154653 263051
rect 154687 263023 154715 263051
rect 154749 263023 154777 263051
rect 154811 263023 154839 263051
rect 154625 262961 154653 262989
rect 154687 262961 154715 262989
rect 154749 262961 154777 262989
rect 154811 262961 154839 262989
rect 48485 257147 48513 257175
rect 48547 257147 48575 257175
rect 48609 257147 48637 257175
rect 48671 257147 48699 257175
rect 48485 257085 48513 257113
rect 48547 257085 48575 257113
rect 48609 257085 48637 257113
rect 48671 257085 48699 257113
rect 48485 257023 48513 257051
rect 48547 257023 48575 257051
rect 48609 257023 48637 257051
rect 48671 257023 48699 257051
rect 48485 256961 48513 256989
rect 48547 256961 48575 256989
rect 48609 256961 48637 256989
rect 48671 256961 48699 256989
rect 59939 257147 59967 257175
rect 60001 257147 60029 257175
rect 59939 257085 59967 257113
rect 60001 257085 60029 257113
rect 59939 257023 59967 257051
rect 60001 257023 60029 257051
rect 59939 256961 59967 256989
rect 60001 256961 60029 256989
rect 75299 257147 75327 257175
rect 75361 257147 75389 257175
rect 75299 257085 75327 257113
rect 75361 257085 75389 257113
rect 75299 257023 75327 257051
rect 75361 257023 75389 257051
rect 75299 256961 75327 256989
rect 75361 256961 75389 256989
rect 90659 257147 90687 257175
rect 90721 257147 90749 257175
rect 90659 257085 90687 257113
rect 90721 257085 90749 257113
rect 90659 257023 90687 257051
rect 90721 257023 90749 257051
rect 90659 256961 90687 256989
rect 90721 256961 90749 256989
rect 106019 257147 106047 257175
rect 106081 257147 106109 257175
rect 106019 257085 106047 257113
rect 106081 257085 106109 257113
rect 106019 257023 106047 257051
rect 106081 257023 106109 257051
rect 106019 256961 106047 256989
rect 106081 256961 106109 256989
rect 121379 257147 121407 257175
rect 121441 257147 121469 257175
rect 121379 257085 121407 257113
rect 121441 257085 121469 257113
rect 121379 257023 121407 257051
rect 121441 257023 121469 257051
rect 121379 256961 121407 256989
rect 121441 256961 121469 256989
rect 136739 257147 136767 257175
rect 136801 257147 136829 257175
rect 136739 257085 136767 257113
rect 136801 257085 136829 257113
rect 136739 257023 136767 257051
rect 136801 257023 136829 257051
rect 136739 256961 136767 256989
rect 136801 256961 136829 256989
rect 52259 254147 52287 254175
rect 52321 254147 52349 254175
rect 52259 254085 52287 254113
rect 52321 254085 52349 254113
rect 52259 254023 52287 254051
rect 52321 254023 52349 254051
rect 52259 253961 52287 253989
rect 52321 253961 52349 253989
rect 67619 254147 67647 254175
rect 67681 254147 67709 254175
rect 67619 254085 67647 254113
rect 67681 254085 67709 254113
rect 67619 254023 67647 254051
rect 67681 254023 67709 254051
rect 67619 253961 67647 253989
rect 67681 253961 67709 253989
rect 82979 254147 83007 254175
rect 83041 254147 83069 254175
rect 82979 254085 83007 254113
rect 83041 254085 83069 254113
rect 82979 254023 83007 254051
rect 83041 254023 83069 254051
rect 82979 253961 83007 253989
rect 83041 253961 83069 253989
rect 98339 254147 98367 254175
rect 98401 254147 98429 254175
rect 98339 254085 98367 254113
rect 98401 254085 98429 254113
rect 98339 254023 98367 254051
rect 98401 254023 98429 254051
rect 98339 253961 98367 253989
rect 98401 253961 98429 253989
rect 113699 254147 113727 254175
rect 113761 254147 113789 254175
rect 113699 254085 113727 254113
rect 113761 254085 113789 254113
rect 113699 254023 113727 254051
rect 113761 254023 113789 254051
rect 113699 253961 113727 253989
rect 113761 253961 113789 253989
rect 129059 254147 129087 254175
rect 129121 254147 129149 254175
rect 129059 254085 129087 254113
rect 129121 254085 129149 254113
rect 129059 254023 129087 254051
rect 129121 254023 129149 254051
rect 129059 253961 129087 253989
rect 129121 253961 129149 253989
rect 144419 254147 144447 254175
rect 144481 254147 144509 254175
rect 144419 254085 144447 254113
rect 144481 254085 144509 254113
rect 144419 254023 144447 254051
rect 144481 254023 144509 254051
rect 144419 253961 144447 253989
rect 144481 253961 144509 253989
rect 154625 254147 154653 254175
rect 154687 254147 154715 254175
rect 154749 254147 154777 254175
rect 154811 254147 154839 254175
rect 154625 254085 154653 254113
rect 154687 254085 154715 254113
rect 154749 254085 154777 254113
rect 154811 254085 154839 254113
rect 154625 254023 154653 254051
rect 154687 254023 154715 254051
rect 154749 254023 154777 254051
rect 154811 254023 154839 254051
rect 154625 253961 154653 253989
rect 154687 253961 154715 253989
rect 154749 253961 154777 253989
rect 154811 253961 154839 253989
rect 48485 248147 48513 248175
rect 48547 248147 48575 248175
rect 48609 248147 48637 248175
rect 48671 248147 48699 248175
rect 48485 248085 48513 248113
rect 48547 248085 48575 248113
rect 48609 248085 48637 248113
rect 48671 248085 48699 248113
rect 48485 248023 48513 248051
rect 48547 248023 48575 248051
rect 48609 248023 48637 248051
rect 48671 248023 48699 248051
rect 48485 247961 48513 247989
rect 48547 247961 48575 247989
rect 48609 247961 48637 247989
rect 48671 247961 48699 247989
rect 59939 248147 59967 248175
rect 60001 248147 60029 248175
rect 59939 248085 59967 248113
rect 60001 248085 60029 248113
rect 59939 248023 59967 248051
rect 60001 248023 60029 248051
rect 59939 247961 59967 247989
rect 60001 247961 60029 247989
rect 75299 248147 75327 248175
rect 75361 248147 75389 248175
rect 75299 248085 75327 248113
rect 75361 248085 75389 248113
rect 75299 248023 75327 248051
rect 75361 248023 75389 248051
rect 75299 247961 75327 247989
rect 75361 247961 75389 247989
rect 90659 248147 90687 248175
rect 90721 248147 90749 248175
rect 90659 248085 90687 248113
rect 90721 248085 90749 248113
rect 90659 248023 90687 248051
rect 90721 248023 90749 248051
rect 90659 247961 90687 247989
rect 90721 247961 90749 247989
rect 106019 248147 106047 248175
rect 106081 248147 106109 248175
rect 106019 248085 106047 248113
rect 106081 248085 106109 248113
rect 106019 248023 106047 248051
rect 106081 248023 106109 248051
rect 106019 247961 106047 247989
rect 106081 247961 106109 247989
rect 121379 248147 121407 248175
rect 121441 248147 121469 248175
rect 121379 248085 121407 248113
rect 121441 248085 121469 248113
rect 121379 248023 121407 248051
rect 121441 248023 121469 248051
rect 121379 247961 121407 247989
rect 121441 247961 121469 247989
rect 136739 248147 136767 248175
rect 136801 248147 136829 248175
rect 136739 248085 136767 248113
rect 136801 248085 136829 248113
rect 136739 248023 136767 248051
rect 136801 248023 136829 248051
rect 136739 247961 136767 247989
rect 136801 247961 136829 247989
rect 52259 245147 52287 245175
rect 52321 245147 52349 245175
rect 52259 245085 52287 245113
rect 52321 245085 52349 245113
rect 52259 245023 52287 245051
rect 52321 245023 52349 245051
rect 52259 244961 52287 244989
rect 52321 244961 52349 244989
rect 67619 245147 67647 245175
rect 67681 245147 67709 245175
rect 67619 245085 67647 245113
rect 67681 245085 67709 245113
rect 67619 245023 67647 245051
rect 67681 245023 67709 245051
rect 67619 244961 67647 244989
rect 67681 244961 67709 244989
rect 82979 245147 83007 245175
rect 83041 245147 83069 245175
rect 82979 245085 83007 245113
rect 83041 245085 83069 245113
rect 82979 245023 83007 245051
rect 83041 245023 83069 245051
rect 82979 244961 83007 244989
rect 83041 244961 83069 244989
rect 98339 245147 98367 245175
rect 98401 245147 98429 245175
rect 98339 245085 98367 245113
rect 98401 245085 98429 245113
rect 98339 245023 98367 245051
rect 98401 245023 98429 245051
rect 98339 244961 98367 244989
rect 98401 244961 98429 244989
rect 113699 245147 113727 245175
rect 113761 245147 113789 245175
rect 113699 245085 113727 245113
rect 113761 245085 113789 245113
rect 113699 245023 113727 245051
rect 113761 245023 113789 245051
rect 113699 244961 113727 244989
rect 113761 244961 113789 244989
rect 129059 245147 129087 245175
rect 129121 245147 129149 245175
rect 129059 245085 129087 245113
rect 129121 245085 129149 245113
rect 129059 245023 129087 245051
rect 129121 245023 129149 245051
rect 129059 244961 129087 244989
rect 129121 244961 129149 244989
rect 144419 245147 144447 245175
rect 144481 245147 144509 245175
rect 144419 245085 144447 245113
rect 144481 245085 144509 245113
rect 144419 245023 144447 245051
rect 144481 245023 144509 245051
rect 144419 244961 144447 244989
rect 144481 244961 144509 244989
rect 154625 245147 154653 245175
rect 154687 245147 154715 245175
rect 154749 245147 154777 245175
rect 154811 245147 154839 245175
rect 154625 245085 154653 245113
rect 154687 245085 154715 245113
rect 154749 245085 154777 245113
rect 154811 245085 154839 245113
rect 154625 245023 154653 245051
rect 154687 245023 154715 245051
rect 154749 245023 154777 245051
rect 154811 245023 154839 245051
rect 154625 244961 154653 244989
rect 154687 244961 154715 244989
rect 154749 244961 154777 244989
rect 154811 244961 154839 244989
rect 48485 239147 48513 239175
rect 48547 239147 48575 239175
rect 48609 239147 48637 239175
rect 48671 239147 48699 239175
rect 48485 239085 48513 239113
rect 48547 239085 48575 239113
rect 48609 239085 48637 239113
rect 48671 239085 48699 239113
rect 48485 239023 48513 239051
rect 48547 239023 48575 239051
rect 48609 239023 48637 239051
rect 48671 239023 48699 239051
rect 48485 238961 48513 238989
rect 48547 238961 48575 238989
rect 48609 238961 48637 238989
rect 48671 238961 48699 238989
rect 59939 239147 59967 239175
rect 60001 239147 60029 239175
rect 59939 239085 59967 239113
rect 60001 239085 60029 239113
rect 59939 239023 59967 239051
rect 60001 239023 60029 239051
rect 59939 238961 59967 238989
rect 60001 238961 60029 238989
rect 75299 239147 75327 239175
rect 75361 239147 75389 239175
rect 75299 239085 75327 239113
rect 75361 239085 75389 239113
rect 75299 239023 75327 239051
rect 75361 239023 75389 239051
rect 75299 238961 75327 238989
rect 75361 238961 75389 238989
rect 90659 239147 90687 239175
rect 90721 239147 90749 239175
rect 90659 239085 90687 239113
rect 90721 239085 90749 239113
rect 90659 239023 90687 239051
rect 90721 239023 90749 239051
rect 90659 238961 90687 238989
rect 90721 238961 90749 238989
rect 106019 239147 106047 239175
rect 106081 239147 106109 239175
rect 106019 239085 106047 239113
rect 106081 239085 106109 239113
rect 106019 239023 106047 239051
rect 106081 239023 106109 239051
rect 106019 238961 106047 238989
rect 106081 238961 106109 238989
rect 121379 239147 121407 239175
rect 121441 239147 121469 239175
rect 121379 239085 121407 239113
rect 121441 239085 121469 239113
rect 121379 239023 121407 239051
rect 121441 239023 121469 239051
rect 121379 238961 121407 238989
rect 121441 238961 121469 238989
rect 136739 239147 136767 239175
rect 136801 239147 136829 239175
rect 136739 239085 136767 239113
rect 136801 239085 136829 239113
rect 136739 239023 136767 239051
rect 136801 239023 136829 239051
rect 136739 238961 136767 238989
rect 136801 238961 136829 238989
rect 52259 236147 52287 236175
rect 52321 236147 52349 236175
rect 52259 236085 52287 236113
rect 52321 236085 52349 236113
rect 52259 236023 52287 236051
rect 52321 236023 52349 236051
rect 52259 235961 52287 235989
rect 52321 235961 52349 235989
rect 67619 236147 67647 236175
rect 67681 236147 67709 236175
rect 67619 236085 67647 236113
rect 67681 236085 67709 236113
rect 67619 236023 67647 236051
rect 67681 236023 67709 236051
rect 67619 235961 67647 235989
rect 67681 235961 67709 235989
rect 82979 236147 83007 236175
rect 83041 236147 83069 236175
rect 82979 236085 83007 236113
rect 83041 236085 83069 236113
rect 82979 236023 83007 236051
rect 83041 236023 83069 236051
rect 82979 235961 83007 235989
rect 83041 235961 83069 235989
rect 98339 236147 98367 236175
rect 98401 236147 98429 236175
rect 98339 236085 98367 236113
rect 98401 236085 98429 236113
rect 98339 236023 98367 236051
rect 98401 236023 98429 236051
rect 98339 235961 98367 235989
rect 98401 235961 98429 235989
rect 113699 236147 113727 236175
rect 113761 236147 113789 236175
rect 113699 236085 113727 236113
rect 113761 236085 113789 236113
rect 113699 236023 113727 236051
rect 113761 236023 113789 236051
rect 113699 235961 113727 235989
rect 113761 235961 113789 235989
rect 129059 236147 129087 236175
rect 129121 236147 129149 236175
rect 129059 236085 129087 236113
rect 129121 236085 129149 236113
rect 129059 236023 129087 236051
rect 129121 236023 129149 236051
rect 129059 235961 129087 235989
rect 129121 235961 129149 235989
rect 144419 236147 144447 236175
rect 144481 236147 144509 236175
rect 144419 236085 144447 236113
rect 144481 236085 144509 236113
rect 144419 236023 144447 236051
rect 144481 236023 144509 236051
rect 144419 235961 144447 235989
rect 144481 235961 144509 235989
rect 154625 236147 154653 236175
rect 154687 236147 154715 236175
rect 154749 236147 154777 236175
rect 154811 236147 154839 236175
rect 154625 236085 154653 236113
rect 154687 236085 154715 236113
rect 154749 236085 154777 236113
rect 154811 236085 154839 236113
rect 154625 236023 154653 236051
rect 154687 236023 154715 236051
rect 154749 236023 154777 236051
rect 154811 236023 154839 236051
rect 154625 235961 154653 235989
rect 154687 235961 154715 235989
rect 154749 235961 154777 235989
rect 154811 235961 154839 235989
rect 48485 230147 48513 230175
rect 48547 230147 48575 230175
rect 48609 230147 48637 230175
rect 48671 230147 48699 230175
rect 48485 230085 48513 230113
rect 48547 230085 48575 230113
rect 48609 230085 48637 230113
rect 48671 230085 48699 230113
rect 48485 230023 48513 230051
rect 48547 230023 48575 230051
rect 48609 230023 48637 230051
rect 48671 230023 48699 230051
rect 48485 229961 48513 229989
rect 48547 229961 48575 229989
rect 48609 229961 48637 229989
rect 48671 229961 48699 229989
rect 59939 230147 59967 230175
rect 60001 230147 60029 230175
rect 59939 230085 59967 230113
rect 60001 230085 60029 230113
rect 59939 230023 59967 230051
rect 60001 230023 60029 230051
rect 59939 229961 59967 229989
rect 60001 229961 60029 229989
rect 75299 230147 75327 230175
rect 75361 230147 75389 230175
rect 75299 230085 75327 230113
rect 75361 230085 75389 230113
rect 75299 230023 75327 230051
rect 75361 230023 75389 230051
rect 75299 229961 75327 229989
rect 75361 229961 75389 229989
rect 90659 230147 90687 230175
rect 90721 230147 90749 230175
rect 90659 230085 90687 230113
rect 90721 230085 90749 230113
rect 90659 230023 90687 230051
rect 90721 230023 90749 230051
rect 90659 229961 90687 229989
rect 90721 229961 90749 229989
rect 106019 230147 106047 230175
rect 106081 230147 106109 230175
rect 106019 230085 106047 230113
rect 106081 230085 106109 230113
rect 106019 230023 106047 230051
rect 106081 230023 106109 230051
rect 106019 229961 106047 229989
rect 106081 229961 106109 229989
rect 121379 230147 121407 230175
rect 121441 230147 121469 230175
rect 121379 230085 121407 230113
rect 121441 230085 121469 230113
rect 121379 230023 121407 230051
rect 121441 230023 121469 230051
rect 121379 229961 121407 229989
rect 121441 229961 121469 229989
rect 136739 230147 136767 230175
rect 136801 230147 136829 230175
rect 136739 230085 136767 230113
rect 136801 230085 136829 230113
rect 136739 230023 136767 230051
rect 136801 230023 136829 230051
rect 136739 229961 136767 229989
rect 136801 229961 136829 229989
rect 52259 227147 52287 227175
rect 52321 227147 52349 227175
rect 52259 227085 52287 227113
rect 52321 227085 52349 227113
rect 52259 227023 52287 227051
rect 52321 227023 52349 227051
rect 52259 226961 52287 226989
rect 52321 226961 52349 226989
rect 67619 227147 67647 227175
rect 67681 227147 67709 227175
rect 67619 227085 67647 227113
rect 67681 227085 67709 227113
rect 67619 227023 67647 227051
rect 67681 227023 67709 227051
rect 67619 226961 67647 226989
rect 67681 226961 67709 226989
rect 82979 227147 83007 227175
rect 83041 227147 83069 227175
rect 82979 227085 83007 227113
rect 83041 227085 83069 227113
rect 82979 227023 83007 227051
rect 83041 227023 83069 227051
rect 82979 226961 83007 226989
rect 83041 226961 83069 226989
rect 98339 227147 98367 227175
rect 98401 227147 98429 227175
rect 98339 227085 98367 227113
rect 98401 227085 98429 227113
rect 98339 227023 98367 227051
rect 98401 227023 98429 227051
rect 98339 226961 98367 226989
rect 98401 226961 98429 226989
rect 113699 227147 113727 227175
rect 113761 227147 113789 227175
rect 113699 227085 113727 227113
rect 113761 227085 113789 227113
rect 113699 227023 113727 227051
rect 113761 227023 113789 227051
rect 113699 226961 113727 226989
rect 113761 226961 113789 226989
rect 129059 227147 129087 227175
rect 129121 227147 129149 227175
rect 129059 227085 129087 227113
rect 129121 227085 129149 227113
rect 129059 227023 129087 227051
rect 129121 227023 129149 227051
rect 129059 226961 129087 226989
rect 129121 226961 129149 226989
rect 144419 227147 144447 227175
rect 144481 227147 144509 227175
rect 144419 227085 144447 227113
rect 144481 227085 144509 227113
rect 144419 227023 144447 227051
rect 144481 227023 144509 227051
rect 144419 226961 144447 226989
rect 144481 226961 144509 226989
rect 154625 227147 154653 227175
rect 154687 227147 154715 227175
rect 154749 227147 154777 227175
rect 154811 227147 154839 227175
rect 154625 227085 154653 227113
rect 154687 227085 154715 227113
rect 154749 227085 154777 227113
rect 154811 227085 154839 227113
rect 154625 227023 154653 227051
rect 154687 227023 154715 227051
rect 154749 227023 154777 227051
rect 154811 227023 154839 227051
rect 154625 226961 154653 226989
rect 154687 226961 154715 226989
rect 154749 226961 154777 226989
rect 154811 226961 154839 226989
rect 48485 221147 48513 221175
rect 48547 221147 48575 221175
rect 48609 221147 48637 221175
rect 48671 221147 48699 221175
rect 48485 221085 48513 221113
rect 48547 221085 48575 221113
rect 48609 221085 48637 221113
rect 48671 221085 48699 221113
rect 48485 221023 48513 221051
rect 48547 221023 48575 221051
rect 48609 221023 48637 221051
rect 48671 221023 48699 221051
rect 48485 220961 48513 220989
rect 48547 220961 48575 220989
rect 48609 220961 48637 220989
rect 48671 220961 48699 220989
rect 59939 221147 59967 221175
rect 60001 221147 60029 221175
rect 59939 221085 59967 221113
rect 60001 221085 60029 221113
rect 59939 221023 59967 221051
rect 60001 221023 60029 221051
rect 59939 220961 59967 220989
rect 60001 220961 60029 220989
rect 75299 221147 75327 221175
rect 75361 221147 75389 221175
rect 75299 221085 75327 221113
rect 75361 221085 75389 221113
rect 75299 221023 75327 221051
rect 75361 221023 75389 221051
rect 75299 220961 75327 220989
rect 75361 220961 75389 220989
rect 90659 221147 90687 221175
rect 90721 221147 90749 221175
rect 90659 221085 90687 221113
rect 90721 221085 90749 221113
rect 90659 221023 90687 221051
rect 90721 221023 90749 221051
rect 90659 220961 90687 220989
rect 90721 220961 90749 220989
rect 106019 221147 106047 221175
rect 106081 221147 106109 221175
rect 106019 221085 106047 221113
rect 106081 221085 106109 221113
rect 106019 221023 106047 221051
rect 106081 221023 106109 221051
rect 106019 220961 106047 220989
rect 106081 220961 106109 220989
rect 121379 221147 121407 221175
rect 121441 221147 121469 221175
rect 121379 221085 121407 221113
rect 121441 221085 121469 221113
rect 121379 221023 121407 221051
rect 121441 221023 121469 221051
rect 121379 220961 121407 220989
rect 121441 220961 121469 220989
rect 136739 221147 136767 221175
rect 136801 221147 136829 221175
rect 136739 221085 136767 221113
rect 136801 221085 136829 221113
rect 136739 221023 136767 221051
rect 136801 221023 136829 221051
rect 136739 220961 136767 220989
rect 136801 220961 136829 220989
rect 52259 218147 52287 218175
rect 52321 218147 52349 218175
rect 52259 218085 52287 218113
rect 52321 218085 52349 218113
rect 52259 218023 52287 218051
rect 52321 218023 52349 218051
rect 52259 217961 52287 217989
rect 52321 217961 52349 217989
rect 67619 218147 67647 218175
rect 67681 218147 67709 218175
rect 67619 218085 67647 218113
rect 67681 218085 67709 218113
rect 67619 218023 67647 218051
rect 67681 218023 67709 218051
rect 67619 217961 67647 217989
rect 67681 217961 67709 217989
rect 82979 218147 83007 218175
rect 83041 218147 83069 218175
rect 82979 218085 83007 218113
rect 83041 218085 83069 218113
rect 82979 218023 83007 218051
rect 83041 218023 83069 218051
rect 82979 217961 83007 217989
rect 83041 217961 83069 217989
rect 98339 218147 98367 218175
rect 98401 218147 98429 218175
rect 98339 218085 98367 218113
rect 98401 218085 98429 218113
rect 98339 218023 98367 218051
rect 98401 218023 98429 218051
rect 98339 217961 98367 217989
rect 98401 217961 98429 217989
rect 113699 218147 113727 218175
rect 113761 218147 113789 218175
rect 113699 218085 113727 218113
rect 113761 218085 113789 218113
rect 113699 218023 113727 218051
rect 113761 218023 113789 218051
rect 113699 217961 113727 217989
rect 113761 217961 113789 217989
rect 129059 218147 129087 218175
rect 129121 218147 129149 218175
rect 129059 218085 129087 218113
rect 129121 218085 129149 218113
rect 129059 218023 129087 218051
rect 129121 218023 129149 218051
rect 129059 217961 129087 217989
rect 129121 217961 129149 217989
rect 144419 218147 144447 218175
rect 144481 218147 144509 218175
rect 144419 218085 144447 218113
rect 144481 218085 144509 218113
rect 144419 218023 144447 218051
rect 144481 218023 144509 218051
rect 144419 217961 144447 217989
rect 144481 217961 144509 217989
rect 154625 218147 154653 218175
rect 154687 218147 154715 218175
rect 154749 218147 154777 218175
rect 154811 218147 154839 218175
rect 154625 218085 154653 218113
rect 154687 218085 154715 218113
rect 154749 218085 154777 218113
rect 154811 218085 154839 218113
rect 154625 218023 154653 218051
rect 154687 218023 154715 218051
rect 154749 218023 154777 218051
rect 154811 218023 154839 218051
rect 154625 217961 154653 217989
rect 154687 217961 154715 217989
rect 154749 217961 154777 217989
rect 154811 217961 154839 217989
rect 48485 212147 48513 212175
rect 48547 212147 48575 212175
rect 48609 212147 48637 212175
rect 48671 212147 48699 212175
rect 48485 212085 48513 212113
rect 48547 212085 48575 212113
rect 48609 212085 48637 212113
rect 48671 212085 48699 212113
rect 48485 212023 48513 212051
rect 48547 212023 48575 212051
rect 48609 212023 48637 212051
rect 48671 212023 48699 212051
rect 48485 211961 48513 211989
rect 48547 211961 48575 211989
rect 48609 211961 48637 211989
rect 48671 211961 48699 211989
rect 59939 212147 59967 212175
rect 60001 212147 60029 212175
rect 59939 212085 59967 212113
rect 60001 212085 60029 212113
rect 59939 212023 59967 212051
rect 60001 212023 60029 212051
rect 59939 211961 59967 211989
rect 60001 211961 60029 211989
rect 75299 212147 75327 212175
rect 75361 212147 75389 212175
rect 75299 212085 75327 212113
rect 75361 212085 75389 212113
rect 75299 212023 75327 212051
rect 75361 212023 75389 212051
rect 75299 211961 75327 211989
rect 75361 211961 75389 211989
rect 90659 212147 90687 212175
rect 90721 212147 90749 212175
rect 90659 212085 90687 212113
rect 90721 212085 90749 212113
rect 90659 212023 90687 212051
rect 90721 212023 90749 212051
rect 90659 211961 90687 211989
rect 90721 211961 90749 211989
rect 106019 212147 106047 212175
rect 106081 212147 106109 212175
rect 106019 212085 106047 212113
rect 106081 212085 106109 212113
rect 106019 212023 106047 212051
rect 106081 212023 106109 212051
rect 106019 211961 106047 211989
rect 106081 211961 106109 211989
rect 121379 212147 121407 212175
rect 121441 212147 121469 212175
rect 121379 212085 121407 212113
rect 121441 212085 121469 212113
rect 121379 212023 121407 212051
rect 121441 212023 121469 212051
rect 121379 211961 121407 211989
rect 121441 211961 121469 211989
rect 136739 212147 136767 212175
rect 136801 212147 136829 212175
rect 136739 212085 136767 212113
rect 136801 212085 136829 212113
rect 136739 212023 136767 212051
rect 136801 212023 136829 212051
rect 136739 211961 136767 211989
rect 136801 211961 136829 211989
rect 52259 209147 52287 209175
rect 52321 209147 52349 209175
rect 52259 209085 52287 209113
rect 52321 209085 52349 209113
rect 52259 209023 52287 209051
rect 52321 209023 52349 209051
rect 52259 208961 52287 208989
rect 52321 208961 52349 208989
rect 67619 209147 67647 209175
rect 67681 209147 67709 209175
rect 67619 209085 67647 209113
rect 67681 209085 67709 209113
rect 67619 209023 67647 209051
rect 67681 209023 67709 209051
rect 67619 208961 67647 208989
rect 67681 208961 67709 208989
rect 82979 209147 83007 209175
rect 83041 209147 83069 209175
rect 82979 209085 83007 209113
rect 83041 209085 83069 209113
rect 82979 209023 83007 209051
rect 83041 209023 83069 209051
rect 82979 208961 83007 208989
rect 83041 208961 83069 208989
rect 98339 209147 98367 209175
rect 98401 209147 98429 209175
rect 98339 209085 98367 209113
rect 98401 209085 98429 209113
rect 98339 209023 98367 209051
rect 98401 209023 98429 209051
rect 98339 208961 98367 208989
rect 98401 208961 98429 208989
rect 113699 209147 113727 209175
rect 113761 209147 113789 209175
rect 113699 209085 113727 209113
rect 113761 209085 113789 209113
rect 113699 209023 113727 209051
rect 113761 209023 113789 209051
rect 113699 208961 113727 208989
rect 113761 208961 113789 208989
rect 129059 209147 129087 209175
rect 129121 209147 129149 209175
rect 129059 209085 129087 209113
rect 129121 209085 129149 209113
rect 129059 209023 129087 209051
rect 129121 209023 129149 209051
rect 129059 208961 129087 208989
rect 129121 208961 129149 208989
rect 144419 209147 144447 209175
rect 144481 209147 144509 209175
rect 144419 209085 144447 209113
rect 144481 209085 144509 209113
rect 144419 209023 144447 209051
rect 144481 209023 144509 209051
rect 144419 208961 144447 208989
rect 144481 208961 144509 208989
rect 154625 209147 154653 209175
rect 154687 209147 154715 209175
rect 154749 209147 154777 209175
rect 154811 209147 154839 209175
rect 154625 209085 154653 209113
rect 154687 209085 154715 209113
rect 154749 209085 154777 209113
rect 154811 209085 154839 209113
rect 154625 209023 154653 209051
rect 154687 209023 154715 209051
rect 154749 209023 154777 209051
rect 154811 209023 154839 209051
rect 154625 208961 154653 208989
rect 154687 208961 154715 208989
rect 154749 208961 154777 208989
rect 154811 208961 154839 208989
rect 48485 203147 48513 203175
rect 48547 203147 48575 203175
rect 48609 203147 48637 203175
rect 48671 203147 48699 203175
rect 48485 203085 48513 203113
rect 48547 203085 48575 203113
rect 48609 203085 48637 203113
rect 48671 203085 48699 203113
rect 48485 203023 48513 203051
rect 48547 203023 48575 203051
rect 48609 203023 48637 203051
rect 48671 203023 48699 203051
rect 48485 202961 48513 202989
rect 48547 202961 48575 202989
rect 48609 202961 48637 202989
rect 48671 202961 48699 202989
rect 59939 203147 59967 203175
rect 60001 203147 60029 203175
rect 59939 203085 59967 203113
rect 60001 203085 60029 203113
rect 59939 203023 59967 203051
rect 60001 203023 60029 203051
rect 59939 202961 59967 202989
rect 60001 202961 60029 202989
rect 75299 203147 75327 203175
rect 75361 203147 75389 203175
rect 75299 203085 75327 203113
rect 75361 203085 75389 203113
rect 75299 203023 75327 203051
rect 75361 203023 75389 203051
rect 75299 202961 75327 202989
rect 75361 202961 75389 202989
rect 90659 203147 90687 203175
rect 90721 203147 90749 203175
rect 90659 203085 90687 203113
rect 90721 203085 90749 203113
rect 90659 203023 90687 203051
rect 90721 203023 90749 203051
rect 90659 202961 90687 202989
rect 90721 202961 90749 202989
rect 106019 203147 106047 203175
rect 106081 203147 106109 203175
rect 106019 203085 106047 203113
rect 106081 203085 106109 203113
rect 106019 203023 106047 203051
rect 106081 203023 106109 203051
rect 106019 202961 106047 202989
rect 106081 202961 106109 202989
rect 121379 203147 121407 203175
rect 121441 203147 121469 203175
rect 121379 203085 121407 203113
rect 121441 203085 121469 203113
rect 121379 203023 121407 203051
rect 121441 203023 121469 203051
rect 121379 202961 121407 202989
rect 121441 202961 121469 202989
rect 136739 203147 136767 203175
rect 136801 203147 136829 203175
rect 136739 203085 136767 203113
rect 136801 203085 136829 203113
rect 136739 203023 136767 203051
rect 136801 203023 136829 203051
rect 136739 202961 136767 202989
rect 136801 202961 136829 202989
rect 154625 200147 154653 200175
rect 154687 200147 154715 200175
rect 154749 200147 154777 200175
rect 154811 200147 154839 200175
rect 154625 200085 154653 200113
rect 154687 200085 154715 200113
rect 154749 200085 154777 200113
rect 154811 200085 154839 200113
rect 154625 200023 154653 200051
rect 154687 200023 154715 200051
rect 154749 200023 154777 200051
rect 154811 200023 154839 200051
rect 154625 199961 154653 199989
rect 154687 199961 154715 199989
rect 154749 199961 154777 199989
rect 154811 199961 154839 199989
rect 48485 194147 48513 194175
rect 48547 194147 48575 194175
rect 48609 194147 48637 194175
rect 48671 194147 48699 194175
rect 48485 194085 48513 194113
rect 48547 194085 48575 194113
rect 48609 194085 48637 194113
rect 48671 194085 48699 194113
rect 48485 194023 48513 194051
rect 48547 194023 48575 194051
rect 48609 194023 48637 194051
rect 48671 194023 48699 194051
rect 48485 193961 48513 193989
rect 48547 193961 48575 193989
rect 48609 193961 48637 193989
rect 48671 193961 48699 193989
rect 48485 185147 48513 185175
rect 48547 185147 48575 185175
rect 48609 185147 48637 185175
rect 48671 185147 48699 185175
rect 48485 185085 48513 185113
rect 48547 185085 48575 185113
rect 48609 185085 48637 185113
rect 48671 185085 48699 185113
rect 48485 185023 48513 185051
rect 48547 185023 48575 185051
rect 48609 185023 48637 185051
rect 48671 185023 48699 185051
rect 48485 184961 48513 184989
rect 48547 184961 48575 184989
rect 48609 184961 48637 184989
rect 48671 184961 48699 184989
rect 57485 194147 57513 194175
rect 57547 194147 57575 194175
rect 57609 194147 57637 194175
rect 57671 194147 57699 194175
rect 57485 194085 57513 194113
rect 57547 194085 57575 194113
rect 57609 194085 57637 194113
rect 57671 194085 57699 194113
rect 57485 194023 57513 194051
rect 57547 194023 57575 194051
rect 57609 194023 57637 194051
rect 57671 194023 57699 194051
rect 57485 193961 57513 193989
rect 57547 193961 57575 193989
rect 57609 193961 57637 193989
rect 57671 193961 57699 193989
rect 57485 185147 57513 185175
rect 57547 185147 57575 185175
rect 57609 185147 57637 185175
rect 57671 185147 57699 185175
rect 57485 185085 57513 185113
rect 57547 185085 57575 185113
rect 57609 185085 57637 185113
rect 57671 185085 57699 185113
rect 57485 185023 57513 185051
rect 57547 185023 57575 185051
rect 57609 185023 57637 185051
rect 57671 185023 57699 185051
rect 57485 184961 57513 184989
rect 57547 184961 57575 184989
rect 57609 184961 57637 184989
rect 57671 184961 57699 184989
rect 66485 194147 66513 194175
rect 66547 194147 66575 194175
rect 66609 194147 66637 194175
rect 66671 194147 66699 194175
rect 66485 194085 66513 194113
rect 66547 194085 66575 194113
rect 66609 194085 66637 194113
rect 66671 194085 66699 194113
rect 66485 194023 66513 194051
rect 66547 194023 66575 194051
rect 66609 194023 66637 194051
rect 66671 194023 66699 194051
rect 66485 193961 66513 193989
rect 66547 193961 66575 193989
rect 66609 193961 66637 193989
rect 66671 193961 66699 193989
rect 66485 185147 66513 185175
rect 66547 185147 66575 185175
rect 66609 185147 66637 185175
rect 66671 185147 66699 185175
rect 66485 185085 66513 185113
rect 66547 185085 66575 185113
rect 66609 185085 66637 185113
rect 66671 185085 66699 185113
rect 66485 185023 66513 185051
rect 66547 185023 66575 185051
rect 66609 185023 66637 185051
rect 66671 185023 66699 185051
rect 66485 184961 66513 184989
rect 66547 184961 66575 184989
rect 66609 184961 66637 184989
rect 66671 184961 66699 184989
rect 75485 194147 75513 194175
rect 75547 194147 75575 194175
rect 75609 194147 75637 194175
rect 75671 194147 75699 194175
rect 75485 194085 75513 194113
rect 75547 194085 75575 194113
rect 75609 194085 75637 194113
rect 75671 194085 75699 194113
rect 75485 194023 75513 194051
rect 75547 194023 75575 194051
rect 75609 194023 75637 194051
rect 75671 194023 75699 194051
rect 75485 193961 75513 193989
rect 75547 193961 75575 193989
rect 75609 193961 75637 193989
rect 75671 193961 75699 193989
rect 75485 185147 75513 185175
rect 75547 185147 75575 185175
rect 75609 185147 75637 185175
rect 75671 185147 75699 185175
rect 75485 185085 75513 185113
rect 75547 185085 75575 185113
rect 75609 185085 75637 185113
rect 75671 185085 75699 185113
rect 75485 185023 75513 185051
rect 75547 185023 75575 185051
rect 75609 185023 75637 185051
rect 75671 185023 75699 185051
rect 75485 184961 75513 184989
rect 75547 184961 75575 184989
rect 75609 184961 75637 184989
rect 75671 184961 75699 184989
rect 84485 194147 84513 194175
rect 84547 194147 84575 194175
rect 84609 194147 84637 194175
rect 84671 194147 84699 194175
rect 84485 194085 84513 194113
rect 84547 194085 84575 194113
rect 84609 194085 84637 194113
rect 84671 194085 84699 194113
rect 84485 194023 84513 194051
rect 84547 194023 84575 194051
rect 84609 194023 84637 194051
rect 84671 194023 84699 194051
rect 84485 193961 84513 193989
rect 84547 193961 84575 193989
rect 84609 193961 84637 193989
rect 84671 193961 84699 193989
rect 84485 185147 84513 185175
rect 84547 185147 84575 185175
rect 84609 185147 84637 185175
rect 84671 185147 84699 185175
rect 84485 185085 84513 185113
rect 84547 185085 84575 185113
rect 84609 185085 84637 185113
rect 84671 185085 84699 185113
rect 84485 185023 84513 185051
rect 84547 185023 84575 185051
rect 84609 185023 84637 185051
rect 84671 185023 84699 185051
rect 84485 184961 84513 184989
rect 84547 184961 84575 184989
rect 84609 184961 84637 184989
rect 84671 184961 84699 184989
rect 93485 194147 93513 194175
rect 93547 194147 93575 194175
rect 93609 194147 93637 194175
rect 93671 194147 93699 194175
rect 93485 194085 93513 194113
rect 93547 194085 93575 194113
rect 93609 194085 93637 194113
rect 93671 194085 93699 194113
rect 93485 194023 93513 194051
rect 93547 194023 93575 194051
rect 93609 194023 93637 194051
rect 93671 194023 93699 194051
rect 93485 193961 93513 193989
rect 93547 193961 93575 193989
rect 93609 193961 93637 193989
rect 93671 193961 93699 193989
rect 93485 185147 93513 185175
rect 93547 185147 93575 185175
rect 93609 185147 93637 185175
rect 93671 185147 93699 185175
rect 93485 185085 93513 185113
rect 93547 185085 93575 185113
rect 93609 185085 93637 185113
rect 93671 185085 93699 185113
rect 93485 185023 93513 185051
rect 93547 185023 93575 185051
rect 93609 185023 93637 185051
rect 93671 185023 93699 185051
rect 93485 184961 93513 184989
rect 93547 184961 93575 184989
rect 93609 184961 93637 184989
rect 93671 184961 93699 184989
rect 102485 194147 102513 194175
rect 102547 194147 102575 194175
rect 102609 194147 102637 194175
rect 102671 194147 102699 194175
rect 102485 194085 102513 194113
rect 102547 194085 102575 194113
rect 102609 194085 102637 194113
rect 102671 194085 102699 194113
rect 102485 194023 102513 194051
rect 102547 194023 102575 194051
rect 102609 194023 102637 194051
rect 102671 194023 102699 194051
rect 102485 193961 102513 193989
rect 102547 193961 102575 193989
rect 102609 193961 102637 193989
rect 102671 193961 102699 193989
rect 102485 185147 102513 185175
rect 102547 185147 102575 185175
rect 102609 185147 102637 185175
rect 102671 185147 102699 185175
rect 102485 185085 102513 185113
rect 102547 185085 102575 185113
rect 102609 185085 102637 185113
rect 102671 185085 102699 185113
rect 102485 185023 102513 185051
rect 102547 185023 102575 185051
rect 102609 185023 102637 185051
rect 102671 185023 102699 185051
rect 102485 184961 102513 184989
rect 102547 184961 102575 184989
rect 102609 184961 102637 184989
rect 102671 184961 102699 184989
rect 111485 194147 111513 194175
rect 111547 194147 111575 194175
rect 111609 194147 111637 194175
rect 111671 194147 111699 194175
rect 111485 194085 111513 194113
rect 111547 194085 111575 194113
rect 111609 194085 111637 194113
rect 111671 194085 111699 194113
rect 111485 194023 111513 194051
rect 111547 194023 111575 194051
rect 111609 194023 111637 194051
rect 111671 194023 111699 194051
rect 111485 193961 111513 193989
rect 111547 193961 111575 193989
rect 111609 193961 111637 193989
rect 111671 193961 111699 193989
rect 111485 185147 111513 185175
rect 111547 185147 111575 185175
rect 111609 185147 111637 185175
rect 111671 185147 111699 185175
rect 111485 185085 111513 185113
rect 111547 185085 111575 185113
rect 111609 185085 111637 185113
rect 111671 185085 111699 185113
rect 111485 185023 111513 185051
rect 111547 185023 111575 185051
rect 111609 185023 111637 185051
rect 111671 185023 111699 185051
rect 111485 184961 111513 184989
rect 111547 184961 111575 184989
rect 111609 184961 111637 184989
rect 111671 184961 111699 184989
rect 120485 194147 120513 194175
rect 120547 194147 120575 194175
rect 120609 194147 120637 194175
rect 120671 194147 120699 194175
rect 120485 194085 120513 194113
rect 120547 194085 120575 194113
rect 120609 194085 120637 194113
rect 120671 194085 120699 194113
rect 120485 194023 120513 194051
rect 120547 194023 120575 194051
rect 120609 194023 120637 194051
rect 120671 194023 120699 194051
rect 120485 193961 120513 193989
rect 120547 193961 120575 193989
rect 120609 193961 120637 193989
rect 120671 193961 120699 193989
rect 120485 185147 120513 185175
rect 120547 185147 120575 185175
rect 120609 185147 120637 185175
rect 120671 185147 120699 185175
rect 120485 185085 120513 185113
rect 120547 185085 120575 185113
rect 120609 185085 120637 185113
rect 120671 185085 120699 185113
rect 120485 185023 120513 185051
rect 120547 185023 120575 185051
rect 120609 185023 120637 185051
rect 120671 185023 120699 185051
rect 120485 184961 120513 184989
rect 120547 184961 120575 184989
rect 120609 184961 120637 184989
rect 120671 184961 120699 184989
rect 129485 194147 129513 194175
rect 129547 194147 129575 194175
rect 129609 194147 129637 194175
rect 129671 194147 129699 194175
rect 129485 194085 129513 194113
rect 129547 194085 129575 194113
rect 129609 194085 129637 194113
rect 129671 194085 129699 194113
rect 129485 194023 129513 194051
rect 129547 194023 129575 194051
rect 129609 194023 129637 194051
rect 129671 194023 129699 194051
rect 129485 193961 129513 193989
rect 129547 193961 129575 193989
rect 129609 193961 129637 193989
rect 129671 193961 129699 193989
rect 129485 185147 129513 185175
rect 129547 185147 129575 185175
rect 129609 185147 129637 185175
rect 129671 185147 129699 185175
rect 129485 185085 129513 185113
rect 129547 185085 129575 185113
rect 129609 185085 129637 185113
rect 129671 185085 129699 185113
rect 129485 185023 129513 185051
rect 129547 185023 129575 185051
rect 129609 185023 129637 185051
rect 129671 185023 129699 185051
rect 129485 184961 129513 184989
rect 129547 184961 129575 184989
rect 129609 184961 129637 184989
rect 129671 184961 129699 184989
rect 138485 194147 138513 194175
rect 138547 194147 138575 194175
rect 138609 194147 138637 194175
rect 138671 194147 138699 194175
rect 138485 194085 138513 194113
rect 138547 194085 138575 194113
rect 138609 194085 138637 194113
rect 138671 194085 138699 194113
rect 138485 194023 138513 194051
rect 138547 194023 138575 194051
rect 138609 194023 138637 194051
rect 138671 194023 138699 194051
rect 138485 193961 138513 193989
rect 138547 193961 138575 193989
rect 138609 193961 138637 193989
rect 138671 193961 138699 193989
rect 138485 185147 138513 185175
rect 138547 185147 138575 185175
rect 138609 185147 138637 185175
rect 138671 185147 138699 185175
rect 138485 185085 138513 185113
rect 138547 185085 138575 185113
rect 138609 185085 138637 185113
rect 138671 185085 138699 185113
rect 138485 185023 138513 185051
rect 138547 185023 138575 185051
rect 138609 185023 138637 185051
rect 138671 185023 138699 185051
rect 138485 184961 138513 184989
rect 138547 184961 138575 184989
rect 138609 184961 138637 184989
rect 138671 184961 138699 184989
rect 147485 194147 147513 194175
rect 147547 194147 147575 194175
rect 147609 194147 147637 194175
rect 147671 194147 147699 194175
rect 147485 194085 147513 194113
rect 147547 194085 147575 194113
rect 147609 194085 147637 194113
rect 147671 194085 147699 194113
rect 147485 194023 147513 194051
rect 147547 194023 147575 194051
rect 147609 194023 147637 194051
rect 147671 194023 147699 194051
rect 147485 193961 147513 193989
rect 147547 193961 147575 193989
rect 147609 193961 147637 193989
rect 147671 193961 147699 193989
rect 147485 185147 147513 185175
rect 147547 185147 147575 185175
rect 147609 185147 147637 185175
rect 147671 185147 147699 185175
rect 147485 185085 147513 185113
rect 147547 185085 147575 185113
rect 147609 185085 147637 185113
rect 147671 185085 147699 185113
rect 147485 185023 147513 185051
rect 147547 185023 147575 185051
rect 147609 185023 147637 185051
rect 147671 185023 147699 185051
rect 147485 184961 147513 184989
rect 147547 184961 147575 184989
rect 147609 184961 147637 184989
rect 147671 184961 147699 184989
rect 154625 191147 154653 191175
rect 154687 191147 154715 191175
rect 154749 191147 154777 191175
rect 154811 191147 154839 191175
rect 154625 191085 154653 191113
rect 154687 191085 154715 191113
rect 154749 191085 154777 191113
rect 154811 191085 154839 191113
rect 154625 191023 154653 191051
rect 154687 191023 154715 191051
rect 154749 191023 154777 191051
rect 154811 191023 154839 191051
rect 154625 190961 154653 190989
rect 154687 190961 154715 190989
rect 154749 190961 154777 190989
rect 154811 190961 154839 190989
rect 52259 182147 52287 182175
rect 52321 182147 52349 182175
rect 52259 182085 52287 182113
rect 52321 182085 52349 182113
rect 52259 182023 52287 182051
rect 52321 182023 52349 182051
rect 52259 181961 52287 181989
rect 52321 181961 52349 181989
rect 67619 182147 67647 182175
rect 67681 182147 67709 182175
rect 67619 182085 67647 182113
rect 67681 182085 67709 182113
rect 67619 182023 67647 182051
rect 67681 182023 67709 182051
rect 67619 181961 67647 181989
rect 67681 181961 67709 181989
rect 82979 182147 83007 182175
rect 83041 182147 83069 182175
rect 82979 182085 83007 182113
rect 83041 182085 83069 182113
rect 82979 182023 83007 182051
rect 83041 182023 83069 182051
rect 82979 181961 83007 181989
rect 83041 181961 83069 181989
rect 98339 182147 98367 182175
rect 98401 182147 98429 182175
rect 98339 182085 98367 182113
rect 98401 182085 98429 182113
rect 98339 182023 98367 182051
rect 98401 182023 98429 182051
rect 98339 181961 98367 181989
rect 98401 181961 98429 181989
rect 113699 182147 113727 182175
rect 113761 182147 113789 182175
rect 113699 182085 113727 182113
rect 113761 182085 113789 182113
rect 113699 182023 113727 182051
rect 113761 182023 113789 182051
rect 113699 181961 113727 181989
rect 113761 181961 113789 181989
rect 129059 182147 129087 182175
rect 129121 182147 129149 182175
rect 129059 182085 129087 182113
rect 129121 182085 129149 182113
rect 129059 182023 129087 182051
rect 129121 182023 129149 182051
rect 129059 181961 129087 181989
rect 129121 181961 129149 181989
rect 144419 182147 144447 182175
rect 144481 182147 144509 182175
rect 144419 182085 144447 182113
rect 144481 182085 144509 182113
rect 144419 182023 144447 182051
rect 144481 182023 144509 182051
rect 144419 181961 144447 181989
rect 144481 181961 144509 181989
rect 154625 182147 154653 182175
rect 154687 182147 154715 182175
rect 154749 182147 154777 182175
rect 154811 182147 154839 182175
rect 154625 182085 154653 182113
rect 154687 182085 154715 182113
rect 154749 182085 154777 182113
rect 154811 182085 154839 182113
rect 154625 182023 154653 182051
rect 154687 182023 154715 182051
rect 154749 182023 154777 182051
rect 154811 182023 154839 182051
rect 154625 181961 154653 181989
rect 154687 181961 154715 181989
rect 154749 181961 154777 181989
rect 154811 181961 154839 181989
rect 48485 176147 48513 176175
rect 48547 176147 48575 176175
rect 48609 176147 48637 176175
rect 48671 176147 48699 176175
rect 48485 176085 48513 176113
rect 48547 176085 48575 176113
rect 48609 176085 48637 176113
rect 48671 176085 48699 176113
rect 48485 176023 48513 176051
rect 48547 176023 48575 176051
rect 48609 176023 48637 176051
rect 48671 176023 48699 176051
rect 48485 175961 48513 175989
rect 48547 175961 48575 175989
rect 48609 175961 48637 175989
rect 48671 175961 48699 175989
rect 59939 176147 59967 176175
rect 60001 176147 60029 176175
rect 59939 176085 59967 176113
rect 60001 176085 60029 176113
rect 59939 176023 59967 176051
rect 60001 176023 60029 176051
rect 59939 175961 59967 175989
rect 60001 175961 60029 175989
rect 75299 176147 75327 176175
rect 75361 176147 75389 176175
rect 75299 176085 75327 176113
rect 75361 176085 75389 176113
rect 75299 176023 75327 176051
rect 75361 176023 75389 176051
rect 75299 175961 75327 175989
rect 75361 175961 75389 175989
rect 90659 176147 90687 176175
rect 90721 176147 90749 176175
rect 90659 176085 90687 176113
rect 90721 176085 90749 176113
rect 90659 176023 90687 176051
rect 90721 176023 90749 176051
rect 90659 175961 90687 175989
rect 90721 175961 90749 175989
rect 106019 176147 106047 176175
rect 106081 176147 106109 176175
rect 106019 176085 106047 176113
rect 106081 176085 106109 176113
rect 106019 176023 106047 176051
rect 106081 176023 106109 176051
rect 106019 175961 106047 175989
rect 106081 175961 106109 175989
rect 121379 176147 121407 176175
rect 121441 176147 121469 176175
rect 121379 176085 121407 176113
rect 121441 176085 121469 176113
rect 121379 176023 121407 176051
rect 121441 176023 121469 176051
rect 121379 175961 121407 175989
rect 121441 175961 121469 175989
rect 136739 176147 136767 176175
rect 136801 176147 136829 176175
rect 136739 176085 136767 176113
rect 136801 176085 136829 176113
rect 136739 176023 136767 176051
rect 136801 176023 136829 176051
rect 136739 175961 136767 175989
rect 136801 175961 136829 175989
rect 52259 173147 52287 173175
rect 52321 173147 52349 173175
rect 52259 173085 52287 173113
rect 52321 173085 52349 173113
rect 52259 173023 52287 173051
rect 52321 173023 52349 173051
rect 52259 172961 52287 172989
rect 52321 172961 52349 172989
rect 67619 173147 67647 173175
rect 67681 173147 67709 173175
rect 67619 173085 67647 173113
rect 67681 173085 67709 173113
rect 67619 173023 67647 173051
rect 67681 173023 67709 173051
rect 67619 172961 67647 172989
rect 67681 172961 67709 172989
rect 82979 173147 83007 173175
rect 83041 173147 83069 173175
rect 82979 173085 83007 173113
rect 83041 173085 83069 173113
rect 82979 173023 83007 173051
rect 83041 173023 83069 173051
rect 82979 172961 83007 172989
rect 83041 172961 83069 172989
rect 98339 173147 98367 173175
rect 98401 173147 98429 173175
rect 98339 173085 98367 173113
rect 98401 173085 98429 173113
rect 98339 173023 98367 173051
rect 98401 173023 98429 173051
rect 98339 172961 98367 172989
rect 98401 172961 98429 172989
rect 113699 173147 113727 173175
rect 113761 173147 113789 173175
rect 113699 173085 113727 173113
rect 113761 173085 113789 173113
rect 113699 173023 113727 173051
rect 113761 173023 113789 173051
rect 113699 172961 113727 172989
rect 113761 172961 113789 172989
rect 129059 173147 129087 173175
rect 129121 173147 129149 173175
rect 129059 173085 129087 173113
rect 129121 173085 129149 173113
rect 129059 173023 129087 173051
rect 129121 173023 129149 173051
rect 129059 172961 129087 172989
rect 129121 172961 129149 172989
rect 144419 173147 144447 173175
rect 144481 173147 144509 173175
rect 144419 173085 144447 173113
rect 144481 173085 144509 173113
rect 144419 173023 144447 173051
rect 144481 173023 144509 173051
rect 144419 172961 144447 172989
rect 144481 172961 144509 172989
rect 154625 173147 154653 173175
rect 154687 173147 154715 173175
rect 154749 173147 154777 173175
rect 154811 173147 154839 173175
rect 154625 173085 154653 173113
rect 154687 173085 154715 173113
rect 154749 173085 154777 173113
rect 154811 173085 154839 173113
rect 154625 173023 154653 173051
rect 154687 173023 154715 173051
rect 154749 173023 154777 173051
rect 154811 173023 154839 173051
rect 154625 172961 154653 172989
rect 154687 172961 154715 172989
rect 154749 172961 154777 172989
rect 154811 172961 154839 172989
rect 48485 167147 48513 167175
rect 48547 167147 48575 167175
rect 48609 167147 48637 167175
rect 48671 167147 48699 167175
rect 48485 167085 48513 167113
rect 48547 167085 48575 167113
rect 48609 167085 48637 167113
rect 48671 167085 48699 167113
rect 48485 167023 48513 167051
rect 48547 167023 48575 167051
rect 48609 167023 48637 167051
rect 48671 167023 48699 167051
rect 48485 166961 48513 166989
rect 48547 166961 48575 166989
rect 48609 166961 48637 166989
rect 48671 166961 48699 166989
rect 59939 167147 59967 167175
rect 60001 167147 60029 167175
rect 59939 167085 59967 167113
rect 60001 167085 60029 167113
rect 59939 167023 59967 167051
rect 60001 167023 60029 167051
rect 59939 166961 59967 166989
rect 60001 166961 60029 166989
rect 75299 167147 75327 167175
rect 75361 167147 75389 167175
rect 75299 167085 75327 167113
rect 75361 167085 75389 167113
rect 75299 167023 75327 167051
rect 75361 167023 75389 167051
rect 75299 166961 75327 166989
rect 75361 166961 75389 166989
rect 90659 167147 90687 167175
rect 90721 167147 90749 167175
rect 90659 167085 90687 167113
rect 90721 167085 90749 167113
rect 90659 167023 90687 167051
rect 90721 167023 90749 167051
rect 90659 166961 90687 166989
rect 90721 166961 90749 166989
rect 106019 167147 106047 167175
rect 106081 167147 106109 167175
rect 106019 167085 106047 167113
rect 106081 167085 106109 167113
rect 106019 167023 106047 167051
rect 106081 167023 106109 167051
rect 106019 166961 106047 166989
rect 106081 166961 106109 166989
rect 121379 167147 121407 167175
rect 121441 167147 121469 167175
rect 121379 167085 121407 167113
rect 121441 167085 121469 167113
rect 121379 167023 121407 167051
rect 121441 167023 121469 167051
rect 121379 166961 121407 166989
rect 121441 166961 121469 166989
rect 136739 167147 136767 167175
rect 136801 167147 136829 167175
rect 136739 167085 136767 167113
rect 136801 167085 136829 167113
rect 136739 167023 136767 167051
rect 136801 167023 136829 167051
rect 136739 166961 136767 166989
rect 136801 166961 136829 166989
rect 52259 164147 52287 164175
rect 52321 164147 52349 164175
rect 52259 164085 52287 164113
rect 52321 164085 52349 164113
rect 52259 164023 52287 164051
rect 52321 164023 52349 164051
rect 52259 163961 52287 163989
rect 52321 163961 52349 163989
rect 67619 164147 67647 164175
rect 67681 164147 67709 164175
rect 67619 164085 67647 164113
rect 67681 164085 67709 164113
rect 67619 164023 67647 164051
rect 67681 164023 67709 164051
rect 67619 163961 67647 163989
rect 67681 163961 67709 163989
rect 82979 164147 83007 164175
rect 83041 164147 83069 164175
rect 82979 164085 83007 164113
rect 83041 164085 83069 164113
rect 82979 164023 83007 164051
rect 83041 164023 83069 164051
rect 82979 163961 83007 163989
rect 83041 163961 83069 163989
rect 98339 164147 98367 164175
rect 98401 164147 98429 164175
rect 98339 164085 98367 164113
rect 98401 164085 98429 164113
rect 98339 164023 98367 164051
rect 98401 164023 98429 164051
rect 98339 163961 98367 163989
rect 98401 163961 98429 163989
rect 113699 164147 113727 164175
rect 113761 164147 113789 164175
rect 113699 164085 113727 164113
rect 113761 164085 113789 164113
rect 113699 164023 113727 164051
rect 113761 164023 113789 164051
rect 113699 163961 113727 163989
rect 113761 163961 113789 163989
rect 129059 164147 129087 164175
rect 129121 164147 129149 164175
rect 129059 164085 129087 164113
rect 129121 164085 129149 164113
rect 129059 164023 129087 164051
rect 129121 164023 129149 164051
rect 129059 163961 129087 163989
rect 129121 163961 129149 163989
rect 144419 164147 144447 164175
rect 144481 164147 144509 164175
rect 144419 164085 144447 164113
rect 144481 164085 144509 164113
rect 144419 164023 144447 164051
rect 144481 164023 144509 164051
rect 144419 163961 144447 163989
rect 144481 163961 144509 163989
rect 154625 164147 154653 164175
rect 154687 164147 154715 164175
rect 154749 164147 154777 164175
rect 154811 164147 154839 164175
rect 154625 164085 154653 164113
rect 154687 164085 154715 164113
rect 154749 164085 154777 164113
rect 154811 164085 154839 164113
rect 154625 164023 154653 164051
rect 154687 164023 154715 164051
rect 154749 164023 154777 164051
rect 154811 164023 154839 164051
rect 154625 163961 154653 163989
rect 154687 163961 154715 163989
rect 154749 163961 154777 163989
rect 154811 163961 154839 163989
rect 48485 158147 48513 158175
rect 48547 158147 48575 158175
rect 48609 158147 48637 158175
rect 48671 158147 48699 158175
rect 48485 158085 48513 158113
rect 48547 158085 48575 158113
rect 48609 158085 48637 158113
rect 48671 158085 48699 158113
rect 48485 158023 48513 158051
rect 48547 158023 48575 158051
rect 48609 158023 48637 158051
rect 48671 158023 48699 158051
rect 48485 157961 48513 157989
rect 48547 157961 48575 157989
rect 48609 157961 48637 157989
rect 48671 157961 48699 157989
rect 59939 158147 59967 158175
rect 60001 158147 60029 158175
rect 59939 158085 59967 158113
rect 60001 158085 60029 158113
rect 59939 158023 59967 158051
rect 60001 158023 60029 158051
rect 59939 157961 59967 157989
rect 60001 157961 60029 157989
rect 75299 158147 75327 158175
rect 75361 158147 75389 158175
rect 75299 158085 75327 158113
rect 75361 158085 75389 158113
rect 75299 158023 75327 158051
rect 75361 158023 75389 158051
rect 75299 157961 75327 157989
rect 75361 157961 75389 157989
rect 90659 158147 90687 158175
rect 90721 158147 90749 158175
rect 90659 158085 90687 158113
rect 90721 158085 90749 158113
rect 90659 158023 90687 158051
rect 90721 158023 90749 158051
rect 90659 157961 90687 157989
rect 90721 157961 90749 157989
rect 106019 158147 106047 158175
rect 106081 158147 106109 158175
rect 106019 158085 106047 158113
rect 106081 158085 106109 158113
rect 106019 158023 106047 158051
rect 106081 158023 106109 158051
rect 106019 157961 106047 157989
rect 106081 157961 106109 157989
rect 121379 158147 121407 158175
rect 121441 158147 121469 158175
rect 121379 158085 121407 158113
rect 121441 158085 121469 158113
rect 121379 158023 121407 158051
rect 121441 158023 121469 158051
rect 121379 157961 121407 157989
rect 121441 157961 121469 157989
rect 136739 158147 136767 158175
rect 136801 158147 136829 158175
rect 136739 158085 136767 158113
rect 136801 158085 136829 158113
rect 136739 158023 136767 158051
rect 136801 158023 136829 158051
rect 136739 157961 136767 157989
rect 136801 157961 136829 157989
rect 52259 155147 52287 155175
rect 52321 155147 52349 155175
rect 52259 155085 52287 155113
rect 52321 155085 52349 155113
rect 52259 155023 52287 155051
rect 52321 155023 52349 155051
rect 52259 154961 52287 154989
rect 52321 154961 52349 154989
rect 67619 155147 67647 155175
rect 67681 155147 67709 155175
rect 67619 155085 67647 155113
rect 67681 155085 67709 155113
rect 67619 155023 67647 155051
rect 67681 155023 67709 155051
rect 67619 154961 67647 154989
rect 67681 154961 67709 154989
rect 82979 155147 83007 155175
rect 83041 155147 83069 155175
rect 82979 155085 83007 155113
rect 83041 155085 83069 155113
rect 82979 155023 83007 155051
rect 83041 155023 83069 155051
rect 82979 154961 83007 154989
rect 83041 154961 83069 154989
rect 98339 155147 98367 155175
rect 98401 155147 98429 155175
rect 98339 155085 98367 155113
rect 98401 155085 98429 155113
rect 98339 155023 98367 155051
rect 98401 155023 98429 155051
rect 98339 154961 98367 154989
rect 98401 154961 98429 154989
rect 113699 155147 113727 155175
rect 113761 155147 113789 155175
rect 113699 155085 113727 155113
rect 113761 155085 113789 155113
rect 113699 155023 113727 155051
rect 113761 155023 113789 155051
rect 113699 154961 113727 154989
rect 113761 154961 113789 154989
rect 129059 155147 129087 155175
rect 129121 155147 129149 155175
rect 129059 155085 129087 155113
rect 129121 155085 129149 155113
rect 129059 155023 129087 155051
rect 129121 155023 129149 155051
rect 129059 154961 129087 154989
rect 129121 154961 129149 154989
rect 144419 155147 144447 155175
rect 144481 155147 144509 155175
rect 144419 155085 144447 155113
rect 144481 155085 144509 155113
rect 144419 155023 144447 155051
rect 144481 155023 144509 155051
rect 144419 154961 144447 154989
rect 144481 154961 144509 154989
rect 154625 155147 154653 155175
rect 154687 155147 154715 155175
rect 154749 155147 154777 155175
rect 154811 155147 154839 155175
rect 154625 155085 154653 155113
rect 154687 155085 154715 155113
rect 154749 155085 154777 155113
rect 154811 155085 154839 155113
rect 154625 155023 154653 155051
rect 154687 155023 154715 155051
rect 154749 155023 154777 155051
rect 154811 155023 154839 155051
rect 154625 154961 154653 154989
rect 154687 154961 154715 154989
rect 154749 154961 154777 154989
rect 154811 154961 154839 154989
rect 48485 149147 48513 149175
rect 48547 149147 48575 149175
rect 48609 149147 48637 149175
rect 48671 149147 48699 149175
rect 48485 149085 48513 149113
rect 48547 149085 48575 149113
rect 48609 149085 48637 149113
rect 48671 149085 48699 149113
rect 48485 149023 48513 149051
rect 48547 149023 48575 149051
rect 48609 149023 48637 149051
rect 48671 149023 48699 149051
rect 48485 148961 48513 148989
rect 48547 148961 48575 148989
rect 48609 148961 48637 148989
rect 48671 148961 48699 148989
rect 59939 149147 59967 149175
rect 60001 149147 60029 149175
rect 59939 149085 59967 149113
rect 60001 149085 60029 149113
rect 59939 149023 59967 149051
rect 60001 149023 60029 149051
rect 59939 148961 59967 148989
rect 60001 148961 60029 148989
rect 75299 149147 75327 149175
rect 75361 149147 75389 149175
rect 75299 149085 75327 149113
rect 75361 149085 75389 149113
rect 75299 149023 75327 149051
rect 75361 149023 75389 149051
rect 75299 148961 75327 148989
rect 75361 148961 75389 148989
rect 90659 149147 90687 149175
rect 90721 149147 90749 149175
rect 90659 149085 90687 149113
rect 90721 149085 90749 149113
rect 90659 149023 90687 149051
rect 90721 149023 90749 149051
rect 90659 148961 90687 148989
rect 90721 148961 90749 148989
rect 106019 149147 106047 149175
rect 106081 149147 106109 149175
rect 106019 149085 106047 149113
rect 106081 149085 106109 149113
rect 106019 149023 106047 149051
rect 106081 149023 106109 149051
rect 106019 148961 106047 148989
rect 106081 148961 106109 148989
rect 121379 149147 121407 149175
rect 121441 149147 121469 149175
rect 121379 149085 121407 149113
rect 121441 149085 121469 149113
rect 121379 149023 121407 149051
rect 121441 149023 121469 149051
rect 121379 148961 121407 148989
rect 121441 148961 121469 148989
rect 136739 149147 136767 149175
rect 136801 149147 136829 149175
rect 136739 149085 136767 149113
rect 136801 149085 136829 149113
rect 136739 149023 136767 149051
rect 136801 149023 136829 149051
rect 136739 148961 136767 148989
rect 136801 148961 136829 148989
rect 52259 146147 52287 146175
rect 52321 146147 52349 146175
rect 52259 146085 52287 146113
rect 52321 146085 52349 146113
rect 52259 146023 52287 146051
rect 52321 146023 52349 146051
rect 52259 145961 52287 145989
rect 52321 145961 52349 145989
rect 67619 146147 67647 146175
rect 67681 146147 67709 146175
rect 67619 146085 67647 146113
rect 67681 146085 67709 146113
rect 67619 146023 67647 146051
rect 67681 146023 67709 146051
rect 67619 145961 67647 145989
rect 67681 145961 67709 145989
rect 82979 146147 83007 146175
rect 83041 146147 83069 146175
rect 82979 146085 83007 146113
rect 83041 146085 83069 146113
rect 82979 146023 83007 146051
rect 83041 146023 83069 146051
rect 82979 145961 83007 145989
rect 83041 145961 83069 145989
rect 98339 146147 98367 146175
rect 98401 146147 98429 146175
rect 98339 146085 98367 146113
rect 98401 146085 98429 146113
rect 98339 146023 98367 146051
rect 98401 146023 98429 146051
rect 98339 145961 98367 145989
rect 98401 145961 98429 145989
rect 113699 146147 113727 146175
rect 113761 146147 113789 146175
rect 113699 146085 113727 146113
rect 113761 146085 113789 146113
rect 113699 146023 113727 146051
rect 113761 146023 113789 146051
rect 113699 145961 113727 145989
rect 113761 145961 113789 145989
rect 129059 146147 129087 146175
rect 129121 146147 129149 146175
rect 129059 146085 129087 146113
rect 129121 146085 129149 146113
rect 129059 146023 129087 146051
rect 129121 146023 129149 146051
rect 129059 145961 129087 145989
rect 129121 145961 129149 145989
rect 144419 146147 144447 146175
rect 144481 146147 144509 146175
rect 144419 146085 144447 146113
rect 144481 146085 144509 146113
rect 144419 146023 144447 146051
rect 144481 146023 144509 146051
rect 144419 145961 144447 145989
rect 144481 145961 144509 145989
rect 154625 146147 154653 146175
rect 154687 146147 154715 146175
rect 154749 146147 154777 146175
rect 154811 146147 154839 146175
rect 154625 146085 154653 146113
rect 154687 146085 154715 146113
rect 154749 146085 154777 146113
rect 154811 146085 154839 146113
rect 154625 146023 154653 146051
rect 154687 146023 154715 146051
rect 154749 146023 154777 146051
rect 154811 146023 154839 146051
rect 154625 145961 154653 145989
rect 154687 145961 154715 145989
rect 154749 145961 154777 145989
rect 154811 145961 154839 145989
rect 48485 140147 48513 140175
rect 48547 140147 48575 140175
rect 48609 140147 48637 140175
rect 48671 140147 48699 140175
rect 48485 140085 48513 140113
rect 48547 140085 48575 140113
rect 48609 140085 48637 140113
rect 48671 140085 48699 140113
rect 48485 140023 48513 140051
rect 48547 140023 48575 140051
rect 48609 140023 48637 140051
rect 48671 140023 48699 140051
rect 48485 139961 48513 139989
rect 48547 139961 48575 139989
rect 48609 139961 48637 139989
rect 48671 139961 48699 139989
rect 59939 140147 59967 140175
rect 60001 140147 60029 140175
rect 59939 140085 59967 140113
rect 60001 140085 60029 140113
rect 59939 140023 59967 140051
rect 60001 140023 60029 140051
rect 59939 139961 59967 139989
rect 60001 139961 60029 139989
rect 75299 140147 75327 140175
rect 75361 140147 75389 140175
rect 75299 140085 75327 140113
rect 75361 140085 75389 140113
rect 75299 140023 75327 140051
rect 75361 140023 75389 140051
rect 75299 139961 75327 139989
rect 75361 139961 75389 139989
rect 90659 140147 90687 140175
rect 90721 140147 90749 140175
rect 90659 140085 90687 140113
rect 90721 140085 90749 140113
rect 90659 140023 90687 140051
rect 90721 140023 90749 140051
rect 90659 139961 90687 139989
rect 90721 139961 90749 139989
rect 106019 140147 106047 140175
rect 106081 140147 106109 140175
rect 106019 140085 106047 140113
rect 106081 140085 106109 140113
rect 106019 140023 106047 140051
rect 106081 140023 106109 140051
rect 106019 139961 106047 139989
rect 106081 139961 106109 139989
rect 121379 140147 121407 140175
rect 121441 140147 121469 140175
rect 121379 140085 121407 140113
rect 121441 140085 121469 140113
rect 121379 140023 121407 140051
rect 121441 140023 121469 140051
rect 121379 139961 121407 139989
rect 121441 139961 121469 139989
rect 136739 140147 136767 140175
rect 136801 140147 136829 140175
rect 136739 140085 136767 140113
rect 136801 140085 136829 140113
rect 136739 140023 136767 140051
rect 136801 140023 136829 140051
rect 136739 139961 136767 139989
rect 136801 139961 136829 139989
rect 52259 137147 52287 137175
rect 52321 137147 52349 137175
rect 52259 137085 52287 137113
rect 52321 137085 52349 137113
rect 52259 137023 52287 137051
rect 52321 137023 52349 137051
rect 52259 136961 52287 136989
rect 52321 136961 52349 136989
rect 67619 137147 67647 137175
rect 67681 137147 67709 137175
rect 67619 137085 67647 137113
rect 67681 137085 67709 137113
rect 67619 137023 67647 137051
rect 67681 137023 67709 137051
rect 67619 136961 67647 136989
rect 67681 136961 67709 136989
rect 82979 137147 83007 137175
rect 83041 137147 83069 137175
rect 82979 137085 83007 137113
rect 83041 137085 83069 137113
rect 82979 137023 83007 137051
rect 83041 137023 83069 137051
rect 82979 136961 83007 136989
rect 83041 136961 83069 136989
rect 98339 137147 98367 137175
rect 98401 137147 98429 137175
rect 98339 137085 98367 137113
rect 98401 137085 98429 137113
rect 98339 137023 98367 137051
rect 98401 137023 98429 137051
rect 98339 136961 98367 136989
rect 98401 136961 98429 136989
rect 113699 137147 113727 137175
rect 113761 137147 113789 137175
rect 113699 137085 113727 137113
rect 113761 137085 113789 137113
rect 113699 137023 113727 137051
rect 113761 137023 113789 137051
rect 113699 136961 113727 136989
rect 113761 136961 113789 136989
rect 129059 137147 129087 137175
rect 129121 137147 129149 137175
rect 129059 137085 129087 137113
rect 129121 137085 129149 137113
rect 129059 137023 129087 137051
rect 129121 137023 129149 137051
rect 129059 136961 129087 136989
rect 129121 136961 129149 136989
rect 144419 137147 144447 137175
rect 144481 137147 144509 137175
rect 144419 137085 144447 137113
rect 144481 137085 144509 137113
rect 144419 137023 144447 137051
rect 144481 137023 144509 137051
rect 144419 136961 144447 136989
rect 144481 136961 144509 136989
rect 154625 137147 154653 137175
rect 154687 137147 154715 137175
rect 154749 137147 154777 137175
rect 154811 137147 154839 137175
rect 154625 137085 154653 137113
rect 154687 137085 154715 137113
rect 154749 137085 154777 137113
rect 154811 137085 154839 137113
rect 154625 137023 154653 137051
rect 154687 137023 154715 137051
rect 154749 137023 154777 137051
rect 154811 137023 154839 137051
rect 154625 136961 154653 136989
rect 154687 136961 154715 136989
rect 154749 136961 154777 136989
rect 154811 136961 154839 136989
rect 48485 131147 48513 131175
rect 48547 131147 48575 131175
rect 48609 131147 48637 131175
rect 48671 131147 48699 131175
rect 48485 131085 48513 131113
rect 48547 131085 48575 131113
rect 48609 131085 48637 131113
rect 48671 131085 48699 131113
rect 48485 131023 48513 131051
rect 48547 131023 48575 131051
rect 48609 131023 48637 131051
rect 48671 131023 48699 131051
rect 48485 130961 48513 130989
rect 48547 130961 48575 130989
rect 48609 130961 48637 130989
rect 48671 130961 48699 130989
rect 59939 131147 59967 131175
rect 60001 131147 60029 131175
rect 59939 131085 59967 131113
rect 60001 131085 60029 131113
rect 59939 131023 59967 131051
rect 60001 131023 60029 131051
rect 59939 130961 59967 130989
rect 60001 130961 60029 130989
rect 75299 131147 75327 131175
rect 75361 131147 75389 131175
rect 75299 131085 75327 131113
rect 75361 131085 75389 131113
rect 75299 131023 75327 131051
rect 75361 131023 75389 131051
rect 75299 130961 75327 130989
rect 75361 130961 75389 130989
rect 90659 131147 90687 131175
rect 90721 131147 90749 131175
rect 90659 131085 90687 131113
rect 90721 131085 90749 131113
rect 90659 131023 90687 131051
rect 90721 131023 90749 131051
rect 90659 130961 90687 130989
rect 90721 130961 90749 130989
rect 106019 131147 106047 131175
rect 106081 131147 106109 131175
rect 106019 131085 106047 131113
rect 106081 131085 106109 131113
rect 106019 131023 106047 131051
rect 106081 131023 106109 131051
rect 106019 130961 106047 130989
rect 106081 130961 106109 130989
rect 121379 131147 121407 131175
rect 121441 131147 121469 131175
rect 121379 131085 121407 131113
rect 121441 131085 121469 131113
rect 121379 131023 121407 131051
rect 121441 131023 121469 131051
rect 121379 130961 121407 130989
rect 121441 130961 121469 130989
rect 136739 131147 136767 131175
rect 136801 131147 136829 131175
rect 136739 131085 136767 131113
rect 136801 131085 136829 131113
rect 136739 131023 136767 131051
rect 136801 131023 136829 131051
rect 136739 130961 136767 130989
rect 136801 130961 136829 130989
rect 52259 128147 52287 128175
rect 52321 128147 52349 128175
rect 52259 128085 52287 128113
rect 52321 128085 52349 128113
rect 52259 128023 52287 128051
rect 52321 128023 52349 128051
rect 52259 127961 52287 127989
rect 52321 127961 52349 127989
rect 67619 128147 67647 128175
rect 67681 128147 67709 128175
rect 67619 128085 67647 128113
rect 67681 128085 67709 128113
rect 67619 128023 67647 128051
rect 67681 128023 67709 128051
rect 67619 127961 67647 127989
rect 67681 127961 67709 127989
rect 82979 128147 83007 128175
rect 83041 128147 83069 128175
rect 82979 128085 83007 128113
rect 83041 128085 83069 128113
rect 82979 128023 83007 128051
rect 83041 128023 83069 128051
rect 82979 127961 83007 127989
rect 83041 127961 83069 127989
rect 98339 128147 98367 128175
rect 98401 128147 98429 128175
rect 98339 128085 98367 128113
rect 98401 128085 98429 128113
rect 98339 128023 98367 128051
rect 98401 128023 98429 128051
rect 98339 127961 98367 127989
rect 98401 127961 98429 127989
rect 113699 128147 113727 128175
rect 113761 128147 113789 128175
rect 113699 128085 113727 128113
rect 113761 128085 113789 128113
rect 113699 128023 113727 128051
rect 113761 128023 113789 128051
rect 113699 127961 113727 127989
rect 113761 127961 113789 127989
rect 129059 128147 129087 128175
rect 129121 128147 129149 128175
rect 129059 128085 129087 128113
rect 129121 128085 129149 128113
rect 129059 128023 129087 128051
rect 129121 128023 129149 128051
rect 129059 127961 129087 127989
rect 129121 127961 129149 127989
rect 144419 128147 144447 128175
rect 144481 128147 144509 128175
rect 144419 128085 144447 128113
rect 144481 128085 144509 128113
rect 144419 128023 144447 128051
rect 144481 128023 144509 128051
rect 144419 127961 144447 127989
rect 144481 127961 144509 127989
rect 154625 128147 154653 128175
rect 154687 128147 154715 128175
rect 154749 128147 154777 128175
rect 154811 128147 154839 128175
rect 154625 128085 154653 128113
rect 154687 128085 154715 128113
rect 154749 128085 154777 128113
rect 154811 128085 154839 128113
rect 154625 128023 154653 128051
rect 154687 128023 154715 128051
rect 154749 128023 154777 128051
rect 154811 128023 154839 128051
rect 154625 127961 154653 127989
rect 154687 127961 154715 127989
rect 154749 127961 154777 127989
rect 154811 127961 154839 127989
rect 48485 122147 48513 122175
rect 48547 122147 48575 122175
rect 48609 122147 48637 122175
rect 48671 122147 48699 122175
rect 48485 122085 48513 122113
rect 48547 122085 48575 122113
rect 48609 122085 48637 122113
rect 48671 122085 48699 122113
rect 48485 122023 48513 122051
rect 48547 122023 48575 122051
rect 48609 122023 48637 122051
rect 48671 122023 48699 122051
rect 48485 121961 48513 121989
rect 48547 121961 48575 121989
rect 48609 121961 48637 121989
rect 48671 121961 48699 121989
rect 48485 113147 48513 113175
rect 48547 113147 48575 113175
rect 48609 113147 48637 113175
rect 48671 113147 48699 113175
rect 48485 113085 48513 113113
rect 48547 113085 48575 113113
rect 48609 113085 48637 113113
rect 48671 113085 48699 113113
rect 48485 113023 48513 113051
rect 48547 113023 48575 113051
rect 48609 113023 48637 113051
rect 48671 113023 48699 113051
rect 48485 112961 48513 112989
rect 48547 112961 48575 112989
rect 48609 112961 48637 112989
rect 48671 112961 48699 112989
rect 55625 119147 55653 119175
rect 55687 119147 55715 119175
rect 55749 119147 55777 119175
rect 55811 119147 55839 119175
rect 55625 119085 55653 119113
rect 55687 119085 55715 119113
rect 55749 119085 55777 119113
rect 55811 119085 55839 119113
rect 55625 119023 55653 119051
rect 55687 119023 55715 119051
rect 55749 119023 55777 119051
rect 55811 119023 55839 119051
rect 55625 118961 55653 118989
rect 55687 118961 55715 118989
rect 55749 118961 55777 118989
rect 55811 118961 55839 118989
rect 55625 110147 55653 110175
rect 55687 110147 55715 110175
rect 55749 110147 55777 110175
rect 55811 110147 55839 110175
rect 55625 110085 55653 110113
rect 55687 110085 55715 110113
rect 55749 110085 55777 110113
rect 55811 110085 55839 110113
rect 55625 110023 55653 110051
rect 55687 110023 55715 110051
rect 55749 110023 55777 110051
rect 55811 110023 55839 110051
rect 55625 109961 55653 109989
rect 55687 109961 55715 109989
rect 55749 109961 55777 109989
rect 55811 109961 55839 109989
rect 48485 104147 48513 104175
rect 48547 104147 48575 104175
rect 48609 104147 48637 104175
rect 48671 104147 48699 104175
rect 48485 104085 48513 104113
rect 48547 104085 48575 104113
rect 48609 104085 48637 104113
rect 48671 104085 48699 104113
rect 48485 104023 48513 104051
rect 48547 104023 48575 104051
rect 48609 104023 48637 104051
rect 48671 104023 48699 104051
rect 48485 103961 48513 103989
rect 48547 103961 48575 103989
rect 48609 103961 48637 103989
rect 48671 103961 48699 103989
rect 54509 104147 54537 104175
rect 54571 104147 54599 104175
rect 54509 104085 54537 104113
rect 54571 104085 54599 104113
rect 54509 104023 54537 104051
rect 54571 104023 54599 104051
rect 54509 103961 54537 103989
rect 54571 103961 54599 103989
rect 52259 101147 52287 101175
rect 52321 101147 52349 101175
rect 52259 101085 52287 101113
rect 52321 101085 52349 101113
rect 52259 101023 52287 101051
rect 52321 101023 52349 101051
rect 52259 100961 52287 100989
rect 52321 100961 52349 100989
rect 57485 122147 57513 122175
rect 57547 122147 57575 122175
rect 57609 122147 57637 122175
rect 57671 122147 57699 122175
rect 57485 122085 57513 122113
rect 57547 122085 57575 122113
rect 57609 122085 57637 122113
rect 57671 122085 57699 122113
rect 57485 122023 57513 122051
rect 57547 122023 57575 122051
rect 57609 122023 57637 122051
rect 57671 122023 57699 122051
rect 57485 121961 57513 121989
rect 57547 121961 57575 121989
rect 57609 121961 57637 121989
rect 57671 121961 57699 121989
rect 57485 113147 57513 113175
rect 57547 113147 57575 113175
rect 57609 113147 57637 113175
rect 57671 113147 57699 113175
rect 57485 113085 57513 113113
rect 57547 113085 57575 113113
rect 57609 113085 57637 113113
rect 57671 113085 57699 113113
rect 57485 113023 57513 113051
rect 57547 113023 57575 113051
rect 57609 113023 57637 113051
rect 57671 113023 57699 113051
rect 57485 112961 57513 112989
rect 57547 112961 57575 112989
rect 57609 112961 57637 112989
rect 57671 112961 57699 112989
rect 64625 119147 64653 119175
rect 64687 119147 64715 119175
rect 64749 119147 64777 119175
rect 64811 119147 64839 119175
rect 64625 119085 64653 119113
rect 64687 119085 64715 119113
rect 64749 119085 64777 119113
rect 64811 119085 64839 119113
rect 64625 119023 64653 119051
rect 64687 119023 64715 119051
rect 64749 119023 64777 119051
rect 64811 119023 64839 119051
rect 64625 118961 64653 118989
rect 64687 118961 64715 118989
rect 64749 118961 64777 118989
rect 64811 118961 64839 118989
rect 64625 110147 64653 110175
rect 64687 110147 64715 110175
rect 64749 110147 64777 110175
rect 64811 110147 64839 110175
rect 64625 110085 64653 110113
rect 64687 110085 64715 110113
rect 64749 110085 64777 110113
rect 64811 110085 64839 110113
rect 64625 110023 64653 110051
rect 64687 110023 64715 110051
rect 64749 110023 64777 110051
rect 64811 110023 64839 110051
rect 64625 109961 64653 109989
rect 64687 109961 64715 109989
rect 64749 109961 64777 109989
rect 64811 109961 64839 109989
rect 57485 104147 57513 104175
rect 57547 104147 57575 104175
rect 57609 104147 57637 104175
rect 57671 104147 57699 104175
rect 57485 104085 57513 104113
rect 57547 104085 57575 104113
rect 57609 104085 57637 104113
rect 57671 104085 57699 104113
rect 57485 104023 57513 104051
rect 57547 104023 57575 104051
rect 57609 104023 57637 104051
rect 57671 104023 57699 104051
rect 57485 103961 57513 103989
rect 57547 103961 57575 103989
rect 57609 103961 57637 103989
rect 57671 103961 57699 103989
rect 55625 101147 55653 101175
rect 55687 101147 55715 101175
rect 55749 101147 55777 101175
rect 55811 101147 55839 101175
rect 55625 101085 55653 101113
rect 55687 101085 55715 101113
rect 55749 101085 55777 101113
rect 55811 101085 55839 101113
rect 55625 101023 55653 101051
rect 55687 101023 55715 101051
rect 55749 101023 55777 101051
rect 55811 101023 55839 101051
rect 55625 100961 55653 100989
rect 55687 100961 55715 100989
rect 55749 100961 55777 100989
rect 55811 100961 55839 100989
rect 48485 95147 48513 95175
rect 48547 95147 48575 95175
rect 48609 95147 48637 95175
rect 48671 95147 48699 95175
rect 48485 95085 48513 95113
rect 48547 95085 48575 95113
rect 48609 95085 48637 95113
rect 48671 95085 48699 95113
rect 48485 95023 48513 95051
rect 48547 95023 48575 95051
rect 48609 95023 48637 95051
rect 48671 95023 48699 95051
rect 48485 94961 48513 94989
rect 48547 94961 48575 94989
rect 48609 94961 48637 94989
rect 48671 94961 48699 94989
rect 54509 95147 54537 95175
rect 54571 95147 54599 95175
rect 54509 95085 54537 95113
rect 54571 95085 54599 95113
rect 54509 95023 54537 95051
rect 54571 95023 54599 95051
rect 54509 94961 54537 94989
rect 54571 94961 54599 94989
rect 52259 92147 52287 92175
rect 52321 92147 52349 92175
rect 52259 92085 52287 92113
rect 52321 92085 52349 92113
rect 52259 92023 52287 92051
rect 52321 92023 52349 92051
rect 52259 91961 52287 91989
rect 52321 91961 52349 91989
rect 56759 101147 56787 101175
rect 56821 101147 56849 101175
rect 56759 101085 56787 101113
rect 56821 101085 56849 101113
rect 56759 101023 56787 101051
rect 56821 101023 56849 101051
rect 56759 100961 56787 100989
rect 56821 100961 56849 100989
rect 59009 104147 59037 104175
rect 59071 104147 59099 104175
rect 59009 104085 59037 104113
rect 59071 104085 59099 104113
rect 59009 104023 59037 104051
rect 59071 104023 59099 104051
rect 59009 103961 59037 103989
rect 59071 103961 59099 103989
rect 63509 104147 63537 104175
rect 63571 104147 63599 104175
rect 63509 104085 63537 104113
rect 63571 104085 63599 104113
rect 63509 104023 63537 104051
rect 63571 104023 63599 104051
rect 63509 103961 63537 103989
rect 63571 103961 63599 103989
rect 61259 101147 61287 101175
rect 61321 101147 61349 101175
rect 61259 101085 61287 101113
rect 61321 101085 61349 101113
rect 61259 101023 61287 101051
rect 61321 101023 61349 101051
rect 61259 100961 61287 100989
rect 61321 100961 61349 100989
rect 66485 122147 66513 122175
rect 66547 122147 66575 122175
rect 66609 122147 66637 122175
rect 66671 122147 66699 122175
rect 66485 122085 66513 122113
rect 66547 122085 66575 122113
rect 66609 122085 66637 122113
rect 66671 122085 66699 122113
rect 66485 122023 66513 122051
rect 66547 122023 66575 122051
rect 66609 122023 66637 122051
rect 66671 122023 66699 122051
rect 66485 121961 66513 121989
rect 66547 121961 66575 121989
rect 66609 121961 66637 121989
rect 66671 121961 66699 121989
rect 66485 113147 66513 113175
rect 66547 113147 66575 113175
rect 66609 113147 66637 113175
rect 66671 113147 66699 113175
rect 66485 113085 66513 113113
rect 66547 113085 66575 113113
rect 66609 113085 66637 113113
rect 66671 113085 66699 113113
rect 66485 113023 66513 113051
rect 66547 113023 66575 113051
rect 66609 113023 66637 113051
rect 66671 113023 66699 113051
rect 66485 112961 66513 112989
rect 66547 112961 66575 112989
rect 66609 112961 66637 112989
rect 66671 112961 66699 112989
rect 73625 119147 73653 119175
rect 73687 119147 73715 119175
rect 73749 119147 73777 119175
rect 73811 119147 73839 119175
rect 73625 119085 73653 119113
rect 73687 119085 73715 119113
rect 73749 119085 73777 119113
rect 73811 119085 73839 119113
rect 73625 119023 73653 119051
rect 73687 119023 73715 119051
rect 73749 119023 73777 119051
rect 73811 119023 73839 119051
rect 73625 118961 73653 118989
rect 73687 118961 73715 118989
rect 73749 118961 73777 118989
rect 73811 118961 73839 118989
rect 73625 110147 73653 110175
rect 73687 110147 73715 110175
rect 73749 110147 73777 110175
rect 73811 110147 73839 110175
rect 73625 110085 73653 110113
rect 73687 110085 73715 110113
rect 73749 110085 73777 110113
rect 73811 110085 73839 110113
rect 73625 110023 73653 110051
rect 73687 110023 73715 110051
rect 73749 110023 73777 110051
rect 73811 110023 73839 110051
rect 73625 109961 73653 109989
rect 73687 109961 73715 109989
rect 73749 109961 73777 109989
rect 73811 109961 73839 109989
rect 66485 104147 66513 104175
rect 66547 104147 66575 104175
rect 66609 104147 66637 104175
rect 66671 104147 66699 104175
rect 66485 104085 66513 104113
rect 66547 104085 66575 104113
rect 66609 104085 66637 104113
rect 66671 104085 66699 104113
rect 66485 104023 66513 104051
rect 66547 104023 66575 104051
rect 66609 104023 66637 104051
rect 66671 104023 66699 104051
rect 66485 103961 66513 103989
rect 66547 103961 66575 103989
rect 66609 103961 66637 103989
rect 66671 103961 66699 103989
rect 64625 101147 64653 101175
rect 64687 101147 64715 101175
rect 64749 101147 64777 101175
rect 64811 101147 64839 101175
rect 64625 101085 64653 101113
rect 64687 101085 64715 101113
rect 64749 101085 64777 101113
rect 64811 101085 64839 101113
rect 64625 101023 64653 101051
rect 64687 101023 64715 101051
rect 64749 101023 64777 101051
rect 64811 101023 64839 101051
rect 64625 100961 64653 100989
rect 64687 100961 64715 100989
rect 64749 100961 64777 100989
rect 64811 100961 64839 100989
rect 57485 95147 57513 95175
rect 57547 95147 57575 95175
rect 57609 95147 57637 95175
rect 57671 95147 57699 95175
rect 57485 95085 57513 95113
rect 57547 95085 57575 95113
rect 57609 95085 57637 95113
rect 57671 95085 57699 95113
rect 57485 95023 57513 95051
rect 57547 95023 57575 95051
rect 57609 95023 57637 95051
rect 57671 95023 57699 95051
rect 57485 94961 57513 94989
rect 57547 94961 57575 94989
rect 57609 94961 57637 94989
rect 57671 94961 57699 94989
rect 55625 92147 55653 92175
rect 55687 92147 55715 92175
rect 55749 92147 55777 92175
rect 55811 92147 55839 92175
rect 55625 92085 55653 92113
rect 55687 92085 55715 92113
rect 55749 92085 55777 92113
rect 55811 92085 55839 92113
rect 55625 92023 55653 92051
rect 55687 92023 55715 92051
rect 55749 92023 55777 92051
rect 55811 92023 55839 92051
rect 55625 91961 55653 91989
rect 55687 91961 55715 91989
rect 55749 91961 55777 91989
rect 55811 91961 55839 91989
rect 48485 86147 48513 86175
rect 48547 86147 48575 86175
rect 48609 86147 48637 86175
rect 48671 86147 48699 86175
rect 48485 86085 48513 86113
rect 48547 86085 48575 86113
rect 48609 86085 48637 86113
rect 48671 86085 48699 86113
rect 48485 86023 48513 86051
rect 48547 86023 48575 86051
rect 48609 86023 48637 86051
rect 48671 86023 48699 86051
rect 48485 85961 48513 85989
rect 48547 85961 48575 85989
rect 48609 85961 48637 85989
rect 48671 85961 48699 85989
rect 54509 86147 54537 86175
rect 54571 86147 54599 86175
rect 54509 86085 54537 86113
rect 54571 86085 54599 86113
rect 54509 86023 54537 86051
rect 54571 86023 54599 86051
rect 54509 85961 54537 85989
rect 54571 85961 54599 85989
rect 52259 83147 52287 83175
rect 52321 83147 52349 83175
rect 52259 83085 52287 83113
rect 52321 83085 52349 83113
rect 52259 83023 52287 83051
rect 52321 83023 52349 83051
rect 52259 82961 52287 82989
rect 52321 82961 52349 82989
rect 56759 92147 56787 92175
rect 56821 92147 56849 92175
rect 56759 92085 56787 92113
rect 56821 92085 56849 92113
rect 56759 92023 56787 92051
rect 56821 92023 56849 92051
rect 56759 91961 56787 91989
rect 56821 91961 56849 91989
rect 59009 95147 59037 95175
rect 59071 95147 59099 95175
rect 59009 95085 59037 95113
rect 59071 95085 59099 95113
rect 59009 95023 59037 95051
rect 59071 95023 59099 95051
rect 59009 94961 59037 94989
rect 59071 94961 59099 94989
rect 63509 95147 63537 95175
rect 63571 95147 63599 95175
rect 63509 95085 63537 95113
rect 63571 95085 63599 95113
rect 63509 95023 63537 95051
rect 63571 95023 63599 95051
rect 63509 94961 63537 94989
rect 63571 94961 63599 94989
rect 61259 92147 61287 92175
rect 61321 92147 61349 92175
rect 61259 92085 61287 92113
rect 61321 92085 61349 92113
rect 61259 92023 61287 92051
rect 61321 92023 61349 92051
rect 61259 91961 61287 91989
rect 61321 91961 61349 91989
rect 65759 101147 65787 101175
rect 65821 101147 65849 101175
rect 65759 101085 65787 101113
rect 65821 101085 65849 101113
rect 65759 101023 65787 101051
rect 65821 101023 65849 101051
rect 65759 100961 65787 100989
rect 65821 100961 65849 100989
rect 68009 104147 68037 104175
rect 68071 104147 68099 104175
rect 68009 104085 68037 104113
rect 68071 104085 68099 104113
rect 68009 104023 68037 104051
rect 68071 104023 68099 104051
rect 68009 103961 68037 103989
rect 68071 103961 68099 103989
rect 72509 104147 72537 104175
rect 72571 104147 72599 104175
rect 72509 104085 72537 104113
rect 72571 104085 72599 104113
rect 72509 104023 72537 104051
rect 72571 104023 72599 104051
rect 72509 103961 72537 103989
rect 72571 103961 72599 103989
rect 70259 101147 70287 101175
rect 70321 101147 70349 101175
rect 70259 101085 70287 101113
rect 70321 101085 70349 101113
rect 70259 101023 70287 101051
rect 70321 101023 70349 101051
rect 70259 100961 70287 100989
rect 70321 100961 70349 100989
rect 75485 122147 75513 122175
rect 75547 122147 75575 122175
rect 75609 122147 75637 122175
rect 75671 122147 75699 122175
rect 75485 122085 75513 122113
rect 75547 122085 75575 122113
rect 75609 122085 75637 122113
rect 75671 122085 75699 122113
rect 75485 122023 75513 122051
rect 75547 122023 75575 122051
rect 75609 122023 75637 122051
rect 75671 122023 75699 122051
rect 75485 121961 75513 121989
rect 75547 121961 75575 121989
rect 75609 121961 75637 121989
rect 75671 121961 75699 121989
rect 75485 113147 75513 113175
rect 75547 113147 75575 113175
rect 75609 113147 75637 113175
rect 75671 113147 75699 113175
rect 75485 113085 75513 113113
rect 75547 113085 75575 113113
rect 75609 113085 75637 113113
rect 75671 113085 75699 113113
rect 75485 113023 75513 113051
rect 75547 113023 75575 113051
rect 75609 113023 75637 113051
rect 75671 113023 75699 113051
rect 75485 112961 75513 112989
rect 75547 112961 75575 112989
rect 75609 112961 75637 112989
rect 75671 112961 75699 112989
rect 82625 119147 82653 119175
rect 82687 119147 82715 119175
rect 82749 119147 82777 119175
rect 82811 119147 82839 119175
rect 82625 119085 82653 119113
rect 82687 119085 82715 119113
rect 82749 119085 82777 119113
rect 82811 119085 82839 119113
rect 82625 119023 82653 119051
rect 82687 119023 82715 119051
rect 82749 119023 82777 119051
rect 82811 119023 82839 119051
rect 82625 118961 82653 118989
rect 82687 118961 82715 118989
rect 82749 118961 82777 118989
rect 82811 118961 82839 118989
rect 82625 110147 82653 110175
rect 82687 110147 82715 110175
rect 82749 110147 82777 110175
rect 82811 110147 82839 110175
rect 82625 110085 82653 110113
rect 82687 110085 82715 110113
rect 82749 110085 82777 110113
rect 82811 110085 82839 110113
rect 82625 110023 82653 110051
rect 82687 110023 82715 110051
rect 82749 110023 82777 110051
rect 82811 110023 82839 110051
rect 82625 109961 82653 109989
rect 82687 109961 82715 109989
rect 82749 109961 82777 109989
rect 82811 109961 82839 109989
rect 75485 104147 75513 104175
rect 75547 104147 75575 104175
rect 75609 104147 75637 104175
rect 75671 104147 75699 104175
rect 75485 104085 75513 104113
rect 75547 104085 75575 104113
rect 75609 104085 75637 104113
rect 75671 104085 75699 104113
rect 75485 104023 75513 104051
rect 75547 104023 75575 104051
rect 75609 104023 75637 104051
rect 75671 104023 75699 104051
rect 75485 103961 75513 103989
rect 75547 103961 75575 103989
rect 75609 103961 75637 103989
rect 75671 103961 75699 103989
rect 73625 101147 73653 101175
rect 73687 101147 73715 101175
rect 73749 101147 73777 101175
rect 73811 101147 73839 101175
rect 73625 101085 73653 101113
rect 73687 101085 73715 101113
rect 73749 101085 73777 101113
rect 73811 101085 73839 101113
rect 73625 101023 73653 101051
rect 73687 101023 73715 101051
rect 73749 101023 73777 101051
rect 73811 101023 73839 101051
rect 73625 100961 73653 100989
rect 73687 100961 73715 100989
rect 73749 100961 73777 100989
rect 73811 100961 73839 100989
rect 66485 95147 66513 95175
rect 66547 95147 66575 95175
rect 66609 95147 66637 95175
rect 66671 95147 66699 95175
rect 66485 95085 66513 95113
rect 66547 95085 66575 95113
rect 66609 95085 66637 95113
rect 66671 95085 66699 95113
rect 66485 95023 66513 95051
rect 66547 95023 66575 95051
rect 66609 95023 66637 95051
rect 66671 95023 66699 95051
rect 66485 94961 66513 94989
rect 66547 94961 66575 94989
rect 66609 94961 66637 94989
rect 66671 94961 66699 94989
rect 64625 92147 64653 92175
rect 64687 92147 64715 92175
rect 64749 92147 64777 92175
rect 64811 92147 64839 92175
rect 64625 92085 64653 92113
rect 64687 92085 64715 92113
rect 64749 92085 64777 92113
rect 64811 92085 64839 92113
rect 64625 92023 64653 92051
rect 64687 92023 64715 92051
rect 64749 92023 64777 92051
rect 64811 92023 64839 92051
rect 64625 91961 64653 91989
rect 64687 91961 64715 91989
rect 64749 91961 64777 91989
rect 64811 91961 64839 91989
rect 57485 86147 57513 86175
rect 57547 86147 57575 86175
rect 57609 86147 57637 86175
rect 57671 86147 57699 86175
rect 57485 86085 57513 86113
rect 57547 86085 57575 86113
rect 57609 86085 57637 86113
rect 57671 86085 57699 86113
rect 57485 86023 57513 86051
rect 57547 86023 57575 86051
rect 57609 86023 57637 86051
rect 57671 86023 57699 86051
rect 57485 85961 57513 85989
rect 57547 85961 57575 85989
rect 57609 85961 57637 85989
rect 57671 85961 57699 85989
rect 55625 83147 55653 83175
rect 55687 83147 55715 83175
rect 55749 83147 55777 83175
rect 55811 83147 55839 83175
rect 55625 83085 55653 83113
rect 55687 83085 55715 83113
rect 55749 83085 55777 83113
rect 55811 83085 55839 83113
rect 55625 83023 55653 83051
rect 55687 83023 55715 83051
rect 55749 83023 55777 83051
rect 55811 83023 55839 83051
rect 55625 82961 55653 82989
rect 55687 82961 55715 82989
rect 55749 82961 55777 82989
rect 55811 82961 55839 82989
rect 48485 77147 48513 77175
rect 48547 77147 48575 77175
rect 48609 77147 48637 77175
rect 48671 77147 48699 77175
rect 48485 77085 48513 77113
rect 48547 77085 48575 77113
rect 48609 77085 48637 77113
rect 48671 77085 48699 77113
rect 48485 77023 48513 77051
rect 48547 77023 48575 77051
rect 48609 77023 48637 77051
rect 48671 77023 48699 77051
rect 48485 76961 48513 76989
rect 48547 76961 48575 76989
rect 48609 76961 48637 76989
rect 48671 76961 48699 76989
rect 54509 77147 54537 77175
rect 54571 77147 54599 77175
rect 54509 77085 54537 77113
rect 54571 77085 54599 77113
rect 54509 77023 54537 77051
rect 54571 77023 54599 77051
rect 54509 76961 54537 76989
rect 54571 76961 54599 76989
rect 52259 74147 52287 74175
rect 52321 74147 52349 74175
rect 52259 74085 52287 74113
rect 52321 74085 52349 74113
rect 52259 74023 52287 74051
rect 52321 74023 52349 74051
rect 52259 73961 52287 73989
rect 52321 73961 52349 73989
rect 56759 83147 56787 83175
rect 56821 83147 56849 83175
rect 56759 83085 56787 83113
rect 56821 83085 56849 83113
rect 56759 83023 56787 83051
rect 56821 83023 56849 83051
rect 56759 82961 56787 82989
rect 56821 82961 56849 82989
rect 59009 86147 59037 86175
rect 59071 86147 59099 86175
rect 59009 86085 59037 86113
rect 59071 86085 59099 86113
rect 59009 86023 59037 86051
rect 59071 86023 59099 86051
rect 59009 85961 59037 85989
rect 59071 85961 59099 85989
rect 63509 86147 63537 86175
rect 63571 86147 63599 86175
rect 63509 86085 63537 86113
rect 63571 86085 63599 86113
rect 63509 86023 63537 86051
rect 63571 86023 63599 86051
rect 63509 85961 63537 85989
rect 63571 85961 63599 85989
rect 61259 83147 61287 83175
rect 61321 83147 61349 83175
rect 61259 83085 61287 83113
rect 61321 83085 61349 83113
rect 61259 83023 61287 83051
rect 61321 83023 61349 83051
rect 61259 82961 61287 82989
rect 61321 82961 61349 82989
rect 65759 92147 65787 92175
rect 65821 92147 65849 92175
rect 65759 92085 65787 92113
rect 65821 92085 65849 92113
rect 65759 92023 65787 92051
rect 65821 92023 65849 92051
rect 65759 91961 65787 91989
rect 65821 91961 65849 91989
rect 68009 95147 68037 95175
rect 68071 95147 68099 95175
rect 68009 95085 68037 95113
rect 68071 95085 68099 95113
rect 68009 95023 68037 95051
rect 68071 95023 68099 95051
rect 68009 94961 68037 94989
rect 68071 94961 68099 94989
rect 72509 95147 72537 95175
rect 72571 95147 72599 95175
rect 72509 95085 72537 95113
rect 72571 95085 72599 95113
rect 72509 95023 72537 95051
rect 72571 95023 72599 95051
rect 72509 94961 72537 94989
rect 72571 94961 72599 94989
rect 70259 92147 70287 92175
rect 70321 92147 70349 92175
rect 70259 92085 70287 92113
rect 70321 92085 70349 92113
rect 70259 92023 70287 92051
rect 70321 92023 70349 92051
rect 70259 91961 70287 91989
rect 70321 91961 70349 91989
rect 74759 101147 74787 101175
rect 74821 101147 74849 101175
rect 74759 101085 74787 101113
rect 74821 101085 74849 101113
rect 74759 101023 74787 101051
rect 74821 101023 74849 101051
rect 74759 100961 74787 100989
rect 74821 100961 74849 100989
rect 77009 104147 77037 104175
rect 77071 104147 77099 104175
rect 77009 104085 77037 104113
rect 77071 104085 77099 104113
rect 77009 104023 77037 104051
rect 77071 104023 77099 104051
rect 77009 103961 77037 103989
rect 77071 103961 77099 103989
rect 81509 104147 81537 104175
rect 81571 104147 81599 104175
rect 81509 104085 81537 104113
rect 81571 104085 81599 104113
rect 81509 104023 81537 104051
rect 81571 104023 81599 104051
rect 81509 103961 81537 103989
rect 81571 103961 81599 103989
rect 79259 101147 79287 101175
rect 79321 101147 79349 101175
rect 79259 101085 79287 101113
rect 79321 101085 79349 101113
rect 79259 101023 79287 101051
rect 79321 101023 79349 101051
rect 79259 100961 79287 100989
rect 79321 100961 79349 100989
rect 84485 122147 84513 122175
rect 84547 122147 84575 122175
rect 84609 122147 84637 122175
rect 84671 122147 84699 122175
rect 84485 122085 84513 122113
rect 84547 122085 84575 122113
rect 84609 122085 84637 122113
rect 84671 122085 84699 122113
rect 84485 122023 84513 122051
rect 84547 122023 84575 122051
rect 84609 122023 84637 122051
rect 84671 122023 84699 122051
rect 84485 121961 84513 121989
rect 84547 121961 84575 121989
rect 84609 121961 84637 121989
rect 84671 121961 84699 121989
rect 84485 113147 84513 113175
rect 84547 113147 84575 113175
rect 84609 113147 84637 113175
rect 84671 113147 84699 113175
rect 84485 113085 84513 113113
rect 84547 113085 84575 113113
rect 84609 113085 84637 113113
rect 84671 113085 84699 113113
rect 84485 113023 84513 113051
rect 84547 113023 84575 113051
rect 84609 113023 84637 113051
rect 84671 113023 84699 113051
rect 84485 112961 84513 112989
rect 84547 112961 84575 112989
rect 84609 112961 84637 112989
rect 84671 112961 84699 112989
rect 91625 119147 91653 119175
rect 91687 119147 91715 119175
rect 91749 119147 91777 119175
rect 91811 119147 91839 119175
rect 91625 119085 91653 119113
rect 91687 119085 91715 119113
rect 91749 119085 91777 119113
rect 91811 119085 91839 119113
rect 91625 119023 91653 119051
rect 91687 119023 91715 119051
rect 91749 119023 91777 119051
rect 91811 119023 91839 119051
rect 91625 118961 91653 118989
rect 91687 118961 91715 118989
rect 91749 118961 91777 118989
rect 91811 118961 91839 118989
rect 91625 110147 91653 110175
rect 91687 110147 91715 110175
rect 91749 110147 91777 110175
rect 91811 110147 91839 110175
rect 91625 110085 91653 110113
rect 91687 110085 91715 110113
rect 91749 110085 91777 110113
rect 91811 110085 91839 110113
rect 91625 110023 91653 110051
rect 91687 110023 91715 110051
rect 91749 110023 91777 110051
rect 91811 110023 91839 110051
rect 91625 109961 91653 109989
rect 91687 109961 91715 109989
rect 91749 109961 91777 109989
rect 91811 109961 91839 109989
rect 84485 104147 84513 104175
rect 84547 104147 84575 104175
rect 84609 104147 84637 104175
rect 84671 104147 84699 104175
rect 84485 104085 84513 104113
rect 84547 104085 84575 104113
rect 84609 104085 84637 104113
rect 84671 104085 84699 104113
rect 84485 104023 84513 104051
rect 84547 104023 84575 104051
rect 84609 104023 84637 104051
rect 84671 104023 84699 104051
rect 84485 103961 84513 103989
rect 84547 103961 84575 103989
rect 84609 103961 84637 103989
rect 84671 103961 84699 103989
rect 82625 101147 82653 101175
rect 82687 101147 82715 101175
rect 82749 101147 82777 101175
rect 82811 101147 82839 101175
rect 82625 101085 82653 101113
rect 82687 101085 82715 101113
rect 82749 101085 82777 101113
rect 82811 101085 82839 101113
rect 82625 101023 82653 101051
rect 82687 101023 82715 101051
rect 82749 101023 82777 101051
rect 82811 101023 82839 101051
rect 82625 100961 82653 100989
rect 82687 100961 82715 100989
rect 82749 100961 82777 100989
rect 82811 100961 82839 100989
rect 75485 95147 75513 95175
rect 75547 95147 75575 95175
rect 75609 95147 75637 95175
rect 75671 95147 75699 95175
rect 75485 95085 75513 95113
rect 75547 95085 75575 95113
rect 75609 95085 75637 95113
rect 75671 95085 75699 95113
rect 75485 95023 75513 95051
rect 75547 95023 75575 95051
rect 75609 95023 75637 95051
rect 75671 95023 75699 95051
rect 75485 94961 75513 94989
rect 75547 94961 75575 94989
rect 75609 94961 75637 94989
rect 75671 94961 75699 94989
rect 73625 92147 73653 92175
rect 73687 92147 73715 92175
rect 73749 92147 73777 92175
rect 73811 92147 73839 92175
rect 73625 92085 73653 92113
rect 73687 92085 73715 92113
rect 73749 92085 73777 92113
rect 73811 92085 73839 92113
rect 73625 92023 73653 92051
rect 73687 92023 73715 92051
rect 73749 92023 73777 92051
rect 73811 92023 73839 92051
rect 73625 91961 73653 91989
rect 73687 91961 73715 91989
rect 73749 91961 73777 91989
rect 73811 91961 73839 91989
rect 66485 86147 66513 86175
rect 66547 86147 66575 86175
rect 66609 86147 66637 86175
rect 66671 86147 66699 86175
rect 66485 86085 66513 86113
rect 66547 86085 66575 86113
rect 66609 86085 66637 86113
rect 66671 86085 66699 86113
rect 66485 86023 66513 86051
rect 66547 86023 66575 86051
rect 66609 86023 66637 86051
rect 66671 86023 66699 86051
rect 66485 85961 66513 85989
rect 66547 85961 66575 85989
rect 66609 85961 66637 85989
rect 66671 85961 66699 85989
rect 64625 83147 64653 83175
rect 64687 83147 64715 83175
rect 64749 83147 64777 83175
rect 64811 83147 64839 83175
rect 64625 83085 64653 83113
rect 64687 83085 64715 83113
rect 64749 83085 64777 83113
rect 64811 83085 64839 83113
rect 64625 83023 64653 83051
rect 64687 83023 64715 83051
rect 64749 83023 64777 83051
rect 64811 83023 64839 83051
rect 64625 82961 64653 82989
rect 64687 82961 64715 82989
rect 64749 82961 64777 82989
rect 64811 82961 64839 82989
rect 57485 77147 57513 77175
rect 57547 77147 57575 77175
rect 57609 77147 57637 77175
rect 57671 77147 57699 77175
rect 57485 77085 57513 77113
rect 57547 77085 57575 77113
rect 57609 77085 57637 77113
rect 57671 77085 57699 77113
rect 57485 77023 57513 77051
rect 57547 77023 57575 77051
rect 57609 77023 57637 77051
rect 57671 77023 57699 77051
rect 57485 76961 57513 76989
rect 57547 76961 57575 76989
rect 57609 76961 57637 76989
rect 57671 76961 57699 76989
rect 55625 74147 55653 74175
rect 55687 74147 55715 74175
rect 55749 74147 55777 74175
rect 55811 74147 55839 74175
rect 55625 74085 55653 74113
rect 55687 74085 55715 74113
rect 55749 74085 55777 74113
rect 55811 74085 55839 74113
rect 55625 74023 55653 74051
rect 55687 74023 55715 74051
rect 55749 74023 55777 74051
rect 55811 74023 55839 74051
rect 55625 73961 55653 73989
rect 55687 73961 55715 73989
rect 55749 73961 55777 73989
rect 55811 73961 55839 73989
rect 48485 68147 48513 68175
rect 48547 68147 48575 68175
rect 48609 68147 48637 68175
rect 48671 68147 48699 68175
rect 48485 68085 48513 68113
rect 48547 68085 48575 68113
rect 48609 68085 48637 68113
rect 48671 68085 48699 68113
rect 48485 68023 48513 68051
rect 48547 68023 48575 68051
rect 48609 68023 48637 68051
rect 48671 68023 48699 68051
rect 48485 67961 48513 67989
rect 48547 67961 48575 67989
rect 48609 67961 48637 67989
rect 48671 67961 48699 67989
rect 54509 68147 54537 68175
rect 54571 68147 54599 68175
rect 54509 68085 54537 68113
rect 54571 68085 54599 68113
rect 54509 68023 54537 68051
rect 54571 68023 54599 68051
rect 54509 67961 54537 67989
rect 54571 67961 54599 67989
rect 52259 65147 52287 65175
rect 52321 65147 52349 65175
rect 52259 65085 52287 65113
rect 52321 65085 52349 65113
rect 52259 65023 52287 65051
rect 52321 65023 52349 65051
rect 52259 64961 52287 64989
rect 52321 64961 52349 64989
rect 56759 74147 56787 74175
rect 56821 74147 56849 74175
rect 56759 74085 56787 74113
rect 56821 74085 56849 74113
rect 56759 74023 56787 74051
rect 56821 74023 56849 74051
rect 56759 73961 56787 73989
rect 56821 73961 56849 73989
rect 59009 77147 59037 77175
rect 59071 77147 59099 77175
rect 59009 77085 59037 77113
rect 59071 77085 59099 77113
rect 59009 77023 59037 77051
rect 59071 77023 59099 77051
rect 59009 76961 59037 76989
rect 59071 76961 59099 76989
rect 63509 77147 63537 77175
rect 63571 77147 63599 77175
rect 63509 77085 63537 77113
rect 63571 77085 63599 77113
rect 63509 77023 63537 77051
rect 63571 77023 63599 77051
rect 63509 76961 63537 76989
rect 63571 76961 63599 76989
rect 61259 74147 61287 74175
rect 61321 74147 61349 74175
rect 61259 74085 61287 74113
rect 61321 74085 61349 74113
rect 61259 74023 61287 74051
rect 61321 74023 61349 74051
rect 61259 73961 61287 73989
rect 61321 73961 61349 73989
rect 65759 83147 65787 83175
rect 65821 83147 65849 83175
rect 65759 83085 65787 83113
rect 65821 83085 65849 83113
rect 65759 83023 65787 83051
rect 65821 83023 65849 83051
rect 65759 82961 65787 82989
rect 65821 82961 65849 82989
rect 68009 86147 68037 86175
rect 68071 86147 68099 86175
rect 68009 86085 68037 86113
rect 68071 86085 68099 86113
rect 68009 86023 68037 86051
rect 68071 86023 68099 86051
rect 68009 85961 68037 85989
rect 68071 85961 68099 85989
rect 72509 86147 72537 86175
rect 72571 86147 72599 86175
rect 72509 86085 72537 86113
rect 72571 86085 72599 86113
rect 72509 86023 72537 86051
rect 72571 86023 72599 86051
rect 72509 85961 72537 85989
rect 72571 85961 72599 85989
rect 70259 83147 70287 83175
rect 70321 83147 70349 83175
rect 70259 83085 70287 83113
rect 70321 83085 70349 83113
rect 70259 83023 70287 83051
rect 70321 83023 70349 83051
rect 70259 82961 70287 82989
rect 70321 82961 70349 82989
rect 74759 92147 74787 92175
rect 74821 92147 74849 92175
rect 74759 92085 74787 92113
rect 74821 92085 74849 92113
rect 74759 92023 74787 92051
rect 74821 92023 74849 92051
rect 74759 91961 74787 91989
rect 74821 91961 74849 91989
rect 77009 95147 77037 95175
rect 77071 95147 77099 95175
rect 77009 95085 77037 95113
rect 77071 95085 77099 95113
rect 77009 95023 77037 95051
rect 77071 95023 77099 95051
rect 77009 94961 77037 94989
rect 77071 94961 77099 94989
rect 81509 95147 81537 95175
rect 81571 95147 81599 95175
rect 81509 95085 81537 95113
rect 81571 95085 81599 95113
rect 81509 95023 81537 95051
rect 81571 95023 81599 95051
rect 81509 94961 81537 94989
rect 81571 94961 81599 94989
rect 79259 92147 79287 92175
rect 79321 92147 79349 92175
rect 79259 92085 79287 92113
rect 79321 92085 79349 92113
rect 79259 92023 79287 92051
rect 79321 92023 79349 92051
rect 79259 91961 79287 91989
rect 79321 91961 79349 91989
rect 83759 101147 83787 101175
rect 83821 101147 83849 101175
rect 83759 101085 83787 101113
rect 83821 101085 83849 101113
rect 83759 101023 83787 101051
rect 83821 101023 83849 101051
rect 83759 100961 83787 100989
rect 83821 100961 83849 100989
rect 86009 104147 86037 104175
rect 86071 104147 86099 104175
rect 86009 104085 86037 104113
rect 86071 104085 86099 104113
rect 86009 104023 86037 104051
rect 86071 104023 86099 104051
rect 86009 103961 86037 103989
rect 86071 103961 86099 103989
rect 90509 104147 90537 104175
rect 90571 104147 90599 104175
rect 90509 104085 90537 104113
rect 90571 104085 90599 104113
rect 90509 104023 90537 104051
rect 90571 104023 90599 104051
rect 90509 103961 90537 103989
rect 90571 103961 90599 103989
rect 88259 101147 88287 101175
rect 88321 101147 88349 101175
rect 88259 101085 88287 101113
rect 88321 101085 88349 101113
rect 88259 101023 88287 101051
rect 88321 101023 88349 101051
rect 88259 100961 88287 100989
rect 88321 100961 88349 100989
rect 93485 122147 93513 122175
rect 93547 122147 93575 122175
rect 93609 122147 93637 122175
rect 93671 122147 93699 122175
rect 93485 122085 93513 122113
rect 93547 122085 93575 122113
rect 93609 122085 93637 122113
rect 93671 122085 93699 122113
rect 93485 122023 93513 122051
rect 93547 122023 93575 122051
rect 93609 122023 93637 122051
rect 93671 122023 93699 122051
rect 93485 121961 93513 121989
rect 93547 121961 93575 121989
rect 93609 121961 93637 121989
rect 93671 121961 93699 121989
rect 93485 113147 93513 113175
rect 93547 113147 93575 113175
rect 93609 113147 93637 113175
rect 93671 113147 93699 113175
rect 93485 113085 93513 113113
rect 93547 113085 93575 113113
rect 93609 113085 93637 113113
rect 93671 113085 93699 113113
rect 93485 113023 93513 113051
rect 93547 113023 93575 113051
rect 93609 113023 93637 113051
rect 93671 113023 93699 113051
rect 93485 112961 93513 112989
rect 93547 112961 93575 112989
rect 93609 112961 93637 112989
rect 93671 112961 93699 112989
rect 100625 119147 100653 119175
rect 100687 119147 100715 119175
rect 100749 119147 100777 119175
rect 100811 119147 100839 119175
rect 100625 119085 100653 119113
rect 100687 119085 100715 119113
rect 100749 119085 100777 119113
rect 100811 119085 100839 119113
rect 100625 119023 100653 119051
rect 100687 119023 100715 119051
rect 100749 119023 100777 119051
rect 100811 119023 100839 119051
rect 100625 118961 100653 118989
rect 100687 118961 100715 118989
rect 100749 118961 100777 118989
rect 100811 118961 100839 118989
rect 100625 110147 100653 110175
rect 100687 110147 100715 110175
rect 100749 110147 100777 110175
rect 100811 110147 100839 110175
rect 100625 110085 100653 110113
rect 100687 110085 100715 110113
rect 100749 110085 100777 110113
rect 100811 110085 100839 110113
rect 100625 110023 100653 110051
rect 100687 110023 100715 110051
rect 100749 110023 100777 110051
rect 100811 110023 100839 110051
rect 100625 109961 100653 109989
rect 100687 109961 100715 109989
rect 100749 109961 100777 109989
rect 100811 109961 100839 109989
rect 93485 104147 93513 104175
rect 93547 104147 93575 104175
rect 93609 104147 93637 104175
rect 93671 104147 93699 104175
rect 93485 104085 93513 104113
rect 93547 104085 93575 104113
rect 93609 104085 93637 104113
rect 93671 104085 93699 104113
rect 93485 104023 93513 104051
rect 93547 104023 93575 104051
rect 93609 104023 93637 104051
rect 93671 104023 93699 104051
rect 93485 103961 93513 103989
rect 93547 103961 93575 103989
rect 93609 103961 93637 103989
rect 93671 103961 93699 103989
rect 91625 101147 91653 101175
rect 91687 101147 91715 101175
rect 91749 101147 91777 101175
rect 91811 101147 91839 101175
rect 91625 101085 91653 101113
rect 91687 101085 91715 101113
rect 91749 101085 91777 101113
rect 91811 101085 91839 101113
rect 91625 101023 91653 101051
rect 91687 101023 91715 101051
rect 91749 101023 91777 101051
rect 91811 101023 91839 101051
rect 91625 100961 91653 100989
rect 91687 100961 91715 100989
rect 91749 100961 91777 100989
rect 91811 100961 91839 100989
rect 84485 95147 84513 95175
rect 84547 95147 84575 95175
rect 84609 95147 84637 95175
rect 84671 95147 84699 95175
rect 84485 95085 84513 95113
rect 84547 95085 84575 95113
rect 84609 95085 84637 95113
rect 84671 95085 84699 95113
rect 84485 95023 84513 95051
rect 84547 95023 84575 95051
rect 84609 95023 84637 95051
rect 84671 95023 84699 95051
rect 84485 94961 84513 94989
rect 84547 94961 84575 94989
rect 84609 94961 84637 94989
rect 84671 94961 84699 94989
rect 82625 92147 82653 92175
rect 82687 92147 82715 92175
rect 82749 92147 82777 92175
rect 82811 92147 82839 92175
rect 82625 92085 82653 92113
rect 82687 92085 82715 92113
rect 82749 92085 82777 92113
rect 82811 92085 82839 92113
rect 82625 92023 82653 92051
rect 82687 92023 82715 92051
rect 82749 92023 82777 92051
rect 82811 92023 82839 92051
rect 82625 91961 82653 91989
rect 82687 91961 82715 91989
rect 82749 91961 82777 91989
rect 82811 91961 82839 91989
rect 75485 86147 75513 86175
rect 75547 86147 75575 86175
rect 75609 86147 75637 86175
rect 75671 86147 75699 86175
rect 75485 86085 75513 86113
rect 75547 86085 75575 86113
rect 75609 86085 75637 86113
rect 75671 86085 75699 86113
rect 75485 86023 75513 86051
rect 75547 86023 75575 86051
rect 75609 86023 75637 86051
rect 75671 86023 75699 86051
rect 75485 85961 75513 85989
rect 75547 85961 75575 85989
rect 75609 85961 75637 85989
rect 75671 85961 75699 85989
rect 73625 83147 73653 83175
rect 73687 83147 73715 83175
rect 73749 83147 73777 83175
rect 73811 83147 73839 83175
rect 73625 83085 73653 83113
rect 73687 83085 73715 83113
rect 73749 83085 73777 83113
rect 73811 83085 73839 83113
rect 73625 83023 73653 83051
rect 73687 83023 73715 83051
rect 73749 83023 73777 83051
rect 73811 83023 73839 83051
rect 73625 82961 73653 82989
rect 73687 82961 73715 82989
rect 73749 82961 73777 82989
rect 73811 82961 73839 82989
rect 66485 77147 66513 77175
rect 66547 77147 66575 77175
rect 66609 77147 66637 77175
rect 66671 77147 66699 77175
rect 66485 77085 66513 77113
rect 66547 77085 66575 77113
rect 66609 77085 66637 77113
rect 66671 77085 66699 77113
rect 66485 77023 66513 77051
rect 66547 77023 66575 77051
rect 66609 77023 66637 77051
rect 66671 77023 66699 77051
rect 66485 76961 66513 76989
rect 66547 76961 66575 76989
rect 66609 76961 66637 76989
rect 66671 76961 66699 76989
rect 64625 74147 64653 74175
rect 64687 74147 64715 74175
rect 64749 74147 64777 74175
rect 64811 74147 64839 74175
rect 64625 74085 64653 74113
rect 64687 74085 64715 74113
rect 64749 74085 64777 74113
rect 64811 74085 64839 74113
rect 64625 74023 64653 74051
rect 64687 74023 64715 74051
rect 64749 74023 64777 74051
rect 64811 74023 64839 74051
rect 64625 73961 64653 73989
rect 64687 73961 64715 73989
rect 64749 73961 64777 73989
rect 64811 73961 64839 73989
rect 57485 68147 57513 68175
rect 57547 68147 57575 68175
rect 57609 68147 57637 68175
rect 57671 68147 57699 68175
rect 57485 68085 57513 68113
rect 57547 68085 57575 68113
rect 57609 68085 57637 68113
rect 57671 68085 57699 68113
rect 57485 68023 57513 68051
rect 57547 68023 57575 68051
rect 57609 68023 57637 68051
rect 57671 68023 57699 68051
rect 57485 67961 57513 67989
rect 57547 67961 57575 67989
rect 57609 67961 57637 67989
rect 57671 67961 57699 67989
rect 55625 65147 55653 65175
rect 55687 65147 55715 65175
rect 55749 65147 55777 65175
rect 55811 65147 55839 65175
rect 55625 65085 55653 65113
rect 55687 65085 55715 65113
rect 55749 65085 55777 65113
rect 55811 65085 55839 65113
rect 55625 65023 55653 65051
rect 55687 65023 55715 65051
rect 55749 65023 55777 65051
rect 55811 65023 55839 65051
rect 55625 64961 55653 64989
rect 55687 64961 55715 64989
rect 55749 64961 55777 64989
rect 55811 64961 55839 64989
rect 48485 59147 48513 59175
rect 48547 59147 48575 59175
rect 48609 59147 48637 59175
rect 48671 59147 48699 59175
rect 48485 59085 48513 59113
rect 48547 59085 48575 59113
rect 48609 59085 48637 59113
rect 48671 59085 48699 59113
rect 48485 59023 48513 59051
rect 48547 59023 48575 59051
rect 48609 59023 48637 59051
rect 48671 59023 48699 59051
rect 48485 58961 48513 58989
rect 48547 58961 48575 58989
rect 48609 58961 48637 58989
rect 48671 58961 48699 58989
rect 54509 59147 54537 59175
rect 54571 59147 54599 59175
rect 54509 59085 54537 59113
rect 54571 59085 54599 59113
rect 54509 59023 54537 59051
rect 54571 59023 54599 59051
rect 54509 58961 54537 58989
rect 54571 58961 54599 58989
rect 52259 56147 52287 56175
rect 52321 56147 52349 56175
rect 52259 56085 52287 56113
rect 52321 56085 52349 56113
rect 52259 56023 52287 56051
rect 52321 56023 52349 56051
rect 52259 55961 52287 55989
rect 52321 55961 52349 55989
rect 56759 65147 56787 65175
rect 56821 65147 56849 65175
rect 56759 65085 56787 65113
rect 56821 65085 56849 65113
rect 56759 65023 56787 65051
rect 56821 65023 56849 65051
rect 56759 64961 56787 64989
rect 56821 64961 56849 64989
rect 59009 68147 59037 68175
rect 59071 68147 59099 68175
rect 59009 68085 59037 68113
rect 59071 68085 59099 68113
rect 59009 68023 59037 68051
rect 59071 68023 59099 68051
rect 59009 67961 59037 67989
rect 59071 67961 59099 67989
rect 63509 68147 63537 68175
rect 63571 68147 63599 68175
rect 63509 68085 63537 68113
rect 63571 68085 63599 68113
rect 63509 68023 63537 68051
rect 63571 68023 63599 68051
rect 63509 67961 63537 67989
rect 63571 67961 63599 67989
rect 61259 65147 61287 65175
rect 61321 65147 61349 65175
rect 61259 65085 61287 65113
rect 61321 65085 61349 65113
rect 61259 65023 61287 65051
rect 61321 65023 61349 65051
rect 61259 64961 61287 64989
rect 61321 64961 61349 64989
rect 65759 74147 65787 74175
rect 65821 74147 65849 74175
rect 65759 74085 65787 74113
rect 65821 74085 65849 74113
rect 65759 74023 65787 74051
rect 65821 74023 65849 74051
rect 65759 73961 65787 73989
rect 65821 73961 65849 73989
rect 68009 77147 68037 77175
rect 68071 77147 68099 77175
rect 68009 77085 68037 77113
rect 68071 77085 68099 77113
rect 68009 77023 68037 77051
rect 68071 77023 68099 77051
rect 68009 76961 68037 76989
rect 68071 76961 68099 76989
rect 72509 77147 72537 77175
rect 72571 77147 72599 77175
rect 72509 77085 72537 77113
rect 72571 77085 72599 77113
rect 72509 77023 72537 77051
rect 72571 77023 72599 77051
rect 72509 76961 72537 76989
rect 72571 76961 72599 76989
rect 70259 74147 70287 74175
rect 70321 74147 70349 74175
rect 70259 74085 70287 74113
rect 70321 74085 70349 74113
rect 70259 74023 70287 74051
rect 70321 74023 70349 74051
rect 70259 73961 70287 73989
rect 70321 73961 70349 73989
rect 74759 83147 74787 83175
rect 74821 83147 74849 83175
rect 74759 83085 74787 83113
rect 74821 83085 74849 83113
rect 74759 83023 74787 83051
rect 74821 83023 74849 83051
rect 74759 82961 74787 82989
rect 74821 82961 74849 82989
rect 77009 86147 77037 86175
rect 77071 86147 77099 86175
rect 77009 86085 77037 86113
rect 77071 86085 77099 86113
rect 77009 86023 77037 86051
rect 77071 86023 77099 86051
rect 77009 85961 77037 85989
rect 77071 85961 77099 85989
rect 81509 86147 81537 86175
rect 81571 86147 81599 86175
rect 81509 86085 81537 86113
rect 81571 86085 81599 86113
rect 81509 86023 81537 86051
rect 81571 86023 81599 86051
rect 81509 85961 81537 85989
rect 81571 85961 81599 85989
rect 79259 83147 79287 83175
rect 79321 83147 79349 83175
rect 79259 83085 79287 83113
rect 79321 83085 79349 83113
rect 79259 83023 79287 83051
rect 79321 83023 79349 83051
rect 79259 82961 79287 82989
rect 79321 82961 79349 82989
rect 83759 92147 83787 92175
rect 83821 92147 83849 92175
rect 83759 92085 83787 92113
rect 83821 92085 83849 92113
rect 83759 92023 83787 92051
rect 83821 92023 83849 92051
rect 83759 91961 83787 91989
rect 83821 91961 83849 91989
rect 86009 95147 86037 95175
rect 86071 95147 86099 95175
rect 86009 95085 86037 95113
rect 86071 95085 86099 95113
rect 86009 95023 86037 95051
rect 86071 95023 86099 95051
rect 86009 94961 86037 94989
rect 86071 94961 86099 94989
rect 90509 95147 90537 95175
rect 90571 95147 90599 95175
rect 90509 95085 90537 95113
rect 90571 95085 90599 95113
rect 90509 95023 90537 95051
rect 90571 95023 90599 95051
rect 90509 94961 90537 94989
rect 90571 94961 90599 94989
rect 88259 92147 88287 92175
rect 88321 92147 88349 92175
rect 88259 92085 88287 92113
rect 88321 92085 88349 92113
rect 88259 92023 88287 92051
rect 88321 92023 88349 92051
rect 88259 91961 88287 91989
rect 88321 91961 88349 91989
rect 92759 101147 92787 101175
rect 92821 101147 92849 101175
rect 92759 101085 92787 101113
rect 92821 101085 92849 101113
rect 92759 101023 92787 101051
rect 92821 101023 92849 101051
rect 92759 100961 92787 100989
rect 92821 100961 92849 100989
rect 95009 104147 95037 104175
rect 95071 104147 95099 104175
rect 95009 104085 95037 104113
rect 95071 104085 95099 104113
rect 95009 104023 95037 104051
rect 95071 104023 95099 104051
rect 95009 103961 95037 103989
rect 95071 103961 95099 103989
rect 99509 104147 99537 104175
rect 99571 104147 99599 104175
rect 99509 104085 99537 104113
rect 99571 104085 99599 104113
rect 99509 104023 99537 104051
rect 99571 104023 99599 104051
rect 99509 103961 99537 103989
rect 99571 103961 99599 103989
rect 97259 101147 97287 101175
rect 97321 101147 97349 101175
rect 97259 101085 97287 101113
rect 97321 101085 97349 101113
rect 97259 101023 97287 101051
rect 97321 101023 97349 101051
rect 97259 100961 97287 100989
rect 97321 100961 97349 100989
rect 102485 122147 102513 122175
rect 102547 122147 102575 122175
rect 102609 122147 102637 122175
rect 102671 122147 102699 122175
rect 102485 122085 102513 122113
rect 102547 122085 102575 122113
rect 102609 122085 102637 122113
rect 102671 122085 102699 122113
rect 102485 122023 102513 122051
rect 102547 122023 102575 122051
rect 102609 122023 102637 122051
rect 102671 122023 102699 122051
rect 102485 121961 102513 121989
rect 102547 121961 102575 121989
rect 102609 121961 102637 121989
rect 102671 121961 102699 121989
rect 102485 113147 102513 113175
rect 102547 113147 102575 113175
rect 102609 113147 102637 113175
rect 102671 113147 102699 113175
rect 102485 113085 102513 113113
rect 102547 113085 102575 113113
rect 102609 113085 102637 113113
rect 102671 113085 102699 113113
rect 102485 113023 102513 113051
rect 102547 113023 102575 113051
rect 102609 113023 102637 113051
rect 102671 113023 102699 113051
rect 102485 112961 102513 112989
rect 102547 112961 102575 112989
rect 102609 112961 102637 112989
rect 102671 112961 102699 112989
rect 109625 119147 109653 119175
rect 109687 119147 109715 119175
rect 109749 119147 109777 119175
rect 109811 119147 109839 119175
rect 109625 119085 109653 119113
rect 109687 119085 109715 119113
rect 109749 119085 109777 119113
rect 109811 119085 109839 119113
rect 109625 119023 109653 119051
rect 109687 119023 109715 119051
rect 109749 119023 109777 119051
rect 109811 119023 109839 119051
rect 109625 118961 109653 118989
rect 109687 118961 109715 118989
rect 109749 118961 109777 118989
rect 109811 118961 109839 118989
rect 109625 110147 109653 110175
rect 109687 110147 109715 110175
rect 109749 110147 109777 110175
rect 109811 110147 109839 110175
rect 109625 110085 109653 110113
rect 109687 110085 109715 110113
rect 109749 110085 109777 110113
rect 109811 110085 109839 110113
rect 109625 110023 109653 110051
rect 109687 110023 109715 110051
rect 109749 110023 109777 110051
rect 109811 110023 109839 110051
rect 109625 109961 109653 109989
rect 109687 109961 109715 109989
rect 109749 109961 109777 109989
rect 109811 109961 109839 109989
rect 102485 104147 102513 104175
rect 102547 104147 102575 104175
rect 102609 104147 102637 104175
rect 102671 104147 102699 104175
rect 102485 104085 102513 104113
rect 102547 104085 102575 104113
rect 102609 104085 102637 104113
rect 102671 104085 102699 104113
rect 102485 104023 102513 104051
rect 102547 104023 102575 104051
rect 102609 104023 102637 104051
rect 102671 104023 102699 104051
rect 102485 103961 102513 103989
rect 102547 103961 102575 103989
rect 102609 103961 102637 103989
rect 102671 103961 102699 103989
rect 100625 101147 100653 101175
rect 100687 101147 100715 101175
rect 100749 101147 100777 101175
rect 100811 101147 100839 101175
rect 100625 101085 100653 101113
rect 100687 101085 100715 101113
rect 100749 101085 100777 101113
rect 100811 101085 100839 101113
rect 100625 101023 100653 101051
rect 100687 101023 100715 101051
rect 100749 101023 100777 101051
rect 100811 101023 100839 101051
rect 100625 100961 100653 100989
rect 100687 100961 100715 100989
rect 100749 100961 100777 100989
rect 100811 100961 100839 100989
rect 101759 101147 101787 101175
rect 101821 101147 101849 101175
rect 101759 101085 101787 101113
rect 101821 101085 101849 101113
rect 101759 101023 101787 101051
rect 101821 101023 101849 101051
rect 101759 100961 101787 100989
rect 101821 100961 101849 100989
rect 104009 104147 104037 104175
rect 104071 104147 104099 104175
rect 104009 104085 104037 104113
rect 104071 104085 104099 104113
rect 104009 104023 104037 104051
rect 104071 104023 104099 104051
rect 104009 103961 104037 103989
rect 104071 103961 104099 103989
rect 108509 104147 108537 104175
rect 108571 104147 108599 104175
rect 108509 104085 108537 104113
rect 108571 104085 108599 104113
rect 108509 104023 108537 104051
rect 108571 104023 108599 104051
rect 108509 103961 108537 103989
rect 108571 103961 108599 103989
rect 106259 101147 106287 101175
rect 106321 101147 106349 101175
rect 106259 101085 106287 101113
rect 106321 101085 106349 101113
rect 106259 101023 106287 101051
rect 106321 101023 106349 101051
rect 106259 100961 106287 100989
rect 106321 100961 106349 100989
rect 111485 122147 111513 122175
rect 111547 122147 111575 122175
rect 111609 122147 111637 122175
rect 111671 122147 111699 122175
rect 111485 122085 111513 122113
rect 111547 122085 111575 122113
rect 111609 122085 111637 122113
rect 111671 122085 111699 122113
rect 111485 122023 111513 122051
rect 111547 122023 111575 122051
rect 111609 122023 111637 122051
rect 111671 122023 111699 122051
rect 111485 121961 111513 121989
rect 111547 121961 111575 121989
rect 111609 121961 111637 121989
rect 111671 121961 111699 121989
rect 111485 113147 111513 113175
rect 111547 113147 111575 113175
rect 111609 113147 111637 113175
rect 111671 113147 111699 113175
rect 111485 113085 111513 113113
rect 111547 113085 111575 113113
rect 111609 113085 111637 113113
rect 111671 113085 111699 113113
rect 111485 113023 111513 113051
rect 111547 113023 111575 113051
rect 111609 113023 111637 113051
rect 111671 113023 111699 113051
rect 111485 112961 111513 112989
rect 111547 112961 111575 112989
rect 111609 112961 111637 112989
rect 111671 112961 111699 112989
rect 118625 119147 118653 119175
rect 118687 119147 118715 119175
rect 118749 119147 118777 119175
rect 118811 119147 118839 119175
rect 118625 119085 118653 119113
rect 118687 119085 118715 119113
rect 118749 119085 118777 119113
rect 118811 119085 118839 119113
rect 118625 119023 118653 119051
rect 118687 119023 118715 119051
rect 118749 119023 118777 119051
rect 118811 119023 118839 119051
rect 118625 118961 118653 118989
rect 118687 118961 118715 118989
rect 118749 118961 118777 118989
rect 118811 118961 118839 118989
rect 118625 110147 118653 110175
rect 118687 110147 118715 110175
rect 118749 110147 118777 110175
rect 118811 110147 118839 110175
rect 118625 110085 118653 110113
rect 118687 110085 118715 110113
rect 118749 110085 118777 110113
rect 118811 110085 118839 110113
rect 118625 110023 118653 110051
rect 118687 110023 118715 110051
rect 118749 110023 118777 110051
rect 118811 110023 118839 110051
rect 118625 109961 118653 109989
rect 118687 109961 118715 109989
rect 118749 109961 118777 109989
rect 118811 109961 118839 109989
rect 111485 104147 111513 104175
rect 111547 104147 111575 104175
rect 111609 104147 111637 104175
rect 111671 104147 111699 104175
rect 111485 104085 111513 104113
rect 111547 104085 111575 104113
rect 111609 104085 111637 104113
rect 111671 104085 111699 104113
rect 111485 104023 111513 104051
rect 111547 104023 111575 104051
rect 111609 104023 111637 104051
rect 111671 104023 111699 104051
rect 111485 103961 111513 103989
rect 111547 103961 111575 103989
rect 111609 103961 111637 103989
rect 111671 103961 111699 103989
rect 109625 101147 109653 101175
rect 109687 101147 109715 101175
rect 109749 101147 109777 101175
rect 109811 101147 109839 101175
rect 109625 101085 109653 101113
rect 109687 101085 109715 101113
rect 109749 101085 109777 101113
rect 109811 101085 109839 101113
rect 109625 101023 109653 101051
rect 109687 101023 109715 101051
rect 109749 101023 109777 101051
rect 109811 101023 109839 101051
rect 109625 100961 109653 100989
rect 109687 100961 109715 100989
rect 109749 100961 109777 100989
rect 109811 100961 109839 100989
rect 110759 101147 110787 101175
rect 110821 101147 110849 101175
rect 110759 101085 110787 101113
rect 110821 101085 110849 101113
rect 110759 101023 110787 101051
rect 110821 101023 110849 101051
rect 110759 100961 110787 100989
rect 110821 100961 110849 100989
rect 113009 104147 113037 104175
rect 113071 104147 113099 104175
rect 113009 104085 113037 104113
rect 113071 104085 113099 104113
rect 113009 104023 113037 104051
rect 113071 104023 113099 104051
rect 113009 103961 113037 103989
rect 113071 103961 113099 103989
rect 117509 104147 117537 104175
rect 117571 104147 117599 104175
rect 117509 104085 117537 104113
rect 117571 104085 117599 104113
rect 117509 104023 117537 104051
rect 117571 104023 117599 104051
rect 117509 103961 117537 103989
rect 117571 103961 117599 103989
rect 115259 101147 115287 101175
rect 115321 101147 115349 101175
rect 115259 101085 115287 101113
rect 115321 101085 115349 101113
rect 115259 101023 115287 101051
rect 115321 101023 115349 101051
rect 115259 100961 115287 100989
rect 115321 100961 115349 100989
rect 118625 101147 118653 101175
rect 118687 101147 118715 101175
rect 118749 101147 118777 101175
rect 118811 101147 118839 101175
rect 118625 101085 118653 101113
rect 118687 101085 118715 101113
rect 118749 101085 118777 101113
rect 118811 101085 118839 101113
rect 118625 101023 118653 101051
rect 118687 101023 118715 101051
rect 118749 101023 118777 101051
rect 118811 101023 118839 101051
rect 118625 100961 118653 100989
rect 118687 100961 118715 100989
rect 118749 100961 118777 100989
rect 118811 100961 118839 100989
rect 120485 122147 120513 122175
rect 120547 122147 120575 122175
rect 120609 122147 120637 122175
rect 120671 122147 120699 122175
rect 120485 122085 120513 122113
rect 120547 122085 120575 122113
rect 120609 122085 120637 122113
rect 120671 122085 120699 122113
rect 120485 122023 120513 122051
rect 120547 122023 120575 122051
rect 120609 122023 120637 122051
rect 120671 122023 120699 122051
rect 120485 121961 120513 121989
rect 120547 121961 120575 121989
rect 120609 121961 120637 121989
rect 120671 121961 120699 121989
rect 120485 113147 120513 113175
rect 120547 113147 120575 113175
rect 120609 113147 120637 113175
rect 120671 113147 120699 113175
rect 120485 113085 120513 113113
rect 120547 113085 120575 113113
rect 120609 113085 120637 113113
rect 120671 113085 120699 113113
rect 120485 113023 120513 113051
rect 120547 113023 120575 113051
rect 120609 113023 120637 113051
rect 120671 113023 120699 113051
rect 120485 112961 120513 112989
rect 120547 112961 120575 112989
rect 120609 112961 120637 112989
rect 120671 112961 120699 112989
rect 120485 104147 120513 104175
rect 120547 104147 120575 104175
rect 120609 104147 120637 104175
rect 120671 104147 120699 104175
rect 120485 104085 120513 104113
rect 120547 104085 120575 104113
rect 120609 104085 120637 104113
rect 120671 104085 120699 104113
rect 120485 104023 120513 104051
rect 120547 104023 120575 104051
rect 120609 104023 120637 104051
rect 120671 104023 120699 104051
rect 120485 103961 120513 103989
rect 120547 103961 120575 103989
rect 120609 103961 120637 103989
rect 120671 103961 120699 103989
rect 95009 95147 95037 95175
rect 95071 95147 95099 95175
rect 95009 95085 95037 95113
rect 95071 95085 95099 95113
rect 95009 95023 95037 95051
rect 95071 95023 95099 95051
rect 95009 94961 95037 94989
rect 95071 94961 95099 94989
rect 99509 95147 99537 95175
rect 99571 95147 99599 95175
rect 99509 95085 99537 95113
rect 99571 95085 99599 95113
rect 99509 95023 99537 95051
rect 99571 95023 99599 95051
rect 99509 94961 99537 94989
rect 99571 94961 99599 94989
rect 104009 95147 104037 95175
rect 104071 95147 104099 95175
rect 104009 95085 104037 95113
rect 104071 95085 104099 95113
rect 104009 95023 104037 95051
rect 104071 95023 104099 95051
rect 104009 94961 104037 94989
rect 104071 94961 104099 94989
rect 108509 95147 108537 95175
rect 108571 95147 108599 95175
rect 108509 95085 108537 95113
rect 108571 95085 108599 95113
rect 108509 95023 108537 95051
rect 108571 95023 108599 95051
rect 108509 94961 108537 94989
rect 108571 94961 108599 94989
rect 113009 95147 113037 95175
rect 113071 95147 113099 95175
rect 113009 95085 113037 95113
rect 113071 95085 113099 95113
rect 113009 95023 113037 95051
rect 113071 95023 113099 95051
rect 113009 94961 113037 94989
rect 113071 94961 113099 94989
rect 117509 95147 117537 95175
rect 117571 95147 117599 95175
rect 117509 95085 117537 95113
rect 117571 95085 117599 95113
rect 117509 95023 117537 95051
rect 117571 95023 117599 95051
rect 117509 94961 117537 94989
rect 117571 94961 117599 94989
rect 120485 95147 120513 95175
rect 120547 95147 120575 95175
rect 120609 95147 120637 95175
rect 120671 95147 120699 95175
rect 120485 95085 120513 95113
rect 120547 95085 120575 95113
rect 120609 95085 120637 95113
rect 120671 95085 120699 95113
rect 120485 95023 120513 95051
rect 120547 95023 120575 95051
rect 120609 95023 120637 95051
rect 120671 95023 120699 95051
rect 120485 94961 120513 94989
rect 120547 94961 120575 94989
rect 120609 94961 120637 94989
rect 120671 94961 120699 94989
rect 91625 92147 91653 92175
rect 91687 92147 91715 92175
rect 91749 92147 91777 92175
rect 91811 92147 91839 92175
rect 91625 92085 91653 92113
rect 91687 92085 91715 92113
rect 91749 92085 91777 92113
rect 91811 92085 91839 92113
rect 91625 92023 91653 92051
rect 91687 92023 91715 92051
rect 91749 92023 91777 92051
rect 91811 92023 91839 92051
rect 91625 91961 91653 91989
rect 91687 91961 91715 91989
rect 91749 91961 91777 91989
rect 91811 91961 91839 91989
rect 84485 86147 84513 86175
rect 84547 86147 84575 86175
rect 84609 86147 84637 86175
rect 84671 86147 84699 86175
rect 84485 86085 84513 86113
rect 84547 86085 84575 86113
rect 84609 86085 84637 86113
rect 84671 86085 84699 86113
rect 84485 86023 84513 86051
rect 84547 86023 84575 86051
rect 84609 86023 84637 86051
rect 84671 86023 84699 86051
rect 84485 85961 84513 85989
rect 84547 85961 84575 85989
rect 84609 85961 84637 85989
rect 84671 85961 84699 85989
rect 82625 83147 82653 83175
rect 82687 83147 82715 83175
rect 82749 83147 82777 83175
rect 82811 83147 82839 83175
rect 82625 83085 82653 83113
rect 82687 83085 82715 83113
rect 82749 83085 82777 83113
rect 82811 83085 82839 83113
rect 82625 83023 82653 83051
rect 82687 83023 82715 83051
rect 82749 83023 82777 83051
rect 82811 83023 82839 83051
rect 82625 82961 82653 82989
rect 82687 82961 82715 82989
rect 82749 82961 82777 82989
rect 82811 82961 82839 82989
rect 75485 77147 75513 77175
rect 75547 77147 75575 77175
rect 75609 77147 75637 77175
rect 75671 77147 75699 77175
rect 75485 77085 75513 77113
rect 75547 77085 75575 77113
rect 75609 77085 75637 77113
rect 75671 77085 75699 77113
rect 75485 77023 75513 77051
rect 75547 77023 75575 77051
rect 75609 77023 75637 77051
rect 75671 77023 75699 77051
rect 75485 76961 75513 76989
rect 75547 76961 75575 76989
rect 75609 76961 75637 76989
rect 75671 76961 75699 76989
rect 73625 74147 73653 74175
rect 73687 74147 73715 74175
rect 73749 74147 73777 74175
rect 73811 74147 73839 74175
rect 73625 74085 73653 74113
rect 73687 74085 73715 74113
rect 73749 74085 73777 74113
rect 73811 74085 73839 74113
rect 73625 74023 73653 74051
rect 73687 74023 73715 74051
rect 73749 74023 73777 74051
rect 73811 74023 73839 74051
rect 73625 73961 73653 73989
rect 73687 73961 73715 73989
rect 73749 73961 73777 73989
rect 73811 73961 73839 73989
rect 66485 68147 66513 68175
rect 66547 68147 66575 68175
rect 66609 68147 66637 68175
rect 66671 68147 66699 68175
rect 66485 68085 66513 68113
rect 66547 68085 66575 68113
rect 66609 68085 66637 68113
rect 66671 68085 66699 68113
rect 66485 68023 66513 68051
rect 66547 68023 66575 68051
rect 66609 68023 66637 68051
rect 66671 68023 66699 68051
rect 66485 67961 66513 67989
rect 66547 67961 66575 67989
rect 66609 67961 66637 67989
rect 66671 67961 66699 67989
rect 64625 65147 64653 65175
rect 64687 65147 64715 65175
rect 64749 65147 64777 65175
rect 64811 65147 64839 65175
rect 64625 65085 64653 65113
rect 64687 65085 64715 65113
rect 64749 65085 64777 65113
rect 64811 65085 64839 65113
rect 64625 65023 64653 65051
rect 64687 65023 64715 65051
rect 64749 65023 64777 65051
rect 64811 65023 64839 65051
rect 64625 64961 64653 64989
rect 64687 64961 64715 64989
rect 64749 64961 64777 64989
rect 64811 64961 64839 64989
rect 57485 59147 57513 59175
rect 57547 59147 57575 59175
rect 57609 59147 57637 59175
rect 57671 59147 57699 59175
rect 57485 59085 57513 59113
rect 57547 59085 57575 59113
rect 57609 59085 57637 59113
rect 57671 59085 57699 59113
rect 57485 59023 57513 59051
rect 57547 59023 57575 59051
rect 57609 59023 57637 59051
rect 57671 59023 57699 59051
rect 57485 58961 57513 58989
rect 57547 58961 57575 58989
rect 57609 58961 57637 58989
rect 57671 58961 57699 58989
rect 55625 56147 55653 56175
rect 55687 56147 55715 56175
rect 55749 56147 55777 56175
rect 55811 56147 55839 56175
rect 55625 56085 55653 56113
rect 55687 56085 55715 56113
rect 55749 56085 55777 56113
rect 55811 56085 55839 56113
rect 55625 56023 55653 56051
rect 55687 56023 55715 56051
rect 55749 56023 55777 56051
rect 55811 56023 55839 56051
rect 55625 55961 55653 55989
rect 55687 55961 55715 55989
rect 55749 55961 55777 55989
rect 55811 55961 55839 55989
rect 48485 50147 48513 50175
rect 48547 50147 48575 50175
rect 48609 50147 48637 50175
rect 48671 50147 48699 50175
rect 48485 50085 48513 50113
rect 48547 50085 48575 50113
rect 48609 50085 48637 50113
rect 48671 50085 48699 50113
rect 48485 50023 48513 50051
rect 48547 50023 48575 50051
rect 48609 50023 48637 50051
rect 48671 50023 48699 50051
rect 48485 49961 48513 49989
rect 48547 49961 48575 49989
rect 48609 49961 48637 49989
rect 48671 49961 48699 49989
rect 48485 41147 48513 41175
rect 48547 41147 48575 41175
rect 48609 41147 48637 41175
rect 48671 41147 48699 41175
rect 48485 41085 48513 41113
rect 48547 41085 48575 41113
rect 48609 41085 48637 41113
rect 48671 41085 48699 41113
rect 48485 41023 48513 41051
rect 48547 41023 48575 41051
rect 48609 41023 48637 41051
rect 48671 41023 48699 41051
rect 48485 40961 48513 40989
rect 48547 40961 48575 40989
rect 48609 40961 48637 40989
rect 48671 40961 48699 40989
rect 48485 32147 48513 32175
rect 48547 32147 48575 32175
rect 48609 32147 48637 32175
rect 48671 32147 48699 32175
rect 48485 32085 48513 32113
rect 48547 32085 48575 32113
rect 48609 32085 48637 32113
rect 48671 32085 48699 32113
rect 48485 32023 48513 32051
rect 48547 32023 48575 32051
rect 48609 32023 48637 32051
rect 48671 32023 48699 32051
rect 48485 31961 48513 31989
rect 48547 31961 48575 31989
rect 48609 31961 48637 31989
rect 48671 31961 48699 31989
rect 48485 23147 48513 23175
rect 48547 23147 48575 23175
rect 48609 23147 48637 23175
rect 48671 23147 48699 23175
rect 48485 23085 48513 23113
rect 48547 23085 48575 23113
rect 48609 23085 48637 23113
rect 48671 23085 48699 23113
rect 48485 23023 48513 23051
rect 48547 23023 48575 23051
rect 48609 23023 48637 23051
rect 48671 23023 48699 23051
rect 48485 22961 48513 22989
rect 48547 22961 48575 22989
rect 48609 22961 48637 22989
rect 48671 22961 48699 22989
rect 48485 14147 48513 14175
rect 48547 14147 48575 14175
rect 48609 14147 48637 14175
rect 48671 14147 48699 14175
rect 48485 14085 48513 14113
rect 48547 14085 48575 14113
rect 48609 14085 48637 14113
rect 48671 14085 48699 14113
rect 48485 14023 48513 14051
rect 48547 14023 48575 14051
rect 48609 14023 48637 14051
rect 48671 14023 48699 14051
rect 48485 13961 48513 13989
rect 48547 13961 48575 13989
rect 48609 13961 48637 13989
rect 48671 13961 48699 13989
rect 48485 5147 48513 5175
rect 48547 5147 48575 5175
rect 48609 5147 48637 5175
rect 48671 5147 48699 5175
rect 48485 5085 48513 5113
rect 48547 5085 48575 5113
rect 48609 5085 48637 5113
rect 48671 5085 48699 5113
rect 48485 5023 48513 5051
rect 48547 5023 48575 5051
rect 48609 5023 48637 5051
rect 48671 5023 48699 5051
rect 48485 4961 48513 4989
rect 48547 4961 48575 4989
rect 48609 4961 48637 4989
rect 48671 4961 48699 4989
rect 48485 -588 48513 -560
rect 48547 -588 48575 -560
rect 48609 -588 48637 -560
rect 48671 -588 48699 -560
rect 48485 -650 48513 -622
rect 48547 -650 48575 -622
rect 48609 -650 48637 -622
rect 48671 -650 48699 -622
rect 48485 -712 48513 -684
rect 48547 -712 48575 -684
rect 48609 -712 48637 -684
rect 48671 -712 48699 -684
rect 48485 -774 48513 -746
rect 48547 -774 48575 -746
rect 48609 -774 48637 -746
rect 48671 -774 48699 -746
rect 56759 56147 56787 56175
rect 56821 56147 56849 56175
rect 56759 56085 56787 56113
rect 56821 56085 56849 56113
rect 56759 56023 56787 56051
rect 56821 56023 56849 56051
rect 56759 55961 56787 55989
rect 56821 55961 56849 55989
rect 55625 47147 55653 47175
rect 55687 47147 55715 47175
rect 55749 47147 55777 47175
rect 55811 47147 55839 47175
rect 55625 47085 55653 47113
rect 55687 47085 55715 47113
rect 55749 47085 55777 47113
rect 55811 47085 55839 47113
rect 55625 47023 55653 47051
rect 55687 47023 55715 47051
rect 55749 47023 55777 47051
rect 55811 47023 55839 47051
rect 55625 46961 55653 46989
rect 55687 46961 55715 46989
rect 55749 46961 55777 46989
rect 55811 46961 55839 46989
rect 55625 38147 55653 38175
rect 55687 38147 55715 38175
rect 55749 38147 55777 38175
rect 55811 38147 55839 38175
rect 55625 38085 55653 38113
rect 55687 38085 55715 38113
rect 55749 38085 55777 38113
rect 55811 38085 55839 38113
rect 55625 38023 55653 38051
rect 55687 38023 55715 38051
rect 55749 38023 55777 38051
rect 55811 38023 55839 38051
rect 55625 37961 55653 37989
rect 55687 37961 55715 37989
rect 55749 37961 55777 37989
rect 55811 37961 55839 37989
rect 55625 29147 55653 29175
rect 55687 29147 55715 29175
rect 55749 29147 55777 29175
rect 55811 29147 55839 29175
rect 55625 29085 55653 29113
rect 55687 29085 55715 29113
rect 55749 29085 55777 29113
rect 55811 29085 55839 29113
rect 55625 29023 55653 29051
rect 55687 29023 55715 29051
rect 55749 29023 55777 29051
rect 55811 29023 55839 29051
rect 55625 28961 55653 28989
rect 55687 28961 55715 28989
rect 55749 28961 55777 28989
rect 55811 28961 55839 28989
rect 55625 20147 55653 20175
rect 55687 20147 55715 20175
rect 55749 20147 55777 20175
rect 55811 20147 55839 20175
rect 55625 20085 55653 20113
rect 55687 20085 55715 20113
rect 55749 20085 55777 20113
rect 55811 20085 55839 20113
rect 55625 20023 55653 20051
rect 55687 20023 55715 20051
rect 55749 20023 55777 20051
rect 55811 20023 55839 20051
rect 55625 19961 55653 19989
rect 55687 19961 55715 19989
rect 55749 19961 55777 19989
rect 55811 19961 55839 19989
rect 55625 11147 55653 11175
rect 55687 11147 55715 11175
rect 55749 11147 55777 11175
rect 55811 11147 55839 11175
rect 55625 11085 55653 11113
rect 55687 11085 55715 11113
rect 55749 11085 55777 11113
rect 55811 11085 55839 11113
rect 55625 11023 55653 11051
rect 55687 11023 55715 11051
rect 55749 11023 55777 11051
rect 55811 11023 55839 11051
rect 55625 10961 55653 10989
rect 55687 10961 55715 10989
rect 55749 10961 55777 10989
rect 55811 10961 55839 10989
rect 55625 2147 55653 2175
rect 55687 2147 55715 2175
rect 55749 2147 55777 2175
rect 55811 2147 55839 2175
rect 55625 2085 55653 2113
rect 55687 2085 55715 2113
rect 55749 2085 55777 2113
rect 55811 2085 55839 2113
rect 55625 2023 55653 2051
rect 55687 2023 55715 2051
rect 55749 2023 55777 2051
rect 55811 2023 55839 2051
rect 55625 1961 55653 1989
rect 55687 1961 55715 1989
rect 55749 1961 55777 1989
rect 55811 1961 55839 1989
rect 55625 -108 55653 -80
rect 55687 -108 55715 -80
rect 55749 -108 55777 -80
rect 55811 -108 55839 -80
rect 55625 -170 55653 -142
rect 55687 -170 55715 -142
rect 55749 -170 55777 -142
rect 55811 -170 55839 -142
rect 55625 -232 55653 -204
rect 55687 -232 55715 -204
rect 55749 -232 55777 -204
rect 55811 -232 55839 -204
rect 55625 -294 55653 -266
rect 55687 -294 55715 -266
rect 55749 -294 55777 -266
rect 55811 -294 55839 -266
rect 59009 59147 59037 59175
rect 59071 59147 59099 59175
rect 59009 59085 59037 59113
rect 59071 59085 59099 59113
rect 59009 59023 59037 59051
rect 59071 59023 59099 59051
rect 59009 58961 59037 58989
rect 59071 58961 59099 58989
rect 63509 59147 63537 59175
rect 63571 59147 63599 59175
rect 63509 59085 63537 59113
rect 63571 59085 63599 59113
rect 63509 59023 63537 59051
rect 63571 59023 63599 59051
rect 63509 58961 63537 58989
rect 63571 58961 63599 58989
rect 61259 56147 61287 56175
rect 61321 56147 61349 56175
rect 61259 56085 61287 56113
rect 61321 56085 61349 56113
rect 61259 56023 61287 56051
rect 61321 56023 61349 56051
rect 61259 55961 61287 55989
rect 61321 55961 61349 55989
rect 65759 65147 65787 65175
rect 65821 65147 65849 65175
rect 65759 65085 65787 65113
rect 65821 65085 65849 65113
rect 65759 65023 65787 65051
rect 65821 65023 65849 65051
rect 65759 64961 65787 64989
rect 65821 64961 65849 64989
rect 68009 68147 68037 68175
rect 68071 68147 68099 68175
rect 68009 68085 68037 68113
rect 68071 68085 68099 68113
rect 68009 68023 68037 68051
rect 68071 68023 68099 68051
rect 68009 67961 68037 67989
rect 68071 67961 68099 67989
rect 72509 68147 72537 68175
rect 72571 68147 72599 68175
rect 72509 68085 72537 68113
rect 72571 68085 72599 68113
rect 72509 68023 72537 68051
rect 72571 68023 72599 68051
rect 72509 67961 72537 67989
rect 72571 67961 72599 67989
rect 70259 65147 70287 65175
rect 70321 65147 70349 65175
rect 70259 65085 70287 65113
rect 70321 65085 70349 65113
rect 70259 65023 70287 65051
rect 70321 65023 70349 65051
rect 70259 64961 70287 64989
rect 70321 64961 70349 64989
rect 74759 74147 74787 74175
rect 74821 74147 74849 74175
rect 74759 74085 74787 74113
rect 74821 74085 74849 74113
rect 74759 74023 74787 74051
rect 74821 74023 74849 74051
rect 74759 73961 74787 73989
rect 74821 73961 74849 73989
rect 77009 77147 77037 77175
rect 77071 77147 77099 77175
rect 77009 77085 77037 77113
rect 77071 77085 77099 77113
rect 77009 77023 77037 77051
rect 77071 77023 77099 77051
rect 77009 76961 77037 76989
rect 77071 76961 77099 76989
rect 81509 77147 81537 77175
rect 81571 77147 81599 77175
rect 81509 77085 81537 77113
rect 81571 77085 81599 77113
rect 81509 77023 81537 77051
rect 81571 77023 81599 77051
rect 81509 76961 81537 76989
rect 81571 76961 81599 76989
rect 79259 74147 79287 74175
rect 79321 74147 79349 74175
rect 79259 74085 79287 74113
rect 79321 74085 79349 74113
rect 79259 74023 79287 74051
rect 79321 74023 79349 74051
rect 79259 73961 79287 73989
rect 79321 73961 79349 73989
rect 83759 83147 83787 83175
rect 83821 83147 83849 83175
rect 83759 83085 83787 83113
rect 83821 83085 83849 83113
rect 83759 83023 83787 83051
rect 83821 83023 83849 83051
rect 83759 82961 83787 82989
rect 83821 82961 83849 82989
rect 86009 86147 86037 86175
rect 86071 86147 86099 86175
rect 86009 86085 86037 86113
rect 86071 86085 86099 86113
rect 86009 86023 86037 86051
rect 86071 86023 86099 86051
rect 86009 85961 86037 85989
rect 86071 85961 86099 85989
rect 90509 86147 90537 86175
rect 90571 86147 90599 86175
rect 90509 86085 90537 86113
rect 90571 86085 90599 86113
rect 90509 86023 90537 86051
rect 90571 86023 90599 86051
rect 90509 85961 90537 85989
rect 90571 85961 90599 85989
rect 88259 83147 88287 83175
rect 88321 83147 88349 83175
rect 88259 83085 88287 83113
rect 88321 83085 88349 83113
rect 88259 83023 88287 83051
rect 88321 83023 88349 83051
rect 88259 82961 88287 82989
rect 88321 82961 88349 82989
rect 92759 92147 92787 92175
rect 92821 92147 92849 92175
rect 92759 92085 92787 92113
rect 92821 92085 92849 92113
rect 92759 92023 92787 92051
rect 92821 92023 92849 92051
rect 92759 91961 92787 91989
rect 92821 91961 92849 91989
rect 97259 92147 97287 92175
rect 97321 92147 97349 92175
rect 97259 92085 97287 92113
rect 97321 92085 97349 92113
rect 97259 92023 97287 92051
rect 97321 92023 97349 92051
rect 97259 91961 97287 91989
rect 97321 91961 97349 91989
rect 101759 92147 101787 92175
rect 101821 92147 101849 92175
rect 101759 92085 101787 92113
rect 101821 92085 101849 92113
rect 101759 92023 101787 92051
rect 101821 92023 101849 92051
rect 101759 91961 101787 91989
rect 101821 91961 101849 91989
rect 106259 92147 106287 92175
rect 106321 92147 106349 92175
rect 106259 92085 106287 92113
rect 106321 92085 106349 92113
rect 106259 92023 106287 92051
rect 106321 92023 106349 92051
rect 106259 91961 106287 91989
rect 106321 91961 106349 91989
rect 110759 92147 110787 92175
rect 110821 92147 110849 92175
rect 110759 92085 110787 92113
rect 110821 92085 110849 92113
rect 110759 92023 110787 92051
rect 110821 92023 110849 92051
rect 110759 91961 110787 91989
rect 110821 91961 110849 91989
rect 115259 92147 115287 92175
rect 115321 92147 115349 92175
rect 115259 92085 115287 92113
rect 115321 92085 115349 92113
rect 115259 92023 115287 92051
rect 115321 92023 115349 92051
rect 115259 91961 115287 91989
rect 115321 91961 115349 91989
rect 95009 86147 95037 86175
rect 95071 86147 95099 86175
rect 95009 86085 95037 86113
rect 95071 86085 95099 86113
rect 95009 86023 95037 86051
rect 95071 86023 95099 86051
rect 95009 85961 95037 85989
rect 95071 85961 95099 85989
rect 99509 86147 99537 86175
rect 99571 86147 99599 86175
rect 99509 86085 99537 86113
rect 99571 86085 99599 86113
rect 99509 86023 99537 86051
rect 99571 86023 99599 86051
rect 99509 85961 99537 85989
rect 99571 85961 99599 85989
rect 104009 86147 104037 86175
rect 104071 86147 104099 86175
rect 104009 86085 104037 86113
rect 104071 86085 104099 86113
rect 104009 86023 104037 86051
rect 104071 86023 104099 86051
rect 104009 85961 104037 85989
rect 104071 85961 104099 85989
rect 108509 86147 108537 86175
rect 108571 86147 108599 86175
rect 108509 86085 108537 86113
rect 108571 86085 108599 86113
rect 108509 86023 108537 86051
rect 108571 86023 108599 86051
rect 108509 85961 108537 85989
rect 108571 85961 108599 85989
rect 113009 86147 113037 86175
rect 113071 86147 113099 86175
rect 113009 86085 113037 86113
rect 113071 86085 113099 86113
rect 113009 86023 113037 86051
rect 113071 86023 113099 86051
rect 113009 85961 113037 85989
rect 113071 85961 113099 85989
rect 117509 86147 117537 86175
rect 117571 86147 117599 86175
rect 117509 86085 117537 86113
rect 117571 86085 117599 86113
rect 117509 86023 117537 86051
rect 117571 86023 117599 86051
rect 117509 85961 117537 85989
rect 117571 85961 117599 85989
rect 120485 86147 120513 86175
rect 120547 86147 120575 86175
rect 120609 86147 120637 86175
rect 120671 86147 120699 86175
rect 120485 86085 120513 86113
rect 120547 86085 120575 86113
rect 120609 86085 120637 86113
rect 120671 86085 120699 86113
rect 120485 86023 120513 86051
rect 120547 86023 120575 86051
rect 120609 86023 120637 86051
rect 120671 86023 120699 86051
rect 120485 85961 120513 85989
rect 120547 85961 120575 85989
rect 120609 85961 120637 85989
rect 120671 85961 120699 85989
rect 91625 83147 91653 83175
rect 91687 83147 91715 83175
rect 91749 83147 91777 83175
rect 91811 83147 91839 83175
rect 91625 83085 91653 83113
rect 91687 83085 91715 83113
rect 91749 83085 91777 83113
rect 91811 83085 91839 83113
rect 91625 83023 91653 83051
rect 91687 83023 91715 83051
rect 91749 83023 91777 83051
rect 91811 83023 91839 83051
rect 91625 82961 91653 82989
rect 91687 82961 91715 82989
rect 91749 82961 91777 82989
rect 91811 82961 91839 82989
rect 84485 77147 84513 77175
rect 84547 77147 84575 77175
rect 84609 77147 84637 77175
rect 84671 77147 84699 77175
rect 84485 77085 84513 77113
rect 84547 77085 84575 77113
rect 84609 77085 84637 77113
rect 84671 77085 84699 77113
rect 84485 77023 84513 77051
rect 84547 77023 84575 77051
rect 84609 77023 84637 77051
rect 84671 77023 84699 77051
rect 84485 76961 84513 76989
rect 84547 76961 84575 76989
rect 84609 76961 84637 76989
rect 84671 76961 84699 76989
rect 82625 74147 82653 74175
rect 82687 74147 82715 74175
rect 82749 74147 82777 74175
rect 82811 74147 82839 74175
rect 82625 74085 82653 74113
rect 82687 74085 82715 74113
rect 82749 74085 82777 74113
rect 82811 74085 82839 74113
rect 82625 74023 82653 74051
rect 82687 74023 82715 74051
rect 82749 74023 82777 74051
rect 82811 74023 82839 74051
rect 82625 73961 82653 73989
rect 82687 73961 82715 73989
rect 82749 73961 82777 73989
rect 82811 73961 82839 73989
rect 75485 68147 75513 68175
rect 75547 68147 75575 68175
rect 75609 68147 75637 68175
rect 75671 68147 75699 68175
rect 75485 68085 75513 68113
rect 75547 68085 75575 68113
rect 75609 68085 75637 68113
rect 75671 68085 75699 68113
rect 75485 68023 75513 68051
rect 75547 68023 75575 68051
rect 75609 68023 75637 68051
rect 75671 68023 75699 68051
rect 75485 67961 75513 67989
rect 75547 67961 75575 67989
rect 75609 67961 75637 67989
rect 75671 67961 75699 67989
rect 73625 65147 73653 65175
rect 73687 65147 73715 65175
rect 73749 65147 73777 65175
rect 73811 65147 73839 65175
rect 73625 65085 73653 65113
rect 73687 65085 73715 65113
rect 73749 65085 73777 65113
rect 73811 65085 73839 65113
rect 73625 65023 73653 65051
rect 73687 65023 73715 65051
rect 73749 65023 73777 65051
rect 73811 65023 73839 65051
rect 73625 64961 73653 64989
rect 73687 64961 73715 64989
rect 73749 64961 73777 64989
rect 73811 64961 73839 64989
rect 66485 59147 66513 59175
rect 66547 59147 66575 59175
rect 66609 59147 66637 59175
rect 66671 59147 66699 59175
rect 66485 59085 66513 59113
rect 66547 59085 66575 59113
rect 66609 59085 66637 59113
rect 66671 59085 66699 59113
rect 66485 59023 66513 59051
rect 66547 59023 66575 59051
rect 66609 59023 66637 59051
rect 66671 59023 66699 59051
rect 66485 58961 66513 58989
rect 66547 58961 66575 58989
rect 66609 58961 66637 58989
rect 66671 58961 66699 58989
rect 64625 56147 64653 56175
rect 64687 56147 64715 56175
rect 64749 56147 64777 56175
rect 64811 56147 64839 56175
rect 64625 56085 64653 56113
rect 64687 56085 64715 56113
rect 64749 56085 64777 56113
rect 64811 56085 64839 56113
rect 64625 56023 64653 56051
rect 64687 56023 64715 56051
rect 64749 56023 64777 56051
rect 64811 56023 64839 56051
rect 64625 55961 64653 55989
rect 64687 55961 64715 55989
rect 64749 55961 64777 55989
rect 64811 55961 64839 55989
rect 57485 50147 57513 50175
rect 57547 50147 57575 50175
rect 57609 50147 57637 50175
rect 57671 50147 57699 50175
rect 57485 50085 57513 50113
rect 57547 50085 57575 50113
rect 57609 50085 57637 50113
rect 57671 50085 57699 50113
rect 57485 50023 57513 50051
rect 57547 50023 57575 50051
rect 57609 50023 57637 50051
rect 57671 50023 57699 50051
rect 57485 49961 57513 49989
rect 57547 49961 57575 49989
rect 57609 49961 57637 49989
rect 57671 49961 57699 49989
rect 57485 41147 57513 41175
rect 57547 41147 57575 41175
rect 57609 41147 57637 41175
rect 57671 41147 57699 41175
rect 57485 41085 57513 41113
rect 57547 41085 57575 41113
rect 57609 41085 57637 41113
rect 57671 41085 57699 41113
rect 57485 41023 57513 41051
rect 57547 41023 57575 41051
rect 57609 41023 57637 41051
rect 57671 41023 57699 41051
rect 57485 40961 57513 40989
rect 57547 40961 57575 40989
rect 57609 40961 57637 40989
rect 57671 40961 57699 40989
rect 57485 32147 57513 32175
rect 57547 32147 57575 32175
rect 57609 32147 57637 32175
rect 57671 32147 57699 32175
rect 57485 32085 57513 32113
rect 57547 32085 57575 32113
rect 57609 32085 57637 32113
rect 57671 32085 57699 32113
rect 57485 32023 57513 32051
rect 57547 32023 57575 32051
rect 57609 32023 57637 32051
rect 57671 32023 57699 32051
rect 57485 31961 57513 31989
rect 57547 31961 57575 31989
rect 57609 31961 57637 31989
rect 57671 31961 57699 31989
rect 57485 23147 57513 23175
rect 57547 23147 57575 23175
rect 57609 23147 57637 23175
rect 57671 23147 57699 23175
rect 57485 23085 57513 23113
rect 57547 23085 57575 23113
rect 57609 23085 57637 23113
rect 57671 23085 57699 23113
rect 57485 23023 57513 23051
rect 57547 23023 57575 23051
rect 57609 23023 57637 23051
rect 57671 23023 57699 23051
rect 57485 22961 57513 22989
rect 57547 22961 57575 22989
rect 57609 22961 57637 22989
rect 57671 22961 57699 22989
rect 57485 14147 57513 14175
rect 57547 14147 57575 14175
rect 57609 14147 57637 14175
rect 57671 14147 57699 14175
rect 57485 14085 57513 14113
rect 57547 14085 57575 14113
rect 57609 14085 57637 14113
rect 57671 14085 57699 14113
rect 57485 14023 57513 14051
rect 57547 14023 57575 14051
rect 57609 14023 57637 14051
rect 57671 14023 57699 14051
rect 57485 13961 57513 13989
rect 57547 13961 57575 13989
rect 57609 13961 57637 13989
rect 57671 13961 57699 13989
rect 57485 5147 57513 5175
rect 57547 5147 57575 5175
rect 57609 5147 57637 5175
rect 57671 5147 57699 5175
rect 57485 5085 57513 5113
rect 57547 5085 57575 5113
rect 57609 5085 57637 5113
rect 57671 5085 57699 5113
rect 57485 5023 57513 5051
rect 57547 5023 57575 5051
rect 57609 5023 57637 5051
rect 57671 5023 57699 5051
rect 57485 4961 57513 4989
rect 57547 4961 57575 4989
rect 57609 4961 57637 4989
rect 57671 4961 57699 4989
rect 57485 -588 57513 -560
rect 57547 -588 57575 -560
rect 57609 -588 57637 -560
rect 57671 -588 57699 -560
rect 57485 -650 57513 -622
rect 57547 -650 57575 -622
rect 57609 -650 57637 -622
rect 57671 -650 57699 -622
rect 57485 -712 57513 -684
rect 57547 -712 57575 -684
rect 57609 -712 57637 -684
rect 57671 -712 57699 -684
rect 57485 -774 57513 -746
rect 57547 -774 57575 -746
rect 57609 -774 57637 -746
rect 57671 -774 57699 -746
rect 65759 56147 65787 56175
rect 65821 56147 65849 56175
rect 65759 56085 65787 56113
rect 65821 56085 65849 56113
rect 65759 56023 65787 56051
rect 65821 56023 65849 56051
rect 65759 55961 65787 55989
rect 65821 55961 65849 55989
rect 64625 47147 64653 47175
rect 64687 47147 64715 47175
rect 64749 47147 64777 47175
rect 64811 47147 64839 47175
rect 64625 47085 64653 47113
rect 64687 47085 64715 47113
rect 64749 47085 64777 47113
rect 64811 47085 64839 47113
rect 64625 47023 64653 47051
rect 64687 47023 64715 47051
rect 64749 47023 64777 47051
rect 64811 47023 64839 47051
rect 64625 46961 64653 46989
rect 64687 46961 64715 46989
rect 64749 46961 64777 46989
rect 64811 46961 64839 46989
rect 64625 38147 64653 38175
rect 64687 38147 64715 38175
rect 64749 38147 64777 38175
rect 64811 38147 64839 38175
rect 64625 38085 64653 38113
rect 64687 38085 64715 38113
rect 64749 38085 64777 38113
rect 64811 38085 64839 38113
rect 64625 38023 64653 38051
rect 64687 38023 64715 38051
rect 64749 38023 64777 38051
rect 64811 38023 64839 38051
rect 64625 37961 64653 37989
rect 64687 37961 64715 37989
rect 64749 37961 64777 37989
rect 64811 37961 64839 37989
rect 64625 29147 64653 29175
rect 64687 29147 64715 29175
rect 64749 29147 64777 29175
rect 64811 29147 64839 29175
rect 64625 29085 64653 29113
rect 64687 29085 64715 29113
rect 64749 29085 64777 29113
rect 64811 29085 64839 29113
rect 64625 29023 64653 29051
rect 64687 29023 64715 29051
rect 64749 29023 64777 29051
rect 64811 29023 64839 29051
rect 64625 28961 64653 28989
rect 64687 28961 64715 28989
rect 64749 28961 64777 28989
rect 64811 28961 64839 28989
rect 64625 20147 64653 20175
rect 64687 20147 64715 20175
rect 64749 20147 64777 20175
rect 64811 20147 64839 20175
rect 64625 20085 64653 20113
rect 64687 20085 64715 20113
rect 64749 20085 64777 20113
rect 64811 20085 64839 20113
rect 64625 20023 64653 20051
rect 64687 20023 64715 20051
rect 64749 20023 64777 20051
rect 64811 20023 64839 20051
rect 64625 19961 64653 19989
rect 64687 19961 64715 19989
rect 64749 19961 64777 19989
rect 64811 19961 64839 19989
rect 64625 11147 64653 11175
rect 64687 11147 64715 11175
rect 64749 11147 64777 11175
rect 64811 11147 64839 11175
rect 64625 11085 64653 11113
rect 64687 11085 64715 11113
rect 64749 11085 64777 11113
rect 64811 11085 64839 11113
rect 64625 11023 64653 11051
rect 64687 11023 64715 11051
rect 64749 11023 64777 11051
rect 64811 11023 64839 11051
rect 64625 10961 64653 10989
rect 64687 10961 64715 10989
rect 64749 10961 64777 10989
rect 64811 10961 64839 10989
rect 64625 2147 64653 2175
rect 64687 2147 64715 2175
rect 64749 2147 64777 2175
rect 64811 2147 64839 2175
rect 64625 2085 64653 2113
rect 64687 2085 64715 2113
rect 64749 2085 64777 2113
rect 64811 2085 64839 2113
rect 64625 2023 64653 2051
rect 64687 2023 64715 2051
rect 64749 2023 64777 2051
rect 64811 2023 64839 2051
rect 64625 1961 64653 1989
rect 64687 1961 64715 1989
rect 64749 1961 64777 1989
rect 64811 1961 64839 1989
rect 64625 -108 64653 -80
rect 64687 -108 64715 -80
rect 64749 -108 64777 -80
rect 64811 -108 64839 -80
rect 64625 -170 64653 -142
rect 64687 -170 64715 -142
rect 64749 -170 64777 -142
rect 64811 -170 64839 -142
rect 64625 -232 64653 -204
rect 64687 -232 64715 -204
rect 64749 -232 64777 -204
rect 64811 -232 64839 -204
rect 64625 -294 64653 -266
rect 64687 -294 64715 -266
rect 64749 -294 64777 -266
rect 64811 -294 64839 -266
rect 68009 59147 68037 59175
rect 68071 59147 68099 59175
rect 68009 59085 68037 59113
rect 68071 59085 68099 59113
rect 68009 59023 68037 59051
rect 68071 59023 68099 59051
rect 68009 58961 68037 58989
rect 68071 58961 68099 58989
rect 72509 59147 72537 59175
rect 72571 59147 72599 59175
rect 72509 59085 72537 59113
rect 72571 59085 72599 59113
rect 72509 59023 72537 59051
rect 72571 59023 72599 59051
rect 72509 58961 72537 58989
rect 72571 58961 72599 58989
rect 70259 56147 70287 56175
rect 70321 56147 70349 56175
rect 70259 56085 70287 56113
rect 70321 56085 70349 56113
rect 70259 56023 70287 56051
rect 70321 56023 70349 56051
rect 70259 55961 70287 55989
rect 70321 55961 70349 55989
rect 74759 65147 74787 65175
rect 74821 65147 74849 65175
rect 74759 65085 74787 65113
rect 74821 65085 74849 65113
rect 74759 65023 74787 65051
rect 74821 65023 74849 65051
rect 74759 64961 74787 64989
rect 74821 64961 74849 64989
rect 77009 68147 77037 68175
rect 77071 68147 77099 68175
rect 77009 68085 77037 68113
rect 77071 68085 77099 68113
rect 77009 68023 77037 68051
rect 77071 68023 77099 68051
rect 77009 67961 77037 67989
rect 77071 67961 77099 67989
rect 81509 68147 81537 68175
rect 81571 68147 81599 68175
rect 81509 68085 81537 68113
rect 81571 68085 81599 68113
rect 81509 68023 81537 68051
rect 81571 68023 81599 68051
rect 81509 67961 81537 67989
rect 81571 67961 81599 67989
rect 79259 65147 79287 65175
rect 79321 65147 79349 65175
rect 79259 65085 79287 65113
rect 79321 65085 79349 65113
rect 79259 65023 79287 65051
rect 79321 65023 79349 65051
rect 79259 64961 79287 64989
rect 79321 64961 79349 64989
rect 83759 74147 83787 74175
rect 83821 74147 83849 74175
rect 83759 74085 83787 74113
rect 83821 74085 83849 74113
rect 83759 74023 83787 74051
rect 83821 74023 83849 74051
rect 83759 73961 83787 73989
rect 83821 73961 83849 73989
rect 86009 77147 86037 77175
rect 86071 77147 86099 77175
rect 86009 77085 86037 77113
rect 86071 77085 86099 77113
rect 86009 77023 86037 77051
rect 86071 77023 86099 77051
rect 86009 76961 86037 76989
rect 86071 76961 86099 76989
rect 90509 77147 90537 77175
rect 90571 77147 90599 77175
rect 90509 77085 90537 77113
rect 90571 77085 90599 77113
rect 90509 77023 90537 77051
rect 90571 77023 90599 77051
rect 90509 76961 90537 76989
rect 90571 76961 90599 76989
rect 88259 74147 88287 74175
rect 88321 74147 88349 74175
rect 88259 74085 88287 74113
rect 88321 74085 88349 74113
rect 88259 74023 88287 74051
rect 88321 74023 88349 74051
rect 88259 73961 88287 73989
rect 88321 73961 88349 73989
rect 92759 83147 92787 83175
rect 92821 83147 92849 83175
rect 92759 83085 92787 83113
rect 92821 83085 92849 83113
rect 92759 83023 92787 83051
rect 92821 83023 92849 83051
rect 92759 82961 92787 82989
rect 92821 82961 92849 82989
rect 97259 83147 97287 83175
rect 97321 83147 97349 83175
rect 97259 83085 97287 83113
rect 97321 83085 97349 83113
rect 97259 83023 97287 83051
rect 97321 83023 97349 83051
rect 97259 82961 97287 82989
rect 97321 82961 97349 82989
rect 101759 83147 101787 83175
rect 101821 83147 101849 83175
rect 101759 83085 101787 83113
rect 101821 83085 101849 83113
rect 101759 83023 101787 83051
rect 101821 83023 101849 83051
rect 101759 82961 101787 82989
rect 101821 82961 101849 82989
rect 106259 83147 106287 83175
rect 106321 83147 106349 83175
rect 106259 83085 106287 83113
rect 106321 83085 106349 83113
rect 106259 83023 106287 83051
rect 106321 83023 106349 83051
rect 106259 82961 106287 82989
rect 106321 82961 106349 82989
rect 110759 83147 110787 83175
rect 110821 83147 110849 83175
rect 110759 83085 110787 83113
rect 110821 83085 110849 83113
rect 110759 83023 110787 83051
rect 110821 83023 110849 83051
rect 110759 82961 110787 82989
rect 110821 82961 110849 82989
rect 115259 83147 115287 83175
rect 115321 83147 115349 83175
rect 115259 83085 115287 83113
rect 115321 83085 115349 83113
rect 115259 83023 115287 83051
rect 115321 83023 115349 83051
rect 115259 82961 115287 82989
rect 115321 82961 115349 82989
rect 95009 77147 95037 77175
rect 95071 77147 95099 77175
rect 95009 77085 95037 77113
rect 95071 77085 95099 77113
rect 95009 77023 95037 77051
rect 95071 77023 95099 77051
rect 95009 76961 95037 76989
rect 95071 76961 95099 76989
rect 99509 77147 99537 77175
rect 99571 77147 99599 77175
rect 99509 77085 99537 77113
rect 99571 77085 99599 77113
rect 99509 77023 99537 77051
rect 99571 77023 99599 77051
rect 99509 76961 99537 76989
rect 99571 76961 99599 76989
rect 104009 77147 104037 77175
rect 104071 77147 104099 77175
rect 104009 77085 104037 77113
rect 104071 77085 104099 77113
rect 104009 77023 104037 77051
rect 104071 77023 104099 77051
rect 104009 76961 104037 76989
rect 104071 76961 104099 76989
rect 108509 77147 108537 77175
rect 108571 77147 108599 77175
rect 108509 77085 108537 77113
rect 108571 77085 108599 77113
rect 108509 77023 108537 77051
rect 108571 77023 108599 77051
rect 108509 76961 108537 76989
rect 108571 76961 108599 76989
rect 113009 77147 113037 77175
rect 113071 77147 113099 77175
rect 113009 77085 113037 77113
rect 113071 77085 113099 77113
rect 113009 77023 113037 77051
rect 113071 77023 113099 77051
rect 113009 76961 113037 76989
rect 113071 76961 113099 76989
rect 117509 77147 117537 77175
rect 117571 77147 117599 77175
rect 117509 77085 117537 77113
rect 117571 77085 117599 77113
rect 117509 77023 117537 77051
rect 117571 77023 117599 77051
rect 117509 76961 117537 76989
rect 117571 76961 117599 76989
rect 120485 77147 120513 77175
rect 120547 77147 120575 77175
rect 120609 77147 120637 77175
rect 120671 77147 120699 77175
rect 120485 77085 120513 77113
rect 120547 77085 120575 77113
rect 120609 77085 120637 77113
rect 120671 77085 120699 77113
rect 120485 77023 120513 77051
rect 120547 77023 120575 77051
rect 120609 77023 120637 77051
rect 120671 77023 120699 77051
rect 120485 76961 120513 76989
rect 120547 76961 120575 76989
rect 120609 76961 120637 76989
rect 120671 76961 120699 76989
rect 91625 74147 91653 74175
rect 91687 74147 91715 74175
rect 91749 74147 91777 74175
rect 91811 74147 91839 74175
rect 91625 74085 91653 74113
rect 91687 74085 91715 74113
rect 91749 74085 91777 74113
rect 91811 74085 91839 74113
rect 91625 74023 91653 74051
rect 91687 74023 91715 74051
rect 91749 74023 91777 74051
rect 91811 74023 91839 74051
rect 91625 73961 91653 73989
rect 91687 73961 91715 73989
rect 91749 73961 91777 73989
rect 91811 73961 91839 73989
rect 84485 68147 84513 68175
rect 84547 68147 84575 68175
rect 84609 68147 84637 68175
rect 84671 68147 84699 68175
rect 84485 68085 84513 68113
rect 84547 68085 84575 68113
rect 84609 68085 84637 68113
rect 84671 68085 84699 68113
rect 84485 68023 84513 68051
rect 84547 68023 84575 68051
rect 84609 68023 84637 68051
rect 84671 68023 84699 68051
rect 84485 67961 84513 67989
rect 84547 67961 84575 67989
rect 84609 67961 84637 67989
rect 84671 67961 84699 67989
rect 82625 65147 82653 65175
rect 82687 65147 82715 65175
rect 82749 65147 82777 65175
rect 82811 65147 82839 65175
rect 82625 65085 82653 65113
rect 82687 65085 82715 65113
rect 82749 65085 82777 65113
rect 82811 65085 82839 65113
rect 82625 65023 82653 65051
rect 82687 65023 82715 65051
rect 82749 65023 82777 65051
rect 82811 65023 82839 65051
rect 82625 64961 82653 64989
rect 82687 64961 82715 64989
rect 82749 64961 82777 64989
rect 82811 64961 82839 64989
rect 75485 59147 75513 59175
rect 75547 59147 75575 59175
rect 75609 59147 75637 59175
rect 75671 59147 75699 59175
rect 75485 59085 75513 59113
rect 75547 59085 75575 59113
rect 75609 59085 75637 59113
rect 75671 59085 75699 59113
rect 75485 59023 75513 59051
rect 75547 59023 75575 59051
rect 75609 59023 75637 59051
rect 75671 59023 75699 59051
rect 75485 58961 75513 58989
rect 75547 58961 75575 58989
rect 75609 58961 75637 58989
rect 75671 58961 75699 58989
rect 73625 56147 73653 56175
rect 73687 56147 73715 56175
rect 73749 56147 73777 56175
rect 73811 56147 73839 56175
rect 73625 56085 73653 56113
rect 73687 56085 73715 56113
rect 73749 56085 73777 56113
rect 73811 56085 73839 56113
rect 73625 56023 73653 56051
rect 73687 56023 73715 56051
rect 73749 56023 73777 56051
rect 73811 56023 73839 56051
rect 73625 55961 73653 55989
rect 73687 55961 73715 55989
rect 73749 55961 73777 55989
rect 73811 55961 73839 55989
rect 66485 50147 66513 50175
rect 66547 50147 66575 50175
rect 66609 50147 66637 50175
rect 66671 50147 66699 50175
rect 66485 50085 66513 50113
rect 66547 50085 66575 50113
rect 66609 50085 66637 50113
rect 66671 50085 66699 50113
rect 66485 50023 66513 50051
rect 66547 50023 66575 50051
rect 66609 50023 66637 50051
rect 66671 50023 66699 50051
rect 66485 49961 66513 49989
rect 66547 49961 66575 49989
rect 66609 49961 66637 49989
rect 66671 49961 66699 49989
rect 66485 41147 66513 41175
rect 66547 41147 66575 41175
rect 66609 41147 66637 41175
rect 66671 41147 66699 41175
rect 66485 41085 66513 41113
rect 66547 41085 66575 41113
rect 66609 41085 66637 41113
rect 66671 41085 66699 41113
rect 66485 41023 66513 41051
rect 66547 41023 66575 41051
rect 66609 41023 66637 41051
rect 66671 41023 66699 41051
rect 66485 40961 66513 40989
rect 66547 40961 66575 40989
rect 66609 40961 66637 40989
rect 66671 40961 66699 40989
rect 66485 32147 66513 32175
rect 66547 32147 66575 32175
rect 66609 32147 66637 32175
rect 66671 32147 66699 32175
rect 66485 32085 66513 32113
rect 66547 32085 66575 32113
rect 66609 32085 66637 32113
rect 66671 32085 66699 32113
rect 66485 32023 66513 32051
rect 66547 32023 66575 32051
rect 66609 32023 66637 32051
rect 66671 32023 66699 32051
rect 66485 31961 66513 31989
rect 66547 31961 66575 31989
rect 66609 31961 66637 31989
rect 66671 31961 66699 31989
rect 66485 23147 66513 23175
rect 66547 23147 66575 23175
rect 66609 23147 66637 23175
rect 66671 23147 66699 23175
rect 66485 23085 66513 23113
rect 66547 23085 66575 23113
rect 66609 23085 66637 23113
rect 66671 23085 66699 23113
rect 66485 23023 66513 23051
rect 66547 23023 66575 23051
rect 66609 23023 66637 23051
rect 66671 23023 66699 23051
rect 66485 22961 66513 22989
rect 66547 22961 66575 22989
rect 66609 22961 66637 22989
rect 66671 22961 66699 22989
rect 66485 14147 66513 14175
rect 66547 14147 66575 14175
rect 66609 14147 66637 14175
rect 66671 14147 66699 14175
rect 66485 14085 66513 14113
rect 66547 14085 66575 14113
rect 66609 14085 66637 14113
rect 66671 14085 66699 14113
rect 66485 14023 66513 14051
rect 66547 14023 66575 14051
rect 66609 14023 66637 14051
rect 66671 14023 66699 14051
rect 66485 13961 66513 13989
rect 66547 13961 66575 13989
rect 66609 13961 66637 13989
rect 66671 13961 66699 13989
rect 66485 5147 66513 5175
rect 66547 5147 66575 5175
rect 66609 5147 66637 5175
rect 66671 5147 66699 5175
rect 66485 5085 66513 5113
rect 66547 5085 66575 5113
rect 66609 5085 66637 5113
rect 66671 5085 66699 5113
rect 66485 5023 66513 5051
rect 66547 5023 66575 5051
rect 66609 5023 66637 5051
rect 66671 5023 66699 5051
rect 66485 4961 66513 4989
rect 66547 4961 66575 4989
rect 66609 4961 66637 4989
rect 66671 4961 66699 4989
rect 66485 -588 66513 -560
rect 66547 -588 66575 -560
rect 66609 -588 66637 -560
rect 66671 -588 66699 -560
rect 66485 -650 66513 -622
rect 66547 -650 66575 -622
rect 66609 -650 66637 -622
rect 66671 -650 66699 -622
rect 66485 -712 66513 -684
rect 66547 -712 66575 -684
rect 66609 -712 66637 -684
rect 66671 -712 66699 -684
rect 66485 -774 66513 -746
rect 66547 -774 66575 -746
rect 66609 -774 66637 -746
rect 66671 -774 66699 -746
rect 74759 56147 74787 56175
rect 74821 56147 74849 56175
rect 74759 56085 74787 56113
rect 74821 56085 74849 56113
rect 74759 56023 74787 56051
rect 74821 56023 74849 56051
rect 74759 55961 74787 55989
rect 74821 55961 74849 55989
rect 73625 47147 73653 47175
rect 73687 47147 73715 47175
rect 73749 47147 73777 47175
rect 73811 47147 73839 47175
rect 73625 47085 73653 47113
rect 73687 47085 73715 47113
rect 73749 47085 73777 47113
rect 73811 47085 73839 47113
rect 73625 47023 73653 47051
rect 73687 47023 73715 47051
rect 73749 47023 73777 47051
rect 73811 47023 73839 47051
rect 73625 46961 73653 46989
rect 73687 46961 73715 46989
rect 73749 46961 73777 46989
rect 73811 46961 73839 46989
rect 73625 38147 73653 38175
rect 73687 38147 73715 38175
rect 73749 38147 73777 38175
rect 73811 38147 73839 38175
rect 73625 38085 73653 38113
rect 73687 38085 73715 38113
rect 73749 38085 73777 38113
rect 73811 38085 73839 38113
rect 73625 38023 73653 38051
rect 73687 38023 73715 38051
rect 73749 38023 73777 38051
rect 73811 38023 73839 38051
rect 73625 37961 73653 37989
rect 73687 37961 73715 37989
rect 73749 37961 73777 37989
rect 73811 37961 73839 37989
rect 73625 29147 73653 29175
rect 73687 29147 73715 29175
rect 73749 29147 73777 29175
rect 73811 29147 73839 29175
rect 73625 29085 73653 29113
rect 73687 29085 73715 29113
rect 73749 29085 73777 29113
rect 73811 29085 73839 29113
rect 73625 29023 73653 29051
rect 73687 29023 73715 29051
rect 73749 29023 73777 29051
rect 73811 29023 73839 29051
rect 73625 28961 73653 28989
rect 73687 28961 73715 28989
rect 73749 28961 73777 28989
rect 73811 28961 73839 28989
rect 73625 20147 73653 20175
rect 73687 20147 73715 20175
rect 73749 20147 73777 20175
rect 73811 20147 73839 20175
rect 73625 20085 73653 20113
rect 73687 20085 73715 20113
rect 73749 20085 73777 20113
rect 73811 20085 73839 20113
rect 73625 20023 73653 20051
rect 73687 20023 73715 20051
rect 73749 20023 73777 20051
rect 73811 20023 73839 20051
rect 73625 19961 73653 19989
rect 73687 19961 73715 19989
rect 73749 19961 73777 19989
rect 73811 19961 73839 19989
rect 73625 11147 73653 11175
rect 73687 11147 73715 11175
rect 73749 11147 73777 11175
rect 73811 11147 73839 11175
rect 73625 11085 73653 11113
rect 73687 11085 73715 11113
rect 73749 11085 73777 11113
rect 73811 11085 73839 11113
rect 73625 11023 73653 11051
rect 73687 11023 73715 11051
rect 73749 11023 73777 11051
rect 73811 11023 73839 11051
rect 73625 10961 73653 10989
rect 73687 10961 73715 10989
rect 73749 10961 73777 10989
rect 73811 10961 73839 10989
rect 73625 2147 73653 2175
rect 73687 2147 73715 2175
rect 73749 2147 73777 2175
rect 73811 2147 73839 2175
rect 73625 2085 73653 2113
rect 73687 2085 73715 2113
rect 73749 2085 73777 2113
rect 73811 2085 73839 2113
rect 73625 2023 73653 2051
rect 73687 2023 73715 2051
rect 73749 2023 73777 2051
rect 73811 2023 73839 2051
rect 73625 1961 73653 1989
rect 73687 1961 73715 1989
rect 73749 1961 73777 1989
rect 73811 1961 73839 1989
rect 73625 -108 73653 -80
rect 73687 -108 73715 -80
rect 73749 -108 73777 -80
rect 73811 -108 73839 -80
rect 73625 -170 73653 -142
rect 73687 -170 73715 -142
rect 73749 -170 73777 -142
rect 73811 -170 73839 -142
rect 73625 -232 73653 -204
rect 73687 -232 73715 -204
rect 73749 -232 73777 -204
rect 73811 -232 73839 -204
rect 73625 -294 73653 -266
rect 73687 -294 73715 -266
rect 73749 -294 73777 -266
rect 73811 -294 73839 -266
rect 77009 59147 77037 59175
rect 77071 59147 77099 59175
rect 77009 59085 77037 59113
rect 77071 59085 77099 59113
rect 77009 59023 77037 59051
rect 77071 59023 77099 59051
rect 77009 58961 77037 58989
rect 77071 58961 77099 58989
rect 81509 59147 81537 59175
rect 81571 59147 81599 59175
rect 81509 59085 81537 59113
rect 81571 59085 81599 59113
rect 81509 59023 81537 59051
rect 81571 59023 81599 59051
rect 81509 58961 81537 58989
rect 81571 58961 81599 58989
rect 79259 56147 79287 56175
rect 79321 56147 79349 56175
rect 79259 56085 79287 56113
rect 79321 56085 79349 56113
rect 79259 56023 79287 56051
rect 79321 56023 79349 56051
rect 79259 55961 79287 55989
rect 79321 55961 79349 55989
rect 83759 65147 83787 65175
rect 83821 65147 83849 65175
rect 83759 65085 83787 65113
rect 83821 65085 83849 65113
rect 83759 65023 83787 65051
rect 83821 65023 83849 65051
rect 83759 64961 83787 64989
rect 83821 64961 83849 64989
rect 86009 68147 86037 68175
rect 86071 68147 86099 68175
rect 86009 68085 86037 68113
rect 86071 68085 86099 68113
rect 86009 68023 86037 68051
rect 86071 68023 86099 68051
rect 86009 67961 86037 67989
rect 86071 67961 86099 67989
rect 90509 68147 90537 68175
rect 90571 68147 90599 68175
rect 90509 68085 90537 68113
rect 90571 68085 90599 68113
rect 90509 68023 90537 68051
rect 90571 68023 90599 68051
rect 90509 67961 90537 67989
rect 90571 67961 90599 67989
rect 88259 65147 88287 65175
rect 88321 65147 88349 65175
rect 88259 65085 88287 65113
rect 88321 65085 88349 65113
rect 88259 65023 88287 65051
rect 88321 65023 88349 65051
rect 88259 64961 88287 64989
rect 88321 64961 88349 64989
rect 92759 74147 92787 74175
rect 92821 74147 92849 74175
rect 92759 74085 92787 74113
rect 92821 74085 92849 74113
rect 92759 74023 92787 74051
rect 92821 74023 92849 74051
rect 92759 73961 92787 73989
rect 92821 73961 92849 73989
rect 97259 74147 97287 74175
rect 97321 74147 97349 74175
rect 97259 74085 97287 74113
rect 97321 74085 97349 74113
rect 97259 74023 97287 74051
rect 97321 74023 97349 74051
rect 97259 73961 97287 73989
rect 97321 73961 97349 73989
rect 101759 74147 101787 74175
rect 101821 74147 101849 74175
rect 101759 74085 101787 74113
rect 101821 74085 101849 74113
rect 101759 74023 101787 74051
rect 101821 74023 101849 74051
rect 101759 73961 101787 73989
rect 101821 73961 101849 73989
rect 106259 74147 106287 74175
rect 106321 74147 106349 74175
rect 106259 74085 106287 74113
rect 106321 74085 106349 74113
rect 106259 74023 106287 74051
rect 106321 74023 106349 74051
rect 106259 73961 106287 73989
rect 106321 73961 106349 73989
rect 110759 74147 110787 74175
rect 110821 74147 110849 74175
rect 110759 74085 110787 74113
rect 110821 74085 110849 74113
rect 110759 74023 110787 74051
rect 110821 74023 110849 74051
rect 110759 73961 110787 73989
rect 110821 73961 110849 73989
rect 115259 74147 115287 74175
rect 115321 74147 115349 74175
rect 115259 74085 115287 74113
rect 115321 74085 115349 74113
rect 115259 74023 115287 74051
rect 115321 74023 115349 74051
rect 115259 73961 115287 73989
rect 115321 73961 115349 73989
rect 95009 68147 95037 68175
rect 95071 68147 95099 68175
rect 95009 68085 95037 68113
rect 95071 68085 95099 68113
rect 95009 68023 95037 68051
rect 95071 68023 95099 68051
rect 95009 67961 95037 67989
rect 95071 67961 95099 67989
rect 99509 68147 99537 68175
rect 99571 68147 99599 68175
rect 99509 68085 99537 68113
rect 99571 68085 99599 68113
rect 99509 68023 99537 68051
rect 99571 68023 99599 68051
rect 99509 67961 99537 67989
rect 99571 67961 99599 67989
rect 104009 68147 104037 68175
rect 104071 68147 104099 68175
rect 104009 68085 104037 68113
rect 104071 68085 104099 68113
rect 104009 68023 104037 68051
rect 104071 68023 104099 68051
rect 104009 67961 104037 67989
rect 104071 67961 104099 67989
rect 108509 68147 108537 68175
rect 108571 68147 108599 68175
rect 108509 68085 108537 68113
rect 108571 68085 108599 68113
rect 108509 68023 108537 68051
rect 108571 68023 108599 68051
rect 108509 67961 108537 67989
rect 108571 67961 108599 67989
rect 113009 68147 113037 68175
rect 113071 68147 113099 68175
rect 113009 68085 113037 68113
rect 113071 68085 113099 68113
rect 113009 68023 113037 68051
rect 113071 68023 113099 68051
rect 113009 67961 113037 67989
rect 113071 67961 113099 67989
rect 117509 68147 117537 68175
rect 117571 68147 117599 68175
rect 117509 68085 117537 68113
rect 117571 68085 117599 68113
rect 117509 68023 117537 68051
rect 117571 68023 117599 68051
rect 117509 67961 117537 67989
rect 117571 67961 117599 67989
rect 120485 68147 120513 68175
rect 120547 68147 120575 68175
rect 120609 68147 120637 68175
rect 120671 68147 120699 68175
rect 120485 68085 120513 68113
rect 120547 68085 120575 68113
rect 120609 68085 120637 68113
rect 120671 68085 120699 68113
rect 120485 68023 120513 68051
rect 120547 68023 120575 68051
rect 120609 68023 120637 68051
rect 120671 68023 120699 68051
rect 120485 67961 120513 67989
rect 120547 67961 120575 67989
rect 120609 67961 120637 67989
rect 120671 67961 120699 67989
rect 91625 65147 91653 65175
rect 91687 65147 91715 65175
rect 91749 65147 91777 65175
rect 91811 65147 91839 65175
rect 91625 65085 91653 65113
rect 91687 65085 91715 65113
rect 91749 65085 91777 65113
rect 91811 65085 91839 65113
rect 91625 65023 91653 65051
rect 91687 65023 91715 65051
rect 91749 65023 91777 65051
rect 91811 65023 91839 65051
rect 91625 64961 91653 64989
rect 91687 64961 91715 64989
rect 91749 64961 91777 64989
rect 91811 64961 91839 64989
rect 84485 59147 84513 59175
rect 84547 59147 84575 59175
rect 84609 59147 84637 59175
rect 84671 59147 84699 59175
rect 84485 59085 84513 59113
rect 84547 59085 84575 59113
rect 84609 59085 84637 59113
rect 84671 59085 84699 59113
rect 84485 59023 84513 59051
rect 84547 59023 84575 59051
rect 84609 59023 84637 59051
rect 84671 59023 84699 59051
rect 84485 58961 84513 58989
rect 84547 58961 84575 58989
rect 84609 58961 84637 58989
rect 84671 58961 84699 58989
rect 82625 56147 82653 56175
rect 82687 56147 82715 56175
rect 82749 56147 82777 56175
rect 82811 56147 82839 56175
rect 82625 56085 82653 56113
rect 82687 56085 82715 56113
rect 82749 56085 82777 56113
rect 82811 56085 82839 56113
rect 82625 56023 82653 56051
rect 82687 56023 82715 56051
rect 82749 56023 82777 56051
rect 82811 56023 82839 56051
rect 82625 55961 82653 55989
rect 82687 55961 82715 55989
rect 82749 55961 82777 55989
rect 82811 55961 82839 55989
rect 75485 50147 75513 50175
rect 75547 50147 75575 50175
rect 75609 50147 75637 50175
rect 75671 50147 75699 50175
rect 75485 50085 75513 50113
rect 75547 50085 75575 50113
rect 75609 50085 75637 50113
rect 75671 50085 75699 50113
rect 75485 50023 75513 50051
rect 75547 50023 75575 50051
rect 75609 50023 75637 50051
rect 75671 50023 75699 50051
rect 75485 49961 75513 49989
rect 75547 49961 75575 49989
rect 75609 49961 75637 49989
rect 75671 49961 75699 49989
rect 75485 41147 75513 41175
rect 75547 41147 75575 41175
rect 75609 41147 75637 41175
rect 75671 41147 75699 41175
rect 75485 41085 75513 41113
rect 75547 41085 75575 41113
rect 75609 41085 75637 41113
rect 75671 41085 75699 41113
rect 75485 41023 75513 41051
rect 75547 41023 75575 41051
rect 75609 41023 75637 41051
rect 75671 41023 75699 41051
rect 75485 40961 75513 40989
rect 75547 40961 75575 40989
rect 75609 40961 75637 40989
rect 75671 40961 75699 40989
rect 75485 32147 75513 32175
rect 75547 32147 75575 32175
rect 75609 32147 75637 32175
rect 75671 32147 75699 32175
rect 75485 32085 75513 32113
rect 75547 32085 75575 32113
rect 75609 32085 75637 32113
rect 75671 32085 75699 32113
rect 75485 32023 75513 32051
rect 75547 32023 75575 32051
rect 75609 32023 75637 32051
rect 75671 32023 75699 32051
rect 75485 31961 75513 31989
rect 75547 31961 75575 31989
rect 75609 31961 75637 31989
rect 75671 31961 75699 31989
rect 75485 23147 75513 23175
rect 75547 23147 75575 23175
rect 75609 23147 75637 23175
rect 75671 23147 75699 23175
rect 75485 23085 75513 23113
rect 75547 23085 75575 23113
rect 75609 23085 75637 23113
rect 75671 23085 75699 23113
rect 75485 23023 75513 23051
rect 75547 23023 75575 23051
rect 75609 23023 75637 23051
rect 75671 23023 75699 23051
rect 75485 22961 75513 22989
rect 75547 22961 75575 22989
rect 75609 22961 75637 22989
rect 75671 22961 75699 22989
rect 75485 14147 75513 14175
rect 75547 14147 75575 14175
rect 75609 14147 75637 14175
rect 75671 14147 75699 14175
rect 75485 14085 75513 14113
rect 75547 14085 75575 14113
rect 75609 14085 75637 14113
rect 75671 14085 75699 14113
rect 75485 14023 75513 14051
rect 75547 14023 75575 14051
rect 75609 14023 75637 14051
rect 75671 14023 75699 14051
rect 75485 13961 75513 13989
rect 75547 13961 75575 13989
rect 75609 13961 75637 13989
rect 75671 13961 75699 13989
rect 75485 5147 75513 5175
rect 75547 5147 75575 5175
rect 75609 5147 75637 5175
rect 75671 5147 75699 5175
rect 75485 5085 75513 5113
rect 75547 5085 75575 5113
rect 75609 5085 75637 5113
rect 75671 5085 75699 5113
rect 75485 5023 75513 5051
rect 75547 5023 75575 5051
rect 75609 5023 75637 5051
rect 75671 5023 75699 5051
rect 75485 4961 75513 4989
rect 75547 4961 75575 4989
rect 75609 4961 75637 4989
rect 75671 4961 75699 4989
rect 75485 -588 75513 -560
rect 75547 -588 75575 -560
rect 75609 -588 75637 -560
rect 75671 -588 75699 -560
rect 75485 -650 75513 -622
rect 75547 -650 75575 -622
rect 75609 -650 75637 -622
rect 75671 -650 75699 -622
rect 75485 -712 75513 -684
rect 75547 -712 75575 -684
rect 75609 -712 75637 -684
rect 75671 -712 75699 -684
rect 75485 -774 75513 -746
rect 75547 -774 75575 -746
rect 75609 -774 75637 -746
rect 75671 -774 75699 -746
rect 83759 56147 83787 56175
rect 83821 56147 83849 56175
rect 83759 56085 83787 56113
rect 83821 56085 83849 56113
rect 83759 56023 83787 56051
rect 83821 56023 83849 56051
rect 83759 55961 83787 55989
rect 83821 55961 83849 55989
rect 82625 47147 82653 47175
rect 82687 47147 82715 47175
rect 82749 47147 82777 47175
rect 82811 47147 82839 47175
rect 82625 47085 82653 47113
rect 82687 47085 82715 47113
rect 82749 47085 82777 47113
rect 82811 47085 82839 47113
rect 82625 47023 82653 47051
rect 82687 47023 82715 47051
rect 82749 47023 82777 47051
rect 82811 47023 82839 47051
rect 82625 46961 82653 46989
rect 82687 46961 82715 46989
rect 82749 46961 82777 46989
rect 82811 46961 82839 46989
rect 82625 38147 82653 38175
rect 82687 38147 82715 38175
rect 82749 38147 82777 38175
rect 82811 38147 82839 38175
rect 82625 38085 82653 38113
rect 82687 38085 82715 38113
rect 82749 38085 82777 38113
rect 82811 38085 82839 38113
rect 82625 38023 82653 38051
rect 82687 38023 82715 38051
rect 82749 38023 82777 38051
rect 82811 38023 82839 38051
rect 82625 37961 82653 37989
rect 82687 37961 82715 37989
rect 82749 37961 82777 37989
rect 82811 37961 82839 37989
rect 82625 29147 82653 29175
rect 82687 29147 82715 29175
rect 82749 29147 82777 29175
rect 82811 29147 82839 29175
rect 82625 29085 82653 29113
rect 82687 29085 82715 29113
rect 82749 29085 82777 29113
rect 82811 29085 82839 29113
rect 82625 29023 82653 29051
rect 82687 29023 82715 29051
rect 82749 29023 82777 29051
rect 82811 29023 82839 29051
rect 82625 28961 82653 28989
rect 82687 28961 82715 28989
rect 82749 28961 82777 28989
rect 82811 28961 82839 28989
rect 82625 20147 82653 20175
rect 82687 20147 82715 20175
rect 82749 20147 82777 20175
rect 82811 20147 82839 20175
rect 82625 20085 82653 20113
rect 82687 20085 82715 20113
rect 82749 20085 82777 20113
rect 82811 20085 82839 20113
rect 82625 20023 82653 20051
rect 82687 20023 82715 20051
rect 82749 20023 82777 20051
rect 82811 20023 82839 20051
rect 82625 19961 82653 19989
rect 82687 19961 82715 19989
rect 82749 19961 82777 19989
rect 82811 19961 82839 19989
rect 82625 11147 82653 11175
rect 82687 11147 82715 11175
rect 82749 11147 82777 11175
rect 82811 11147 82839 11175
rect 82625 11085 82653 11113
rect 82687 11085 82715 11113
rect 82749 11085 82777 11113
rect 82811 11085 82839 11113
rect 82625 11023 82653 11051
rect 82687 11023 82715 11051
rect 82749 11023 82777 11051
rect 82811 11023 82839 11051
rect 82625 10961 82653 10989
rect 82687 10961 82715 10989
rect 82749 10961 82777 10989
rect 82811 10961 82839 10989
rect 82625 2147 82653 2175
rect 82687 2147 82715 2175
rect 82749 2147 82777 2175
rect 82811 2147 82839 2175
rect 82625 2085 82653 2113
rect 82687 2085 82715 2113
rect 82749 2085 82777 2113
rect 82811 2085 82839 2113
rect 82625 2023 82653 2051
rect 82687 2023 82715 2051
rect 82749 2023 82777 2051
rect 82811 2023 82839 2051
rect 82625 1961 82653 1989
rect 82687 1961 82715 1989
rect 82749 1961 82777 1989
rect 82811 1961 82839 1989
rect 82625 -108 82653 -80
rect 82687 -108 82715 -80
rect 82749 -108 82777 -80
rect 82811 -108 82839 -80
rect 82625 -170 82653 -142
rect 82687 -170 82715 -142
rect 82749 -170 82777 -142
rect 82811 -170 82839 -142
rect 82625 -232 82653 -204
rect 82687 -232 82715 -204
rect 82749 -232 82777 -204
rect 82811 -232 82839 -204
rect 82625 -294 82653 -266
rect 82687 -294 82715 -266
rect 82749 -294 82777 -266
rect 82811 -294 82839 -266
rect 86009 59147 86037 59175
rect 86071 59147 86099 59175
rect 86009 59085 86037 59113
rect 86071 59085 86099 59113
rect 86009 59023 86037 59051
rect 86071 59023 86099 59051
rect 86009 58961 86037 58989
rect 86071 58961 86099 58989
rect 90509 59147 90537 59175
rect 90571 59147 90599 59175
rect 90509 59085 90537 59113
rect 90571 59085 90599 59113
rect 90509 59023 90537 59051
rect 90571 59023 90599 59051
rect 90509 58961 90537 58989
rect 90571 58961 90599 58989
rect 88259 56147 88287 56175
rect 88321 56147 88349 56175
rect 88259 56085 88287 56113
rect 88321 56085 88349 56113
rect 88259 56023 88287 56051
rect 88321 56023 88349 56051
rect 88259 55961 88287 55989
rect 88321 55961 88349 55989
rect 92759 65147 92787 65175
rect 92821 65147 92849 65175
rect 92759 65085 92787 65113
rect 92821 65085 92849 65113
rect 92759 65023 92787 65051
rect 92821 65023 92849 65051
rect 92759 64961 92787 64989
rect 92821 64961 92849 64989
rect 97259 65147 97287 65175
rect 97321 65147 97349 65175
rect 97259 65085 97287 65113
rect 97321 65085 97349 65113
rect 97259 65023 97287 65051
rect 97321 65023 97349 65051
rect 97259 64961 97287 64989
rect 97321 64961 97349 64989
rect 101759 65147 101787 65175
rect 101821 65147 101849 65175
rect 101759 65085 101787 65113
rect 101821 65085 101849 65113
rect 101759 65023 101787 65051
rect 101821 65023 101849 65051
rect 101759 64961 101787 64989
rect 101821 64961 101849 64989
rect 106259 65147 106287 65175
rect 106321 65147 106349 65175
rect 106259 65085 106287 65113
rect 106321 65085 106349 65113
rect 106259 65023 106287 65051
rect 106321 65023 106349 65051
rect 106259 64961 106287 64989
rect 106321 64961 106349 64989
rect 110759 65147 110787 65175
rect 110821 65147 110849 65175
rect 110759 65085 110787 65113
rect 110821 65085 110849 65113
rect 110759 65023 110787 65051
rect 110821 65023 110849 65051
rect 110759 64961 110787 64989
rect 110821 64961 110849 64989
rect 115259 65147 115287 65175
rect 115321 65147 115349 65175
rect 115259 65085 115287 65113
rect 115321 65085 115349 65113
rect 115259 65023 115287 65051
rect 115321 65023 115349 65051
rect 115259 64961 115287 64989
rect 115321 64961 115349 64989
rect 95009 59147 95037 59175
rect 95071 59147 95099 59175
rect 95009 59085 95037 59113
rect 95071 59085 95099 59113
rect 95009 59023 95037 59051
rect 95071 59023 95099 59051
rect 95009 58961 95037 58989
rect 95071 58961 95099 58989
rect 99509 59147 99537 59175
rect 99571 59147 99599 59175
rect 99509 59085 99537 59113
rect 99571 59085 99599 59113
rect 99509 59023 99537 59051
rect 99571 59023 99599 59051
rect 99509 58961 99537 58989
rect 99571 58961 99599 58989
rect 104009 59147 104037 59175
rect 104071 59147 104099 59175
rect 104009 59085 104037 59113
rect 104071 59085 104099 59113
rect 104009 59023 104037 59051
rect 104071 59023 104099 59051
rect 104009 58961 104037 58989
rect 104071 58961 104099 58989
rect 108509 59147 108537 59175
rect 108571 59147 108599 59175
rect 108509 59085 108537 59113
rect 108571 59085 108599 59113
rect 108509 59023 108537 59051
rect 108571 59023 108599 59051
rect 108509 58961 108537 58989
rect 108571 58961 108599 58989
rect 113009 59147 113037 59175
rect 113071 59147 113099 59175
rect 113009 59085 113037 59113
rect 113071 59085 113099 59113
rect 113009 59023 113037 59051
rect 113071 59023 113099 59051
rect 113009 58961 113037 58989
rect 113071 58961 113099 58989
rect 117509 59147 117537 59175
rect 117571 59147 117599 59175
rect 117509 59085 117537 59113
rect 117571 59085 117599 59113
rect 117509 59023 117537 59051
rect 117571 59023 117599 59051
rect 117509 58961 117537 58989
rect 117571 58961 117599 58989
rect 120485 59147 120513 59175
rect 120547 59147 120575 59175
rect 120609 59147 120637 59175
rect 120671 59147 120699 59175
rect 120485 59085 120513 59113
rect 120547 59085 120575 59113
rect 120609 59085 120637 59113
rect 120671 59085 120699 59113
rect 120485 59023 120513 59051
rect 120547 59023 120575 59051
rect 120609 59023 120637 59051
rect 120671 59023 120699 59051
rect 120485 58961 120513 58989
rect 120547 58961 120575 58989
rect 120609 58961 120637 58989
rect 120671 58961 120699 58989
rect 91625 56147 91653 56175
rect 91687 56147 91715 56175
rect 91749 56147 91777 56175
rect 91811 56147 91839 56175
rect 91625 56085 91653 56113
rect 91687 56085 91715 56113
rect 91749 56085 91777 56113
rect 91811 56085 91839 56113
rect 91625 56023 91653 56051
rect 91687 56023 91715 56051
rect 91749 56023 91777 56051
rect 91811 56023 91839 56051
rect 91625 55961 91653 55989
rect 91687 55961 91715 55989
rect 91749 55961 91777 55989
rect 91811 55961 91839 55989
rect 84485 50147 84513 50175
rect 84547 50147 84575 50175
rect 84609 50147 84637 50175
rect 84671 50147 84699 50175
rect 84485 50085 84513 50113
rect 84547 50085 84575 50113
rect 84609 50085 84637 50113
rect 84671 50085 84699 50113
rect 84485 50023 84513 50051
rect 84547 50023 84575 50051
rect 84609 50023 84637 50051
rect 84671 50023 84699 50051
rect 84485 49961 84513 49989
rect 84547 49961 84575 49989
rect 84609 49961 84637 49989
rect 84671 49961 84699 49989
rect 84485 41147 84513 41175
rect 84547 41147 84575 41175
rect 84609 41147 84637 41175
rect 84671 41147 84699 41175
rect 84485 41085 84513 41113
rect 84547 41085 84575 41113
rect 84609 41085 84637 41113
rect 84671 41085 84699 41113
rect 84485 41023 84513 41051
rect 84547 41023 84575 41051
rect 84609 41023 84637 41051
rect 84671 41023 84699 41051
rect 84485 40961 84513 40989
rect 84547 40961 84575 40989
rect 84609 40961 84637 40989
rect 84671 40961 84699 40989
rect 84485 32147 84513 32175
rect 84547 32147 84575 32175
rect 84609 32147 84637 32175
rect 84671 32147 84699 32175
rect 84485 32085 84513 32113
rect 84547 32085 84575 32113
rect 84609 32085 84637 32113
rect 84671 32085 84699 32113
rect 84485 32023 84513 32051
rect 84547 32023 84575 32051
rect 84609 32023 84637 32051
rect 84671 32023 84699 32051
rect 84485 31961 84513 31989
rect 84547 31961 84575 31989
rect 84609 31961 84637 31989
rect 84671 31961 84699 31989
rect 84485 23147 84513 23175
rect 84547 23147 84575 23175
rect 84609 23147 84637 23175
rect 84671 23147 84699 23175
rect 84485 23085 84513 23113
rect 84547 23085 84575 23113
rect 84609 23085 84637 23113
rect 84671 23085 84699 23113
rect 84485 23023 84513 23051
rect 84547 23023 84575 23051
rect 84609 23023 84637 23051
rect 84671 23023 84699 23051
rect 84485 22961 84513 22989
rect 84547 22961 84575 22989
rect 84609 22961 84637 22989
rect 84671 22961 84699 22989
rect 84485 14147 84513 14175
rect 84547 14147 84575 14175
rect 84609 14147 84637 14175
rect 84671 14147 84699 14175
rect 84485 14085 84513 14113
rect 84547 14085 84575 14113
rect 84609 14085 84637 14113
rect 84671 14085 84699 14113
rect 84485 14023 84513 14051
rect 84547 14023 84575 14051
rect 84609 14023 84637 14051
rect 84671 14023 84699 14051
rect 84485 13961 84513 13989
rect 84547 13961 84575 13989
rect 84609 13961 84637 13989
rect 84671 13961 84699 13989
rect 84485 5147 84513 5175
rect 84547 5147 84575 5175
rect 84609 5147 84637 5175
rect 84671 5147 84699 5175
rect 84485 5085 84513 5113
rect 84547 5085 84575 5113
rect 84609 5085 84637 5113
rect 84671 5085 84699 5113
rect 84485 5023 84513 5051
rect 84547 5023 84575 5051
rect 84609 5023 84637 5051
rect 84671 5023 84699 5051
rect 84485 4961 84513 4989
rect 84547 4961 84575 4989
rect 84609 4961 84637 4989
rect 84671 4961 84699 4989
rect 84485 -588 84513 -560
rect 84547 -588 84575 -560
rect 84609 -588 84637 -560
rect 84671 -588 84699 -560
rect 84485 -650 84513 -622
rect 84547 -650 84575 -622
rect 84609 -650 84637 -622
rect 84671 -650 84699 -622
rect 84485 -712 84513 -684
rect 84547 -712 84575 -684
rect 84609 -712 84637 -684
rect 84671 -712 84699 -684
rect 84485 -774 84513 -746
rect 84547 -774 84575 -746
rect 84609 -774 84637 -746
rect 84671 -774 84699 -746
rect 92759 56147 92787 56175
rect 92821 56147 92849 56175
rect 92759 56085 92787 56113
rect 92821 56085 92849 56113
rect 92759 56023 92787 56051
rect 92821 56023 92849 56051
rect 92759 55961 92787 55989
rect 92821 55961 92849 55989
rect 97259 56147 97287 56175
rect 97321 56147 97349 56175
rect 97259 56085 97287 56113
rect 97321 56085 97349 56113
rect 97259 56023 97287 56051
rect 97321 56023 97349 56051
rect 97259 55961 97287 55989
rect 97321 55961 97349 55989
rect 101759 56147 101787 56175
rect 101821 56147 101849 56175
rect 101759 56085 101787 56113
rect 101821 56085 101849 56113
rect 101759 56023 101787 56051
rect 101821 56023 101849 56051
rect 101759 55961 101787 55989
rect 101821 55961 101849 55989
rect 106259 56147 106287 56175
rect 106321 56147 106349 56175
rect 106259 56085 106287 56113
rect 106321 56085 106349 56113
rect 106259 56023 106287 56051
rect 106321 56023 106349 56051
rect 106259 55961 106287 55989
rect 106321 55961 106349 55989
rect 110759 56147 110787 56175
rect 110821 56147 110849 56175
rect 110759 56085 110787 56113
rect 110821 56085 110849 56113
rect 110759 56023 110787 56051
rect 110821 56023 110849 56051
rect 110759 55961 110787 55989
rect 110821 55961 110849 55989
rect 115259 56147 115287 56175
rect 115321 56147 115349 56175
rect 115259 56085 115287 56113
rect 115321 56085 115349 56113
rect 115259 56023 115287 56051
rect 115321 56023 115349 56051
rect 115259 55961 115287 55989
rect 115321 55961 115349 55989
rect 120485 50147 120513 50175
rect 120547 50147 120575 50175
rect 120609 50147 120637 50175
rect 120671 50147 120699 50175
rect 120485 50085 120513 50113
rect 120547 50085 120575 50113
rect 120609 50085 120637 50113
rect 120671 50085 120699 50113
rect 120485 50023 120513 50051
rect 120547 50023 120575 50051
rect 120609 50023 120637 50051
rect 120671 50023 120699 50051
rect 120485 49961 120513 49989
rect 120547 49961 120575 49989
rect 120609 49961 120637 49989
rect 120671 49961 120699 49989
rect 91625 47147 91653 47175
rect 91687 47147 91715 47175
rect 91749 47147 91777 47175
rect 91811 47147 91839 47175
rect 91625 47085 91653 47113
rect 91687 47085 91715 47113
rect 91749 47085 91777 47113
rect 91811 47085 91839 47113
rect 91625 47023 91653 47051
rect 91687 47023 91715 47051
rect 91749 47023 91777 47051
rect 91811 47023 91839 47051
rect 91625 46961 91653 46989
rect 91687 46961 91715 46989
rect 91749 46961 91777 46989
rect 91811 46961 91839 46989
rect 91625 38147 91653 38175
rect 91687 38147 91715 38175
rect 91749 38147 91777 38175
rect 91811 38147 91839 38175
rect 91625 38085 91653 38113
rect 91687 38085 91715 38113
rect 91749 38085 91777 38113
rect 91811 38085 91839 38113
rect 91625 38023 91653 38051
rect 91687 38023 91715 38051
rect 91749 38023 91777 38051
rect 91811 38023 91839 38051
rect 91625 37961 91653 37989
rect 91687 37961 91715 37989
rect 91749 37961 91777 37989
rect 91811 37961 91839 37989
rect 91625 29147 91653 29175
rect 91687 29147 91715 29175
rect 91749 29147 91777 29175
rect 91811 29147 91839 29175
rect 91625 29085 91653 29113
rect 91687 29085 91715 29113
rect 91749 29085 91777 29113
rect 91811 29085 91839 29113
rect 91625 29023 91653 29051
rect 91687 29023 91715 29051
rect 91749 29023 91777 29051
rect 91811 29023 91839 29051
rect 91625 28961 91653 28989
rect 91687 28961 91715 28989
rect 91749 28961 91777 28989
rect 91811 28961 91839 28989
rect 91625 20147 91653 20175
rect 91687 20147 91715 20175
rect 91749 20147 91777 20175
rect 91811 20147 91839 20175
rect 91625 20085 91653 20113
rect 91687 20085 91715 20113
rect 91749 20085 91777 20113
rect 91811 20085 91839 20113
rect 91625 20023 91653 20051
rect 91687 20023 91715 20051
rect 91749 20023 91777 20051
rect 91811 20023 91839 20051
rect 91625 19961 91653 19989
rect 91687 19961 91715 19989
rect 91749 19961 91777 19989
rect 91811 19961 91839 19989
rect 91625 11147 91653 11175
rect 91687 11147 91715 11175
rect 91749 11147 91777 11175
rect 91811 11147 91839 11175
rect 91625 11085 91653 11113
rect 91687 11085 91715 11113
rect 91749 11085 91777 11113
rect 91811 11085 91839 11113
rect 91625 11023 91653 11051
rect 91687 11023 91715 11051
rect 91749 11023 91777 11051
rect 91811 11023 91839 11051
rect 91625 10961 91653 10989
rect 91687 10961 91715 10989
rect 91749 10961 91777 10989
rect 91811 10961 91839 10989
rect 91625 2147 91653 2175
rect 91687 2147 91715 2175
rect 91749 2147 91777 2175
rect 91811 2147 91839 2175
rect 91625 2085 91653 2113
rect 91687 2085 91715 2113
rect 91749 2085 91777 2113
rect 91811 2085 91839 2113
rect 91625 2023 91653 2051
rect 91687 2023 91715 2051
rect 91749 2023 91777 2051
rect 91811 2023 91839 2051
rect 91625 1961 91653 1989
rect 91687 1961 91715 1989
rect 91749 1961 91777 1989
rect 91811 1961 91839 1989
rect 91625 -108 91653 -80
rect 91687 -108 91715 -80
rect 91749 -108 91777 -80
rect 91811 -108 91839 -80
rect 91625 -170 91653 -142
rect 91687 -170 91715 -142
rect 91749 -170 91777 -142
rect 91811 -170 91839 -142
rect 91625 -232 91653 -204
rect 91687 -232 91715 -204
rect 91749 -232 91777 -204
rect 91811 -232 91839 -204
rect 91625 -294 91653 -266
rect 91687 -294 91715 -266
rect 91749 -294 91777 -266
rect 91811 -294 91839 -266
rect 93485 41147 93513 41175
rect 93547 41147 93575 41175
rect 93609 41147 93637 41175
rect 93671 41147 93699 41175
rect 93485 41085 93513 41113
rect 93547 41085 93575 41113
rect 93609 41085 93637 41113
rect 93671 41085 93699 41113
rect 93485 41023 93513 41051
rect 93547 41023 93575 41051
rect 93609 41023 93637 41051
rect 93671 41023 93699 41051
rect 93485 40961 93513 40989
rect 93547 40961 93575 40989
rect 93609 40961 93637 40989
rect 93671 40961 93699 40989
rect 93485 32147 93513 32175
rect 93547 32147 93575 32175
rect 93609 32147 93637 32175
rect 93671 32147 93699 32175
rect 93485 32085 93513 32113
rect 93547 32085 93575 32113
rect 93609 32085 93637 32113
rect 93671 32085 93699 32113
rect 93485 32023 93513 32051
rect 93547 32023 93575 32051
rect 93609 32023 93637 32051
rect 93671 32023 93699 32051
rect 93485 31961 93513 31989
rect 93547 31961 93575 31989
rect 93609 31961 93637 31989
rect 93671 31961 93699 31989
rect 93485 23147 93513 23175
rect 93547 23147 93575 23175
rect 93609 23147 93637 23175
rect 93671 23147 93699 23175
rect 93485 23085 93513 23113
rect 93547 23085 93575 23113
rect 93609 23085 93637 23113
rect 93671 23085 93699 23113
rect 93485 23023 93513 23051
rect 93547 23023 93575 23051
rect 93609 23023 93637 23051
rect 93671 23023 93699 23051
rect 93485 22961 93513 22989
rect 93547 22961 93575 22989
rect 93609 22961 93637 22989
rect 93671 22961 93699 22989
rect 93485 14147 93513 14175
rect 93547 14147 93575 14175
rect 93609 14147 93637 14175
rect 93671 14147 93699 14175
rect 93485 14085 93513 14113
rect 93547 14085 93575 14113
rect 93609 14085 93637 14113
rect 93671 14085 93699 14113
rect 93485 14023 93513 14051
rect 93547 14023 93575 14051
rect 93609 14023 93637 14051
rect 93671 14023 93699 14051
rect 93485 13961 93513 13989
rect 93547 13961 93575 13989
rect 93609 13961 93637 13989
rect 93671 13961 93699 13989
rect 93485 5147 93513 5175
rect 93547 5147 93575 5175
rect 93609 5147 93637 5175
rect 93671 5147 93699 5175
rect 93485 5085 93513 5113
rect 93547 5085 93575 5113
rect 93609 5085 93637 5113
rect 93671 5085 93699 5113
rect 93485 5023 93513 5051
rect 93547 5023 93575 5051
rect 93609 5023 93637 5051
rect 93671 5023 93699 5051
rect 93485 4961 93513 4989
rect 93547 4961 93575 4989
rect 93609 4961 93637 4989
rect 93671 4961 93699 4989
rect 93485 -588 93513 -560
rect 93547 -588 93575 -560
rect 93609 -588 93637 -560
rect 93671 -588 93699 -560
rect 93485 -650 93513 -622
rect 93547 -650 93575 -622
rect 93609 -650 93637 -622
rect 93671 -650 93699 -622
rect 93485 -712 93513 -684
rect 93547 -712 93575 -684
rect 93609 -712 93637 -684
rect 93671 -712 93699 -684
rect 93485 -774 93513 -746
rect 93547 -774 93575 -746
rect 93609 -774 93637 -746
rect 93671 -774 93699 -746
rect 100625 47147 100653 47175
rect 100687 47147 100715 47175
rect 100749 47147 100777 47175
rect 100811 47147 100839 47175
rect 100625 47085 100653 47113
rect 100687 47085 100715 47113
rect 100749 47085 100777 47113
rect 100811 47085 100839 47113
rect 100625 47023 100653 47051
rect 100687 47023 100715 47051
rect 100749 47023 100777 47051
rect 100811 47023 100839 47051
rect 100625 46961 100653 46989
rect 100687 46961 100715 46989
rect 100749 46961 100777 46989
rect 100811 46961 100839 46989
rect 100625 38147 100653 38175
rect 100687 38147 100715 38175
rect 100749 38147 100777 38175
rect 100811 38147 100839 38175
rect 100625 38085 100653 38113
rect 100687 38085 100715 38113
rect 100749 38085 100777 38113
rect 100811 38085 100839 38113
rect 100625 38023 100653 38051
rect 100687 38023 100715 38051
rect 100749 38023 100777 38051
rect 100811 38023 100839 38051
rect 100625 37961 100653 37989
rect 100687 37961 100715 37989
rect 100749 37961 100777 37989
rect 100811 37961 100839 37989
rect 100625 29147 100653 29175
rect 100687 29147 100715 29175
rect 100749 29147 100777 29175
rect 100811 29147 100839 29175
rect 100625 29085 100653 29113
rect 100687 29085 100715 29113
rect 100749 29085 100777 29113
rect 100811 29085 100839 29113
rect 100625 29023 100653 29051
rect 100687 29023 100715 29051
rect 100749 29023 100777 29051
rect 100811 29023 100839 29051
rect 100625 28961 100653 28989
rect 100687 28961 100715 28989
rect 100749 28961 100777 28989
rect 100811 28961 100839 28989
rect 100625 20147 100653 20175
rect 100687 20147 100715 20175
rect 100749 20147 100777 20175
rect 100811 20147 100839 20175
rect 100625 20085 100653 20113
rect 100687 20085 100715 20113
rect 100749 20085 100777 20113
rect 100811 20085 100839 20113
rect 100625 20023 100653 20051
rect 100687 20023 100715 20051
rect 100749 20023 100777 20051
rect 100811 20023 100839 20051
rect 100625 19961 100653 19989
rect 100687 19961 100715 19989
rect 100749 19961 100777 19989
rect 100811 19961 100839 19989
rect 100625 11147 100653 11175
rect 100687 11147 100715 11175
rect 100749 11147 100777 11175
rect 100811 11147 100839 11175
rect 100625 11085 100653 11113
rect 100687 11085 100715 11113
rect 100749 11085 100777 11113
rect 100811 11085 100839 11113
rect 100625 11023 100653 11051
rect 100687 11023 100715 11051
rect 100749 11023 100777 11051
rect 100811 11023 100839 11051
rect 100625 10961 100653 10989
rect 100687 10961 100715 10989
rect 100749 10961 100777 10989
rect 100811 10961 100839 10989
rect 100625 2147 100653 2175
rect 100687 2147 100715 2175
rect 100749 2147 100777 2175
rect 100811 2147 100839 2175
rect 100625 2085 100653 2113
rect 100687 2085 100715 2113
rect 100749 2085 100777 2113
rect 100811 2085 100839 2113
rect 100625 2023 100653 2051
rect 100687 2023 100715 2051
rect 100749 2023 100777 2051
rect 100811 2023 100839 2051
rect 100625 1961 100653 1989
rect 100687 1961 100715 1989
rect 100749 1961 100777 1989
rect 100811 1961 100839 1989
rect 100625 -108 100653 -80
rect 100687 -108 100715 -80
rect 100749 -108 100777 -80
rect 100811 -108 100839 -80
rect 100625 -170 100653 -142
rect 100687 -170 100715 -142
rect 100749 -170 100777 -142
rect 100811 -170 100839 -142
rect 100625 -232 100653 -204
rect 100687 -232 100715 -204
rect 100749 -232 100777 -204
rect 100811 -232 100839 -204
rect 100625 -294 100653 -266
rect 100687 -294 100715 -266
rect 100749 -294 100777 -266
rect 100811 -294 100839 -266
rect 102485 41147 102513 41175
rect 102547 41147 102575 41175
rect 102609 41147 102637 41175
rect 102671 41147 102699 41175
rect 102485 41085 102513 41113
rect 102547 41085 102575 41113
rect 102609 41085 102637 41113
rect 102671 41085 102699 41113
rect 102485 41023 102513 41051
rect 102547 41023 102575 41051
rect 102609 41023 102637 41051
rect 102671 41023 102699 41051
rect 102485 40961 102513 40989
rect 102547 40961 102575 40989
rect 102609 40961 102637 40989
rect 102671 40961 102699 40989
rect 102485 32147 102513 32175
rect 102547 32147 102575 32175
rect 102609 32147 102637 32175
rect 102671 32147 102699 32175
rect 102485 32085 102513 32113
rect 102547 32085 102575 32113
rect 102609 32085 102637 32113
rect 102671 32085 102699 32113
rect 102485 32023 102513 32051
rect 102547 32023 102575 32051
rect 102609 32023 102637 32051
rect 102671 32023 102699 32051
rect 102485 31961 102513 31989
rect 102547 31961 102575 31989
rect 102609 31961 102637 31989
rect 102671 31961 102699 31989
rect 102485 23147 102513 23175
rect 102547 23147 102575 23175
rect 102609 23147 102637 23175
rect 102671 23147 102699 23175
rect 102485 23085 102513 23113
rect 102547 23085 102575 23113
rect 102609 23085 102637 23113
rect 102671 23085 102699 23113
rect 102485 23023 102513 23051
rect 102547 23023 102575 23051
rect 102609 23023 102637 23051
rect 102671 23023 102699 23051
rect 102485 22961 102513 22989
rect 102547 22961 102575 22989
rect 102609 22961 102637 22989
rect 102671 22961 102699 22989
rect 102485 14147 102513 14175
rect 102547 14147 102575 14175
rect 102609 14147 102637 14175
rect 102671 14147 102699 14175
rect 102485 14085 102513 14113
rect 102547 14085 102575 14113
rect 102609 14085 102637 14113
rect 102671 14085 102699 14113
rect 102485 14023 102513 14051
rect 102547 14023 102575 14051
rect 102609 14023 102637 14051
rect 102671 14023 102699 14051
rect 102485 13961 102513 13989
rect 102547 13961 102575 13989
rect 102609 13961 102637 13989
rect 102671 13961 102699 13989
rect 102485 5147 102513 5175
rect 102547 5147 102575 5175
rect 102609 5147 102637 5175
rect 102671 5147 102699 5175
rect 102485 5085 102513 5113
rect 102547 5085 102575 5113
rect 102609 5085 102637 5113
rect 102671 5085 102699 5113
rect 102485 5023 102513 5051
rect 102547 5023 102575 5051
rect 102609 5023 102637 5051
rect 102671 5023 102699 5051
rect 102485 4961 102513 4989
rect 102547 4961 102575 4989
rect 102609 4961 102637 4989
rect 102671 4961 102699 4989
rect 102485 -588 102513 -560
rect 102547 -588 102575 -560
rect 102609 -588 102637 -560
rect 102671 -588 102699 -560
rect 102485 -650 102513 -622
rect 102547 -650 102575 -622
rect 102609 -650 102637 -622
rect 102671 -650 102699 -622
rect 102485 -712 102513 -684
rect 102547 -712 102575 -684
rect 102609 -712 102637 -684
rect 102671 -712 102699 -684
rect 102485 -774 102513 -746
rect 102547 -774 102575 -746
rect 102609 -774 102637 -746
rect 102671 -774 102699 -746
rect 109625 47147 109653 47175
rect 109687 47147 109715 47175
rect 109749 47147 109777 47175
rect 109811 47147 109839 47175
rect 109625 47085 109653 47113
rect 109687 47085 109715 47113
rect 109749 47085 109777 47113
rect 109811 47085 109839 47113
rect 109625 47023 109653 47051
rect 109687 47023 109715 47051
rect 109749 47023 109777 47051
rect 109811 47023 109839 47051
rect 109625 46961 109653 46989
rect 109687 46961 109715 46989
rect 109749 46961 109777 46989
rect 109811 46961 109839 46989
rect 109625 38147 109653 38175
rect 109687 38147 109715 38175
rect 109749 38147 109777 38175
rect 109811 38147 109839 38175
rect 109625 38085 109653 38113
rect 109687 38085 109715 38113
rect 109749 38085 109777 38113
rect 109811 38085 109839 38113
rect 109625 38023 109653 38051
rect 109687 38023 109715 38051
rect 109749 38023 109777 38051
rect 109811 38023 109839 38051
rect 109625 37961 109653 37989
rect 109687 37961 109715 37989
rect 109749 37961 109777 37989
rect 109811 37961 109839 37989
rect 109625 29147 109653 29175
rect 109687 29147 109715 29175
rect 109749 29147 109777 29175
rect 109811 29147 109839 29175
rect 109625 29085 109653 29113
rect 109687 29085 109715 29113
rect 109749 29085 109777 29113
rect 109811 29085 109839 29113
rect 109625 29023 109653 29051
rect 109687 29023 109715 29051
rect 109749 29023 109777 29051
rect 109811 29023 109839 29051
rect 109625 28961 109653 28989
rect 109687 28961 109715 28989
rect 109749 28961 109777 28989
rect 109811 28961 109839 28989
rect 109625 20147 109653 20175
rect 109687 20147 109715 20175
rect 109749 20147 109777 20175
rect 109811 20147 109839 20175
rect 109625 20085 109653 20113
rect 109687 20085 109715 20113
rect 109749 20085 109777 20113
rect 109811 20085 109839 20113
rect 109625 20023 109653 20051
rect 109687 20023 109715 20051
rect 109749 20023 109777 20051
rect 109811 20023 109839 20051
rect 109625 19961 109653 19989
rect 109687 19961 109715 19989
rect 109749 19961 109777 19989
rect 109811 19961 109839 19989
rect 109625 11147 109653 11175
rect 109687 11147 109715 11175
rect 109749 11147 109777 11175
rect 109811 11147 109839 11175
rect 109625 11085 109653 11113
rect 109687 11085 109715 11113
rect 109749 11085 109777 11113
rect 109811 11085 109839 11113
rect 109625 11023 109653 11051
rect 109687 11023 109715 11051
rect 109749 11023 109777 11051
rect 109811 11023 109839 11051
rect 109625 10961 109653 10989
rect 109687 10961 109715 10989
rect 109749 10961 109777 10989
rect 109811 10961 109839 10989
rect 109625 2147 109653 2175
rect 109687 2147 109715 2175
rect 109749 2147 109777 2175
rect 109811 2147 109839 2175
rect 109625 2085 109653 2113
rect 109687 2085 109715 2113
rect 109749 2085 109777 2113
rect 109811 2085 109839 2113
rect 109625 2023 109653 2051
rect 109687 2023 109715 2051
rect 109749 2023 109777 2051
rect 109811 2023 109839 2051
rect 109625 1961 109653 1989
rect 109687 1961 109715 1989
rect 109749 1961 109777 1989
rect 109811 1961 109839 1989
rect 109625 -108 109653 -80
rect 109687 -108 109715 -80
rect 109749 -108 109777 -80
rect 109811 -108 109839 -80
rect 109625 -170 109653 -142
rect 109687 -170 109715 -142
rect 109749 -170 109777 -142
rect 109811 -170 109839 -142
rect 109625 -232 109653 -204
rect 109687 -232 109715 -204
rect 109749 -232 109777 -204
rect 109811 -232 109839 -204
rect 109625 -294 109653 -266
rect 109687 -294 109715 -266
rect 109749 -294 109777 -266
rect 109811 -294 109839 -266
rect 111485 41147 111513 41175
rect 111547 41147 111575 41175
rect 111609 41147 111637 41175
rect 111671 41147 111699 41175
rect 111485 41085 111513 41113
rect 111547 41085 111575 41113
rect 111609 41085 111637 41113
rect 111671 41085 111699 41113
rect 111485 41023 111513 41051
rect 111547 41023 111575 41051
rect 111609 41023 111637 41051
rect 111671 41023 111699 41051
rect 111485 40961 111513 40989
rect 111547 40961 111575 40989
rect 111609 40961 111637 40989
rect 111671 40961 111699 40989
rect 111485 32147 111513 32175
rect 111547 32147 111575 32175
rect 111609 32147 111637 32175
rect 111671 32147 111699 32175
rect 111485 32085 111513 32113
rect 111547 32085 111575 32113
rect 111609 32085 111637 32113
rect 111671 32085 111699 32113
rect 111485 32023 111513 32051
rect 111547 32023 111575 32051
rect 111609 32023 111637 32051
rect 111671 32023 111699 32051
rect 111485 31961 111513 31989
rect 111547 31961 111575 31989
rect 111609 31961 111637 31989
rect 111671 31961 111699 31989
rect 111485 23147 111513 23175
rect 111547 23147 111575 23175
rect 111609 23147 111637 23175
rect 111671 23147 111699 23175
rect 111485 23085 111513 23113
rect 111547 23085 111575 23113
rect 111609 23085 111637 23113
rect 111671 23085 111699 23113
rect 111485 23023 111513 23051
rect 111547 23023 111575 23051
rect 111609 23023 111637 23051
rect 111671 23023 111699 23051
rect 111485 22961 111513 22989
rect 111547 22961 111575 22989
rect 111609 22961 111637 22989
rect 111671 22961 111699 22989
rect 111485 14147 111513 14175
rect 111547 14147 111575 14175
rect 111609 14147 111637 14175
rect 111671 14147 111699 14175
rect 111485 14085 111513 14113
rect 111547 14085 111575 14113
rect 111609 14085 111637 14113
rect 111671 14085 111699 14113
rect 111485 14023 111513 14051
rect 111547 14023 111575 14051
rect 111609 14023 111637 14051
rect 111671 14023 111699 14051
rect 111485 13961 111513 13989
rect 111547 13961 111575 13989
rect 111609 13961 111637 13989
rect 111671 13961 111699 13989
rect 111485 5147 111513 5175
rect 111547 5147 111575 5175
rect 111609 5147 111637 5175
rect 111671 5147 111699 5175
rect 111485 5085 111513 5113
rect 111547 5085 111575 5113
rect 111609 5085 111637 5113
rect 111671 5085 111699 5113
rect 111485 5023 111513 5051
rect 111547 5023 111575 5051
rect 111609 5023 111637 5051
rect 111671 5023 111699 5051
rect 111485 4961 111513 4989
rect 111547 4961 111575 4989
rect 111609 4961 111637 4989
rect 111671 4961 111699 4989
rect 111485 -588 111513 -560
rect 111547 -588 111575 -560
rect 111609 -588 111637 -560
rect 111671 -588 111699 -560
rect 111485 -650 111513 -622
rect 111547 -650 111575 -622
rect 111609 -650 111637 -622
rect 111671 -650 111699 -622
rect 111485 -712 111513 -684
rect 111547 -712 111575 -684
rect 111609 -712 111637 -684
rect 111671 -712 111699 -684
rect 111485 -774 111513 -746
rect 111547 -774 111575 -746
rect 111609 -774 111637 -746
rect 111671 -774 111699 -746
rect 118625 47147 118653 47175
rect 118687 47147 118715 47175
rect 118749 47147 118777 47175
rect 118811 47147 118839 47175
rect 118625 47085 118653 47113
rect 118687 47085 118715 47113
rect 118749 47085 118777 47113
rect 118811 47085 118839 47113
rect 118625 47023 118653 47051
rect 118687 47023 118715 47051
rect 118749 47023 118777 47051
rect 118811 47023 118839 47051
rect 118625 46961 118653 46989
rect 118687 46961 118715 46989
rect 118749 46961 118777 46989
rect 118811 46961 118839 46989
rect 118625 38147 118653 38175
rect 118687 38147 118715 38175
rect 118749 38147 118777 38175
rect 118811 38147 118839 38175
rect 118625 38085 118653 38113
rect 118687 38085 118715 38113
rect 118749 38085 118777 38113
rect 118811 38085 118839 38113
rect 118625 38023 118653 38051
rect 118687 38023 118715 38051
rect 118749 38023 118777 38051
rect 118811 38023 118839 38051
rect 118625 37961 118653 37989
rect 118687 37961 118715 37989
rect 118749 37961 118777 37989
rect 118811 37961 118839 37989
rect 118625 29147 118653 29175
rect 118687 29147 118715 29175
rect 118749 29147 118777 29175
rect 118811 29147 118839 29175
rect 118625 29085 118653 29113
rect 118687 29085 118715 29113
rect 118749 29085 118777 29113
rect 118811 29085 118839 29113
rect 118625 29023 118653 29051
rect 118687 29023 118715 29051
rect 118749 29023 118777 29051
rect 118811 29023 118839 29051
rect 118625 28961 118653 28989
rect 118687 28961 118715 28989
rect 118749 28961 118777 28989
rect 118811 28961 118839 28989
rect 118625 20147 118653 20175
rect 118687 20147 118715 20175
rect 118749 20147 118777 20175
rect 118811 20147 118839 20175
rect 118625 20085 118653 20113
rect 118687 20085 118715 20113
rect 118749 20085 118777 20113
rect 118811 20085 118839 20113
rect 118625 20023 118653 20051
rect 118687 20023 118715 20051
rect 118749 20023 118777 20051
rect 118811 20023 118839 20051
rect 118625 19961 118653 19989
rect 118687 19961 118715 19989
rect 118749 19961 118777 19989
rect 118811 19961 118839 19989
rect 118625 11147 118653 11175
rect 118687 11147 118715 11175
rect 118749 11147 118777 11175
rect 118811 11147 118839 11175
rect 118625 11085 118653 11113
rect 118687 11085 118715 11113
rect 118749 11085 118777 11113
rect 118811 11085 118839 11113
rect 118625 11023 118653 11051
rect 118687 11023 118715 11051
rect 118749 11023 118777 11051
rect 118811 11023 118839 11051
rect 118625 10961 118653 10989
rect 118687 10961 118715 10989
rect 118749 10961 118777 10989
rect 118811 10961 118839 10989
rect 118625 2147 118653 2175
rect 118687 2147 118715 2175
rect 118749 2147 118777 2175
rect 118811 2147 118839 2175
rect 118625 2085 118653 2113
rect 118687 2085 118715 2113
rect 118749 2085 118777 2113
rect 118811 2085 118839 2113
rect 118625 2023 118653 2051
rect 118687 2023 118715 2051
rect 118749 2023 118777 2051
rect 118811 2023 118839 2051
rect 118625 1961 118653 1989
rect 118687 1961 118715 1989
rect 118749 1961 118777 1989
rect 118811 1961 118839 1989
rect 118625 -108 118653 -80
rect 118687 -108 118715 -80
rect 118749 -108 118777 -80
rect 118811 -108 118839 -80
rect 118625 -170 118653 -142
rect 118687 -170 118715 -142
rect 118749 -170 118777 -142
rect 118811 -170 118839 -142
rect 118625 -232 118653 -204
rect 118687 -232 118715 -204
rect 118749 -232 118777 -204
rect 118811 -232 118839 -204
rect 118625 -294 118653 -266
rect 118687 -294 118715 -266
rect 118749 -294 118777 -266
rect 118811 -294 118839 -266
rect 120485 41147 120513 41175
rect 120547 41147 120575 41175
rect 120609 41147 120637 41175
rect 120671 41147 120699 41175
rect 120485 41085 120513 41113
rect 120547 41085 120575 41113
rect 120609 41085 120637 41113
rect 120671 41085 120699 41113
rect 120485 41023 120513 41051
rect 120547 41023 120575 41051
rect 120609 41023 120637 41051
rect 120671 41023 120699 41051
rect 120485 40961 120513 40989
rect 120547 40961 120575 40989
rect 120609 40961 120637 40989
rect 120671 40961 120699 40989
rect 120485 32147 120513 32175
rect 120547 32147 120575 32175
rect 120609 32147 120637 32175
rect 120671 32147 120699 32175
rect 120485 32085 120513 32113
rect 120547 32085 120575 32113
rect 120609 32085 120637 32113
rect 120671 32085 120699 32113
rect 120485 32023 120513 32051
rect 120547 32023 120575 32051
rect 120609 32023 120637 32051
rect 120671 32023 120699 32051
rect 120485 31961 120513 31989
rect 120547 31961 120575 31989
rect 120609 31961 120637 31989
rect 120671 31961 120699 31989
rect 120485 23147 120513 23175
rect 120547 23147 120575 23175
rect 120609 23147 120637 23175
rect 120671 23147 120699 23175
rect 120485 23085 120513 23113
rect 120547 23085 120575 23113
rect 120609 23085 120637 23113
rect 120671 23085 120699 23113
rect 120485 23023 120513 23051
rect 120547 23023 120575 23051
rect 120609 23023 120637 23051
rect 120671 23023 120699 23051
rect 120485 22961 120513 22989
rect 120547 22961 120575 22989
rect 120609 22961 120637 22989
rect 120671 22961 120699 22989
rect 120485 14147 120513 14175
rect 120547 14147 120575 14175
rect 120609 14147 120637 14175
rect 120671 14147 120699 14175
rect 120485 14085 120513 14113
rect 120547 14085 120575 14113
rect 120609 14085 120637 14113
rect 120671 14085 120699 14113
rect 120485 14023 120513 14051
rect 120547 14023 120575 14051
rect 120609 14023 120637 14051
rect 120671 14023 120699 14051
rect 120485 13961 120513 13989
rect 120547 13961 120575 13989
rect 120609 13961 120637 13989
rect 120671 13961 120699 13989
rect 120485 5147 120513 5175
rect 120547 5147 120575 5175
rect 120609 5147 120637 5175
rect 120671 5147 120699 5175
rect 120485 5085 120513 5113
rect 120547 5085 120575 5113
rect 120609 5085 120637 5113
rect 120671 5085 120699 5113
rect 120485 5023 120513 5051
rect 120547 5023 120575 5051
rect 120609 5023 120637 5051
rect 120671 5023 120699 5051
rect 120485 4961 120513 4989
rect 120547 4961 120575 4989
rect 120609 4961 120637 4989
rect 120671 4961 120699 4989
rect 120485 -588 120513 -560
rect 120547 -588 120575 -560
rect 120609 -588 120637 -560
rect 120671 -588 120699 -560
rect 120485 -650 120513 -622
rect 120547 -650 120575 -622
rect 120609 -650 120637 -622
rect 120671 -650 120699 -622
rect 120485 -712 120513 -684
rect 120547 -712 120575 -684
rect 120609 -712 120637 -684
rect 120671 -712 120699 -684
rect 120485 -774 120513 -746
rect 120547 -774 120575 -746
rect 120609 -774 120637 -746
rect 120671 -774 120699 -746
rect 127625 119147 127653 119175
rect 127687 119147 127715 119175
rect 127749 119147 127777 119175
rect 127811 119147 127839 119175
rect 127625 119085 127653 119113
rect 127687 119085 127715 119113
rect 127749 119085 127777 119113
rect 127811 119085 127839 119113
rect 127625 119023 127653 119051
rect 127687 119023 127715 119051
rect 127749 119023 127777 119051
rect 127811 119023 127839 119051
rect 127625 118961 127653 118989
rect 127687 118961 127715 118989
rect 127749 118961 127777 118989
rect 127811 118961 127839 118989
rect 127625 110147 127653 110175
rect 127687 110147 127715 110175
rect 127749 110147 127777 110175
rect 127811 110147 127839 110175
rect 127625 110085 127653 110113
rect 127687 110085 127715 110113
rect 127749 110085 127777 110113
rect 127811 110085 127839 110113
rect 127625 110023 127653 110051
rect 127687 110023 127715 110051
rect 127749 110023 127777 110051
rect 127811 110023 127839 110051
rect 127625 109961 127653 109989
rect 127687 109961 127715 109989
rect 127749 109961 127777 109989
rect 127811 109961 127839 109989
rect 127625 101147 127653 101175
rect 127687 101147 127715 101175
rect 127749 101147 127777 101175
rect 127811 101147 127839 101175
rect 127625 101085 127653 101113
rect 127687 101085 127715 101113
rect 127749 101085 127777 101113
rect 127811 101085 127839 101113
rect 127625 101023 127653 101051
rect 127687 101023 127715 101051
rect 127749 101023 127777 101051
rect 127811 101023 127839 101051
rect 127625 100961 127653 100989
rect 127687 100961 127715 100989
rect 127749 100961 127777 100989
rect 127811 100961 127839 100989
rect 127625 92147 127653 92175
rect 127687 92147 127715 92175
rect 127749 92147 127777 92175
rect 127811 92147 127839 92175
rect 127625 92085 127653 92113
rect 127687 92085 127715 92113
rect 127749 92085 127777 92113
rect 127811 92085 127839 92113
rect 127625 92023 127653 92051
rect 127687 92023 127715 92051
rect 127749 92023 127777 92051
rect 127811 92023 127839 92051
rect 127625 91961 127653 91989
rect 127687 91961 127715 91989
rect 127749 91961 127777 91989
rect 127811 91961 127839 91989
rect 127625 83147 127653 83175
rect 127687 83147 127715 83175
rect 127749 83147 127777 83175
rect 127811 83147 127839 83175
rect 127625 83085 127653 83113
rect 127687 83085 127715 83113
rect 127749 83085 127777 83113
rect 127811 83085 127839 83113
rect 127625 83023 127653 83051
rect 127687 83023 127715 83051
rect 127749 83023 127777 83051
rect 127811 83023 127839 83051
rect 127625 82961 127653 82989
rect 127687 82961 127715 82989
rect 127749 82961 127777 82989
rect 127811 82961 127839 82989
rect 127625 74147 127653 74175
rect 127687 74147 127715 74175
rect 127749 74147 127777 74175
rect 127811 74147 127839 74175
rect 127625 74085 127653 74113
rect 127687 74085 127715 74113
rect 127749 74085 127777 74113
rect 127811 74085 127839 74113
rect 127625 74023 127653 74051
rect 127687 74023 127715 74051
rect 127749 74023 127777 74051
rect 127811 74023 127839 74051
rect 127625 73961 127653 73989
rect 127687 73961 127715 73989
rect 127749 73961 127777 73989
rect 127811 73961 127839 73989
rect 127625 65147 127653 65175
rect 127687 65147 127715 65175
rect 127749 65147 127777 65175
rect 127811 65147 127839 65175
rect 127625 65085 127653 65113
rect 127687 65085 127715 65113
rect 127749 65085 127777 65113
rect 127811 65085 127839 65113
rect 127625 65023 127653 65051
rect 127687 65023 127715 65051
rect 127749 65023 127777 65051
rect 127811 65023 127839 65051
rect 127625 64961 127653 64989
rect 127687 64961 127715 64989
rect 127749 64961 127777 64989
rect 127811 64961 127839 64989
rect 127625 56147 127653 56175
rect 127687 56147 127715 56175
rect 127749 56147 127777 56175
rect 127811 56147 127839 56175
rect 127625 56085 127653 56113
rect 127687 56085 127715 56113
rect 127749 56085 127777 56113
rect 127811 56085 127839 56113
rect 127625 56023 127653 56051
rect 127687 56023 127715 56051
rect 127749 56023 127777 56051
rect 127811 56023 127839 56051
rect 127625 55961 127653 55989
rect 127687 55961 127715 55989
rect 127749 55961 127777 55989
rect 127811 55961 127839 55989
rect 127625 47147 127653 47175
rect 127687 47147 127715 47175
rect 127749 47147 127777 47175
rect 127811 47147 127839 47175
rect 127625 47085 127653 47113
rect 127687 47085 127715 47113
rect 127749 47085 127777 47113
rect 127811 47085 127839 47113
rect 127625 47023 127653 47051
rect 127687 47023 127715 47051
rect 127749 47023 127777 47051
rect 127811 47023 127839 47051
rect 127625 46961 127653 46989
rect 127687 46961 127715 46989
rect 127749 46961 127777 46989
rect 127811 46961 127839 46989
rect 127625 38147 127653 38175
rect 127687 38147 127715 38175
rect 127749 38147 127777 38175
rect 127811 38147 127839 38175
rect 127625 38085 127653 38113
rect 127687 38085 127715 38113
rect 127749 38085 127777 38113
rect 127811 38085 127839 38113
rect 127625 38023 127653 38051
rect 127687 38023 127715 38051
rect 127749 38023 127777 38051
rect 127811 38023 127839 38051
rect 127625 37961 127653 37989
rect 127687 37961 127715 37989
rect 127749 37961 127777 37989
rect 127811 37961 127839 37989
rect 127625 29147 127653 29175
rect 127687 29147 127715 29175
rect 127749 29147 127777 29175
rect 127811 29147 127839 29175
rect 127625 29085 127653 29113
rect 127687 29085 127715 29113
rect 127749 29085 127777 29113
rect 127811 29085 127839 29113
rect 127625 29023 127653 29051
rect 127687 29023 127715 29051
rect 127749 29023 127777 29051
rect 127811 29023 127839 29051
rect 127625 28961 127653 28989
rect 127687 28961 127715 28989
rect 127749 28961 127777 28989
rect 127811 28961 127839 28989
rect 127625 20147 127653 20175
rect 127687 20147 127715 20175
rect 127749 20147 127777 20175
rect 127811 20147 127839 20175
rect 127625 20085 127653 20113
rect 127687 20085 127715 20113
rect 127749 20085 127777 20113
rect 127811 20085 127839 20113
rect 127625 20023 127653 20051
rect 127687 20023 127715 20051
rect 127749 20023 127777 20051
rect 127811 20023 127839 20051
rect 127625 19961 127653 19989
rect 127687 19961 127715 19989
rect 127749 19961 127777 19989
rect 127811 19961 127839 19989
rect 127625 11147 127653 11175
rect 127687 11147 127715 11175
rect 127749 11147 127777 11175
rect 127811 11147 127839 11175
rect 127625 11085 127653 11113
rect 127687 11085 127715 11113
rect 127749 11085 127777 11113
rect 127811 11085 127839 11113
rect 127625 11023 127653 11051
rect 127687 11023 127715 11051
rect 127749 11023 127777 11051
rect 127811 11023 127839 11051
rect 127625 10961 127653 10989
rect 127687 10961 127715 10989
rect 127749 10961 127777 10989
rect 127811 10961 127839 10989
rect 127625 2147 127653 2175
rect 127687 2147 127715 2175
rect 127749 2147 127777 2175
rect 127811 2147 127839 2175
rect 127625 2085 127653 2113
rect 127687 2085 127715 2113
rect 127749 2085 127777 2113
rect 127811 2085 127839 2113
rect 127625 2023 127653 2051
rect 127687 2023 127715 2051
rect 127749 2023 127777 2051
rect 127811 2023 127839 2051
rect 127625 1961 127653 1989
rect 127687 1961 127715 1989
rect 127749 1961 127777 1989
rect 127811 1961 127839 1989
rect 127625 -108 127653 -80
rect 127687 -108 127715 -80
rect 127749 -108 127777 -80
rect 127811 -108 127839 -80
rect 127625 -170 127653 -142
rect 127687 -170 127715 -142
rect 127749 -170 127777 -142
rect 127811 -170 127839 -142
rect 127625 -232 127653 -204
rect 127687 -232 127715 -204
rect 127749 -232 127777 -204
rect 127811 -232 127839 -204
rect 127625 -294 127653 -266
rect 127687 -294 127715 -266
rect 127749 -294 127777 -266
rect 127811 -294 127839 -266
rect 129485 122147 129513 122175
rect 129547 122147 129575 122175
rect 129609 122147 129637 122175
rect 129671 122147 129699 122175
rect 129485 122085 129513 122113
rect 129547 122085 129575 122113
rect 129609 122085 129637 122113
rect 129671 122085 129699 122113
rect 129485 122023 129513 122051
rect 129547 122023 129575 122051
rect 129609 122023 129637 122051
rect 129671 122023 129699 122051
rect 129485 121961 129513 121989
rect 129547 121961 129575 121989
rect 129609 121961 129637 121989
rect 129671 121961 129699 121989
rect 129485 113147 129513 113175
rect 129547 113147 129575 113175
rect 129609 113147 129637 113175
rect 129671 113147 129699 113175
rect 129485 113085 129513 113113
rect 129547 113085 129575 113113
rect 129609 113085 129637 113113
rect 129671 113085 129699 113113
rect 129485 113023 129513 113051
rect 129547 113023 129575 113051
rect 129609 113023 129637 113051
rect 129671 113023 129699 113051
rect 129485 112961 129513 112989
rect 129547 112961 129575 112989
rect 129609 112961 129637 112989
rect 129671 112961 129699 112989
rect 129485 104147 129513 104175
rect 129547 104147 129575 104175
rect 129609 104147 129637 104175
rect 129671 104147 129699 104175
rect 129485 104085 129513 104113
rect 129547 104085 129575 104113
rect 129609 104085 129637 104113
rect 129671 104085 129699 104113
rect 129485 104023 129513 104051
rect 129547 104023 129575 104051
rect 129609 104023 129637 104051
rect 129671 104023 129699 104051
rect 129485 103961 129513 103989
rect 129547 103961 129575 103989
rect 129609 103961 129637 103989
rect 129671 103961 129699 103989
rect 129485 95147 129513 95175
rect 129547 95147 129575 95175
rect 129609 95147 129637 95175
rect 129671 95147 129699 95175
rect 129485 95085 129513 95113
rect 129547 95085 129575 95113
rect 129609 95085 129637 95113
rect 129671 95085 129699 95113
rect 129485 95023 129513 95051
rect 129547 95023 129575 95051
rect 129609 95023 129637 95051
rect 129671 95023 129699 95051
rect 129485 94961 129513 94989
rect 129547 94961 129575 94989
rect 129609 94961 129637 94989
rect 129671 94961 129699 94989
rect 129485 86147 129513 86175
rect 129547 86147 129575 86175
rect 129609 86147 129637 86175
rect 129671 86147 129699 86175
rect 129485 86085 129513 86113
rect 129547 86085 129575 86113
rect 129609 86085 129637 86113
rect 129671 86085 129699 86113
rect 129485 86023 129513 86051
rect 129547 86023 129575 86051
rect 129609 86023 129637 86051
rect 129671 86023 129699 86051
rect 129485 85961 129513 85989
rect 129547 85961 129575 85989
rect 129609 85961 129637 85989
rect 129671 85961 129699 85989
rect 129485 77147 129513 77175
rect 129547 77147 129575 77175
rect 129609 77147 129637 77175
rect 129671 77147 129699 77175
rect 129485 77085 129513 77113
rect 129547 77085 129575 77113
rect 129609 77085 129637 77113
rect 129671 77085 129699 77113
rect 129485 77023 129513 77051
rect 129547 77023 129575 77051
rect 129609 77023 129637 77051
rect 129671 77023 129699 77051
rect 129485 76961 129513 76989
rect 129547 76961 129575 76989
rect 129609 76961 129637 76989
rect 129671 76961 129699 76989
rect 129485 68147 129513 68175
rect 129547 68147 129575 68175
rect 129609 68147 129637 68175
rect 129671 68147 129699 68175
rect 129485 68085 129513 68113
rect 129547 68085 129575 68113
rect 129609 68085 129637 68113
rect 129671 68085 129699 68113
rect 129485 68023 129513 68051
rect 129547 68023 129575 68051
rect 129609 68023 129637 68051
rect 129671 68023 129699 68051
rect 129485 67961 129513 67989
rect 129547 67961 129575 67989
rect 129609 67961 129637 67989
rect 129671 67961 129699 67989
rect 129485 59147 129513 59175
rect 129547 59147 129575 59175
rect 129609 59147 129637 59175
rect 129671 59147 129699 59175
rect 129485 59085 129513 59113
rect 129547 59085 129575 59113
rect 129609 59085 129637 59113
rect 129671 59085 129699 59113
rect 129485 59023 129513 59051
rect 129547 59023 129575 59051
rect 129609 59023 129637 59051
rect 129671 59023 129699 59051
rect 129485 58961 129513 58989
rect 129547 58961 129575 58989
rect 129609 58961 129637 58989
rect 129671 58961 129699 58989
rect 129485 50147 129513 50175
rect 129547 50147 129575 50175
rect 129609 50147 129637 50175
rect 129671 50147 129699 50175
rect 129485 50085 129513 50113
rect 129547 50085 129575 50113
rect 129609 50085 129637 50113
rect 129671 50085 129699 50113
rect 129485 50023 129513 50051
rect 129547 50023 129575 50051
rect 129609 50023 129637 50051
rect 129671 50023 129699 50051
rect 129485 49961 129513 49989
rect 129547 49961 129575 49989
rect 129609 49961 129637 49989
rect 129671 49961 129699 49989
rect 129485 41147 129513 41175
rect 129547 41147 129575 41175
rect 129609 41147 129637 41175
rect 129671 41147 129699 41175
rect 129485 41085 129513 41113
rect 129547 41085 129575 41113
rect 129609 41085 129637 41113
rect 129671 41085 129699 41113
rect 129485 41023 129513 41051
rect 129547 41023 129575 41051
rect 129609 41023 129637 41051
rect 129671 41023 129699 41051
rect 129485 40961 129513 40989
rect 129547 40961 129575 40989
rect 129609 40961 129637 40989
rect 129671 40961 129699 40989
rect 129485 32147 129513 32175
rect 129547 32147 129575 32175
rect 129609 32147 129637 32175
rect 129671 32147 129699 32175
rect 129485 32085 129513 32113
rect 129547 32085 129575 32113
rect 129609 32085 129637 32113
rect 129671 32085 129699 32113
rect 129485 32023 129513 32051
rect 129547 32023 129575 32051
rect 129609 32023 129637 32051
rect 129671 32023 129699 32051
rect 129485 31961 129513 31989
rect 129547 31961 129575 31989
rect 129609 31961 129637 31989
rect 129671 31961 129699 31989
rect 129485 23147 129513 23175
rect 129547 23147 129575 23175
rect 129609 23147 129637 23175
rect 129671 23147 129699 23175
rect 129485 23085 129513 23113
rect 129547 23085 129575 23113
rect 129609 23085 129637 23113
rect 129671 23085 129699 23113
rect 129485 23023 129513 23051
rect 129547 23023 129575 23051
rect 129609 23023 129637 23051
rect 129671 23023 129699 23051
rect 129485 22961 129513 22989
rect 129547 22961 129575 22989
rect 129609 22961 129637 22989
rect 129671 22961 129699 22989
rect 129485 14147 129513 14175
rect 129547 14147 129575 14175
rect 129609 14147 129637 14175
rect 129671 14147 129699 14175
rect 129485 14085 129513 14113
rect 129547 14085 129575 14113
rect 129609 14085 129637 14113
rect 129671 14085 129699 14113
rect 129485 14023 129513 14051
rect 129547 14023 129575 14051
rect 129609 14023 129637 14051
rect 129671 14023 129699 14051
rect 129485 13961 129513 13989
rect 129547 13961 129575 13989
rect 129609 13961 129637 13989
rect 129671 13961 129699 13989
rect 129485 5147 129513 5175
rect 129547 5147 129575 5175
rect 129609 5147 129637 5175
rect 129671 5147 129699 5175
rect 129485 5085 129513 5113
rect 129547 5085 129575 5113
rect 129609 5085 129637 5113
rect 129671 5085 129699 5113
rect 129485 5023 129513 5051
rect 129547 5023 129575 5051
rect 129609 5023 129637 5051
rect 129671 5023 129699 5051
rect 129485 4961 129513 4989
rect 129547 4961 129575 4989
rect 129609 4961 129637 4989
rect 129671 4961 129699 4989
rect 129485 -588 129513 -560
rect 129547 -588 129575 -560
rect 129609 -588 129637 -560
rect 129671 -588 129699 -560
rect 129485 -650 129513 -622
rect 129547 -650 129575 -622
rect 129609 -650 129637 -622
rect 129671 -650 129699 -622
rect 129485 -712 129513 -684
rect 129547 -712 129575 -684
rect 129609 -712 129637 -684
rect 129671 -712 129699 -684
rect 129485 -774 129513 -746
rect 129547 -774 129575 -746
rect 129609 -774 129637 -746
rect 129671 -774 129699 -746
rect 136625 119147 136653 119175
rect 136687 119147 136715 119175
rect 136749 119147 136777 119175
rect 136811 119147 136839 119175
rect 136625 119085 136653 119113
rect 136687 119085 136715 119113
rect 136749 119085 136777 119113
rect 136811 119085 136839 119113
rect 136625 119023 136653 119051
rect 136687 119023 136715 119051
rect 136749 119023 136777 119051
rect 136811 119023 136839 119051
rect 136625 118961 136653 118989
rect 136687 118961 136715 118989
rect 136749 118961 136777 118989
rect 136811 118961 136839 118989
rect 136625 110147 136653 110175
rect 136687 110147 136715 110175
rect 136749 110147 136777 110175
rect 136811 110147 136839 110175
rect 136625 110085 136653 110113
rect 136687 110085 136715 110113
rect 136749 110085 136777 110113
rect 136811 110085 136839 110113
rect 136625 110023 136653 110051
rect 136687 110023 136715 110051
rect 136749 110023 136777 110051
rect 136811 110023 136839 110051
rect 136625 109961 136653 109989
rect 136687 109961 136715 109989
rect 136749 109961 136777 109989
rect 136811 109961 136839 109989
rect 136625 101147 136653 101175
rect 136687 101147 136715 101175
rect 136749 101147 136777 101175
rect 136811 101147 136839 101175
rect 136625 101085 136653 101113
rect 136687 101085 136715 101113
rect 136749 101085 136777 101113
rect 136811 101085 136839 101113
rect 136625 101023 136653 101051
rect 136687 101023 136715 101051
rect 136749 101023 136777 101051
rect 136811 101023 136839 101051
rect 136625 100961 136653 100989
rect 136687 100961 136715 100989
rect 136749 100961 136777 100989
rect 136811 100961 136839 100989
rect 136625 92147 136653 92175
rect 136687 92147 136715 92175
rect 136749 92147 136777 92175
rect 136811 92147 136839 92175
rect 136625 92085 136653 92113
rect 136687 92085 136715 92113
rect 136749 92085 136777 92113
rect 136811 92085 136839 92113
rect 136625 92023 136653 92051
rect 136687 92023 136715 92051
rect 136749 92023 136777 92051
rect 136811 92023 136839 92051
rect 136625 91961 136653 91989
rect 136687 91961 136715 91989
rect 136749 91961 136777 91989
rect 136811 91961 136839 91989
rect 136625 83147 136653 83175
rect 136687 83147 136715 83175
rect 136749 83147 136777 83175
rect 136811 83147 136839 83175
rect 136625 83085 136653 83113
rect 136687 83085 136715 83113
rect 136749 83085 136777 83113
rect 136811 83085 136839 83113
rect 136625 83023 136653 83051
rect 136687 83023 136715 83051
rect 136749 83023 136777 83051
rect 136811 83023 136839 83051
rect 136625 82961 136653 82989
rect 136687 82961 136715 82989
rect 136749 82961 136777 82989
rect 136811 82961 136839 82989
rect 136625 74147 136653 74175
rect 136687 74147 136715 74175
rect 136749 74147 136777 74175
rect 136811 74147 136839 74175
rect 136625 74085 136653 74113
rect 136687 74085 136715 74113
rect 136749 74085 136777 74113
rect 136811 74085 136839 74113
rect 136625 74023 136653 74051
rect 136687 74023 136715 74051
rect 136749 74023 136777 74051
rect 136811 74023 136839 74051
rect 136625 73961 136653 73989
rect 136687 73961 136715 73989
rect 136749 73961 136777 73989
rect 136811 73961 136839 73989
rect 136625 65147 136653 65175
rect 136687 65147 136715 65175
rect 136749 65147 136777 65175
rect 136811 65147 136839 65175
rect 136625 65085 136653 65113
rect 136687 65085 136715 65113
rect 136749 65085 136777 65113
rect 136811 65085 136839 65113
rect 136625 65023 136653 65051
rect 136687 65023 136715 65051
rect 136749 65023 136777 65051
rect 136811 65023 136839 65051
rect 136625 64961 136653 64989
rect 136687 64961 136715 64989
rect 136749 64961 136777 64989
rect 136811 64961 136839 64989
rect 136625 56147 136653 56175
rect 136687 56147 136715 56175
rect 136749 56147 136777 56175
rect 136811 56147 136839 56175
rect 136625 56085 136653 56113
rect 136687 56085 136715 56113
rect 136749 56085 136777 56113
rect 136811 56085 136839 56113
rect 136625 56023 136653 56051
rect 136687 56023 136715 56051
rect 136749 56023 136777 56051
rect 136811 56023 136839 56051
rect 136625 55961 136653 55989
rect 136687 55961 136715 55989
rect 136749 55961 136777 55989
rect 136811 55961 136839 55989
rect 136625 47147 136653 47175
rect 136687 47147 136715 47175
rect 136749 47147 136777 47175
rect 136811 47147 136839 47175
rect 136625 47085 136653 47113
rect 136687 47085 136715 47113
rect 136749 47085 136777 47113
rect 136811 47085 136839 47113
rect 136625 47023 136653 47051
rect 136687 47023 136715 47051
rect 136749 47023 136777 47051
rect 136811 47023 136839 47051
rect 136625 46961 136653 46989
rect 136687 46961 136715 46989
rect 136749 46961 136777 46989
rect 136811 46961 136839 46989
rect 136625 38147 136653 38175
rect 136687 38147 136715 38175
rect 136749 38147 136777 38175
rect 136811 38147 136839 38175
rect 136625 38085 136653 38113
rect 136687 38085 136715 38113
rect 136749 38085 136777 38113
rect 136811 38085 136839 38113
rect 136625 38023 136653 38051
rect 136687 38023 136715 38051
rect 136749 38023 136777 38051
rect 136811 38023 136839 38051
rect 136625 37961 136653 37989
rect 136687 37961 136715 37989
rect 136749 37961 136777 37989
rect 136811 37961 136839 37989
rect 136625 29147 136653 29175
rect 136687 29147 136715 29175
rect 136749 29147 136777 29175
rect 136811 29147 136839 29175
rect 136625 29085 136653 29113
rect 136687 29085 136715 29113
rect 136749 29085 136777 29113
rect 136811 29085 136839 29113
rect 136625 29023 136653 29051
rect 136687 29023 136715 29051
rect 136749 29023 136777 29051
rect 136811 29023 136839 29051
rect 136625 28961 136653 28989
rect 136687 28961 136715 28989
rect 136749 28961 136777 28989
rect 136811 28961 136839 28989
rect 136625 20147 136653 20175
rect 136687 20147 136715 20175
rect 136749 20147 136777 20175
rect 136811 20147 136839 20175
rect 136625 20085 136653 20113
rect 136687 20085 136715 20113
rect 136749 20085 136777 20113
rect 136811 20085 136839 20113
rect 136625 20023 136653 20051
rect 136687 20023 136715 20051
rect 136749 20023 136777 20051
rect 136811 20023 136839 20051
rect 136625 19961 136653 19989
rect 136687 19961 136715 19989
rect 136749 19961 136777 19989
rect 136811 19961 136839 19989
rect 136625 11147 136653 11175
rect 136687 11147 136715 11175
rect 136749 11147 136777 11175
rect 136811 11147 136839 11175
rect 136625 11085 136653 11113
rect 136687 11085 136715 11113
rect 136749 11085 136777 11113
rect 136811 11085 136839 11113
rect 136625 11023 136653 11051
rect 136687 11023 136715 11051
rect 136749 11023 136777 11051
rect 136811 11023 136839 11051
rect 136625 10961 136653 10989
rect 136687 10961 136715 10989
rect 136749 10961 136777 10989
rect 136811 10961 136839 10989
rect 136625 2147 136653 2175
rect 136687 2147 136715 2175
rect 136749 2147 136777 2175
rect 136811 2147 136839 2175
rect 136625 2085 136653 2113
rect 136687 2085 136715 2113
rect 136749 2085 136777 2113
rect 136811 2085 136839 2113
rect 136625 2023 136653 2051
rect 136687 2023 136715 2051
rect 136749 2023 136777 2051
rect 136811 2023 136839 2051
rect 136625 1961 136653 1989
rect 136687 1961 136715 1989
rect 136749 1961 136777 1989
rect 136811 1961 136839 1989
rect 136625 -108 136653 -80
rect 136687 -108 136715 -80
rect 136749 -108 136777 -80
rect 136811 -108 136839 -80
rect 136625 -170 136653 -142
rect 136687 -170 136715 -142
rect 136749 -170 136777 -142
rect 136811 -170 136839 -142
rect 136625 -232 136653 -204
rect 136687 -232 136715 -204
rect 136749 -232 136777 -204
rect 136811 -232 136839 -204
rect 136625 -294 136653 -266
rect 136687 -294 136715 -266
rect 136749 -294 136777 -266
rect 136811 -294 136839 -266
rect 138485 122147 138513 122175
rect 138547 122147 138575 122175
rect 138609 122147 138637 122175
rect 138671 122147 138699 122175
rect 138485 122085 138513 122113
rect 138547 122085 138575 122113
rect 138609 122085 138637 122113
rect 138671 122085 138699 122113
rect 138485 122023 138513 122051
rect 138547 122023 138575 122051
rect 138609 122023 138637 122051
rect 138671 122023 138699 122051
rect 138485 121961 138513 121989
rect 138547 121961 138575 121989
rect 138609 121961 138637 121989
rect 138671 121961 138699 121989
rect 138485 113147 138513 113175
rect 138547 113147 138575 113175
rect 138609 113147 138637 113175
rect 138671 113147 138699 113175
rect 138485 113085 138513 113113
rect 138547 113085 138575 113113
rect 138609 113085 138637 113113
rect 138671 113085 138699 113113
rect 138485 113023 138513 113051
rect 138547 113023 138575 113051
rect 138609 113023 138637 113051
rect 138671 113023 138699 113051
rect 138485 112961 138513 112989
rect 138547 112961 138575 112989
rect 138609 112961 138637 112989
rect 138671 112961 138699 112989
rect 138485 104147 138513 104175
rect 138547 104147 138575 104175
rect 138609 104147 138637 104175
rect 138671 104147 138699 104175
rect 138485 104085 138513 104113
rect 138547 104085 138575 104113
rect 138609 104085 138637 104113
rect 138671 104085 138699 104113
rect 138485 104023 138513 104051
rect 138547 104023 138575 104051
rect 138609 104023 138637 104051
rect 138671 104023 138699 104051
rect 138485 103961 138513 103989
rect 138547 103961 138575 103989
rect 138609 103961 138637 103989
rect 138671 103961 138699 103989
rect 138485 95147 138513 95175
rect 138547 95147 138575 95175
rect 138609 95147 138637 95175
rect 138671 95147 138699 95175
rect 138485 95085 138513 95113
rect 138547 95085 138575 95113
rect 138609 95085 138637 95113
rect 138671 95085 138699 95113
rect 138485 95023 138513 95051
rect 138547 95023 138575 95051
rect 138609 95023 138637 95051
rect 138671 95023 138699 95051
rect 138485 94961 138513 94989
rect 138547 94961 138575 94989
rect 138609 94961 138637 94989
rect 138671 94961 138699 94989
rect 138485 86147 138513 86175
rect 138547 86147 138575 86175
rect 138609 86147 138637 86175
rect 138671 86147 138699 86175
rect 138485 86085 138513 86113
rect 138547 86085 138575 86113
rect 138609 86085 138637 86113
rect 138671 86085 138699 86113
rect 138485 86023 138513 86051
rect 138547 86023 138575 86051
rect 138609 86023 138637 86051
rect 138671 86023 138699 86051
rect 138485 85961 138513 85989
rect 138547 85961 138575 85989
rect 138609 85961 138637 85989
rect 138671 85961 138699 85989
rect 138485 77147 138513 77175
rect 138547 77147 138575 77175
rect 138609 77147 138637 77175
rect 138671 77147 138699 77175
rect 138485 77085 138513 77113
rect 138547 77085 138575 77113
rect 138609 77085 138637 77113
rect 138671 77085 138699 77113
rect 138485 77023 138513 77051
rect 138547 77023 138575 77051
rect 138609 77023 138637 77051
rect 138671 77023 138699 77051
rect 138485 76961 138513 76989
rect 138547 76961 138575 76989
rect 138609 76961 138637 76989
rect 138671 76961 138699 76989
rect 138485 68147 138513 68175
rect 138547 68147 138575 68175
rect 138609 68147 138637 68175
rect 138671 68147 138699 68175
rect 138485 68085 138513 68113
rect 138547 68085 138575 68113
rect 138609 68085 138637 68113
rect 138671 68085 138699 68113
rect 138485 68023 138513 68051
rect 138547 68023 138575 68051
rect 138609 68023 138637 68051
rect 138671 68023 138699 68051
rect 138485 67961 138513 67989
rect 138547 67961 138575 67989
rect 138609 67961 138637 67989
rect 138671 67961 138699 67989
rect 138485 59147 138513 59175
rect 138547 59147 138575 59175
rect 138609 59147 138637 59175
rect 138671 59147 138699 59175
rect 138485 59085 138513 59113
rect 138547 59085 138575 59113
rect 138609 59085 138637 59113
rect 138671 59085 138699 59113
rect 138485 59023 138513 59051
rect 138547 59023 138575 59051
rect 138609 59023 138637 59051
rect 138671 59023 138699 59051
rect 138485 58961 138513 58989
rect 138547 58961 138575 58989
rect 138609 58961 138637 58989
rect 138671 58961 138699 58989
rect 138485 50147 138513 50175
rect 138547 50147 138575 50175
rect 138609 50147 138637 50175
rect 138671 50147 138699 50175
rect 138485 50085 138513 50113
rect 138547 50085 138575 50113
rect 138609 50085 138637 50113
rect 138671 50085 138699 50113
rect 138485 50023 138513 50051
rect 138547 50023 138575 50051
rect 138609 50023 138637 50051
rect 138671 50023 138699 50051
rect 138485 49961 138513 49989
rect 138547 49961 138575 49989
rect 138609 49961 138637 49989
rect 138671 49961 138699 49989
rect 138485 41147 138513 41175
rect 138547 41147 138575 41175
rect 138609 41147 138637 41175
rect 138671 41147 138699 41175
rect 138485 41085 138513 41113
rect 138547 41085 138575 41113
rect 138609 41085 138637 41113
rect 138671 41085 138699 41113
rect 138485 41023 138513 41051
rect 138547 41023 138575 41051
rect 138609 41023 138637 41051
rect 138671 41023 138699 41051
rect 138485 40961 138513 40989
rect 138547 40961 138575 40989
rect 138609 40961 138637 40989
rect 138671 40961 138699 40989
rect 138485 32147 138513 32175
rect 138547 32147 138575 32175
rect 138609 32147 138637 32175
rect 138671 32147 138699 32175
rect 138485 32085 138513 32113
rect 138547 32085 138575 32113
rect 138609 32085 138637 32113
rect 138671 32085 138699 32113
rect 138485 32023 138513 32051
rect 138547 32023 138575 32051
rect 138609 32023 138637 32051
rect 138671 32023 138699 32051
rect 138485 31961 138513 31989
rect 138547 31961 138575 31989
rect 138609 31961 138637 31989
rect 138671 31961 138699 31989
rect 138485 23147 138513 23175
rect 138547 23147 138575 23175
rect 138609 23147 138637 23175
rect 138671 23147 138699 23175
rect 138485 23085 138513 23113
rect 138547 23085 138575 23113
rect 138609 23085 138637 23113
rect 138671 23085 138699 23113
rect 138485 23023 138513 23051
rect 138547 23023 138575 23051
rect 138609 23023 138637 23051
rect 138671 23023 138699 23051
rect 138485 22961 138513 22989
rect 138547 22961 138575 22989
rect 138609 22961 138637 22989
rect 138671 22961 138699 22989
rect 138485 14147 138513 14175
rect 138547 14147 138575 14175
rect 138609 14147 138637 14175
rect 138671 14147 138699 14175
rect 138485 14085 138513 14113
rect 138547 14085 138575 14113
rect 138609 14085 138637 14113
rect 138671 14085 138699 14113
rect 138485 14023 138513 14051
rect 138547 14023 138575 14051
rect 138609 14023 138637 14051
rect 138671 14023 138699 14051
rect 138485 13961 138513 13989
rect 138547 13961 138575 13989
rect 138609 13961 138637 13989
rect 138671 13961 138699 13989
rect 138485 5147 138513 5175
rect 138547 5147 138575 5175
rect 138609 5147 138637 5175
rect 138671 5147 138699 5175
rect 138485 5085 138513 5113
rect 138547 5085 138575 5113
rect 138609 5085 138637 5113
rect 138671 5085 138699 5113
rect 138485 5023 138513 5051
rect 138547 5023 138575 5051
rect 138609 5023 138637 5051
rect 138671 5023 138699 5051
rect 138485 4961 138513 4989
rect 138547 4961 138575 4989
rect 138609 4961 138637 4989
rect 138671 4961 138699 4989
rect 138485 -588 138513 -560
rect 138547 -588 138575 -560
rect 138609 -588 138637 -560
rect 138671 -588 138699 -560
rect 138485 -650 138513 -622
rect 138547 -650 138575 -622
rect 138609 -650 138637 -622
rect 138671 -650 138699 -622
rect 138485 -712 138513 -684
rect 138547 -712 138575 -684
rect 138609 -712 138637 -684
rect 138671 -712 138699 -684
rect 138485 -774 138513 -746
rect 138547 -774 138575 -746
rect 138609 -774 138637 -746
rect 138671 -774 138699 -746
rect 145625 119147 145653 119175
rect 145687 119147 145715 119175
rect 145749 119147 145777 119175
rect 145811 119147 145839 119175
rect 145625 119085 145653 119113
rect 145687 119085 145715 119113
rect 145749 119085 145777 119113
rect 145811 119085 145839 119113
rect 145625 119023 145653 119051
rect 145687 119023 145715 119051
rect 145749 119023 145777 119051
rect 145811 119023 145839 119051
rect 145625 118961 145653 118989
rect 145687 118961 145715 118989
rect 145749 118961 145777 118989
rect 145811 118961 145839 118989
rect 145625 110147 145653 110175
rect 145687 110147 145715 110175
rect 145749 110147 145777 110175
rect 145811 110147 145839 110175
rect 145625 110085 145653 110113
rect 145687 110085 145715 110113
rect 145749 110085 145777 110113
rect 145811 110085 145839 110113
rect 145625 110023 145653 110051
rect 145687 110023 145715 110051
rect 145749 110023 145777 110051
rect 145811 110023 145839 110051
rect 145625 109961 145653 109989
rect 145687 109961 145715 109989
rect 145749 109961 145777 109989
rect 145811 109961 145839 109989
rect 145625 101147 145653 101175
rect 145687 101147 145715 101175
rect 145749 101147 145777 101175
rect 145811 101147 145839 101175
rect 145625 101085 145653 101113
rect 145687 101085 145715 101113
rect 145749 101085 145777 101113
rect 145811 101085 145839 101113
rect 145625 101023 145653 101051
rect 145687 101023 145715 101051
rect 145749 101023 145777 101051
rect 145811 101023 145839 101051
rect 145625 100961 145653 100989
rect 145687 100961 145715 100989
rect 145749 100961 145777 100989
rect 145811 100961 145839 100989
rect 145625 92147 145653 92175
rect 145687 92147 145715 92175
rect 145749 92147 145777 92175
rect 145811 92147 145839 92175
rect 145625 92085 145653 92113
rect 145687 92085 145715 92113
rect 145749 92085 145777 92113
rect 145811 92085 145839 92113
rect 145625 92023 145653 92051
rect 145687 92023 145715 92051
rect 145749 92023 145777 92051
rect 145811 92023 145839 92051
rect 145625 91961 145653 91989
rect 145687 91961 145715 91989
rect 145749 91961 145777 91989
rect 145811 91961 145839 91989
rect 145625 83147 145653 83175
rect 145687 83147 145715 83175
rect 145749 83147 145777 83175
rect 145811 83147 145839 83175
rect 145625 83085 145653 83113
rect 145687 83085 145715 83113
rect 145749 83085 145777 83113
rect 145811 83085 145839 83113
rect 145625 83023 145653 83051
rect 145687 83023 145715 83051
rect 145749 83023 145777 83051
rect 145811 83023 145839 83051
rect 145625 82961 145653 82989
rect 145687 82961 145715 82989
rect 145749 82961 145777 82989
rect 145811 82961 145839 82989
rect 145625 74147 145653 74175
rect 145687 74147 145715 74175
rect 145749 74147 145777 74175
rect 145811 74147 145839 74175
rect 145625 74085 145653 74113
rect 145687 74085 145715 74113
rect 145749 74085 145777 74113
rect 145811 74085 145839 74113
rect 145625 74023 145653 74051
rect 145687 74023 145715 74051
rect 145749 74023 145777 74051
rect 145811 74023 145839 74051
rect 145625 73961 145653 73989
rect 145687 73961 145715 73989
rect 145749 73961 145777 73989
rect 145811 73961 145839 73989
rect 145625 65147 145653 65175
rect 145687 65147 145715 65175
rect 145749 65147 145777 65175
rect 145811 65147 145839 65175
rect 145625 65085 145653 65113
rect 145687 65085 145715 65113
rect 145749 65085 145777 65113
rect 145811 65085 145839 65113
rect 145625 65023 145653 65051
rect 145687 65023 145715 65051
rect 145749 65023 145777 65051
rect 145811 65023 145839 65051
rect 145625 64961 145653 64989
rect 145687 64961 145715 64989
rect 145749 64961 145777 64989
rect 145811 64961 145839 64989
rect 145625 56147 145653 56175
rect 145687 56147 145715 56175
rect 145749 56147 145777 56175
rect 145811 56147 145839 56175
rect 145625 56085 145653 56113
rect 145687 56085 145715 56113
rect 145749 56085 145777 56113
rect 145811 56085 145839 56113
rect 145625 56023 145653 56051
rect 145687 56023 145715 56051
rect 145749 56023 145777 56051
rect 145811 56023 145839 56051
rect 145625 55961 145653 55989
rect 145687 55961 145715 55989
rect 145749 55961 145777 55989
rect 145811 55961 145839 55989
rect 145625 47147 145653 47175
rect 145687 47147 145715 47175
rect 145749 47147 145777 47175
rect 145811 47147 145839 47175
rect 145625 47085 145653 47113
rect 145687 47085 145715 47113
rect 145749 47085 145777 47113
rect 145811 47085 145839 47113
rect 145625 47023 145653 47051
rect 145687 47023 145715 47051
rect 145749 47023 145777 47051
rect 145811 47023 145839 47051
rect 145625 46961 145653 46989
rect 145687 46961 145715 46989
rect 145749 46961 145777 46989
rect 145811 46961 145839 46989
rect 145625 38147 145653 38175
rect 145687 38147 145715 38175
rect 145749 38147 145777 38175
rect 145811 38147 145839 38175
rect 145625 38085 145653 38113
rect 145687 38085 145715 38113
rect 145749 38085 145777 38113
rect 145811 38085 145839 38113
rect 145625 38023 145653 38051
rect 145687 38023 145715 38051
rect 145749 38023 145777 38051
rect 145811 38023 145839 38051
rect 145625 37961 145653 37989
rect 145687 37961 145715 37989
rect 145749 37961 145777 37989
rect 145811 37961 145839 37989
rect 145625 29147 145653 29175
rect 145687 29147 145715 29175
rect 145749 29147 145777 29175
rect 145811 29147 145839 29175
rect 145625 29085 145653 29113
rect 145687 29085 145715 29113
rect 145749 29085 145777 29113
rect 145811 29085 145839 29113
rect 145625 29023 145653 29051
rect 145687 29023 145715 29051
rect 145749 29023 145777 29051
rect 145811 29023 145839 29051
rect 145625 28961 145653 28989
rect 145687 28961 145715 28989
rect 145749 28961 145777 28989
rect 145811 28961 145839 28989
rect 145625 20147 145653 20175
rect 145687 20147 145715 20175
rect 145749 20147 145777 20175
rect 145811 20147 145839 20175
rect 145625 20085 145653 20113
rect 145687 20085 145715 20113
rect 145749 20085 145777 20113
rect 145811 20085 145839 20113
rect 145625 20023 145653 20051
rect 145687 20023 145715 20051
rect 145749 20023 145777 20051
rect 145811 20023 145839 20051
rect 145625 19961 145653 19989
rect 145687 19961 145715 19989
rect 145749 19961 145777 19989
rect 145811 19961 145839 19989
rect 145625 11147 145653 11175
rect 145687 11147 145715 11175
rect 145749 11147 145777 11175
rect 145811 11147 145839 11175
rect 145625 11085 145653 11113
rect 145687 11085 145715 11113
rect 145749 11085 145777 11113
rect 145811 11085 145839 11113
rect 145625 11023 145653 11051
rect 145687 11023 145715 11051
rect 145749 11023 145777 11051
rect 145811 11023 145839 11051
rect 145625 10961 145653 10989
rect 145687 10961 145715 10989
rect 145749 10961 145777 10989
rect 145811 10961 145839 10989
rect 145625 2147 145653 2175
rect 145687 2147 145715 2175
rect 145749 2147 145777 2175
rect 145811 2147 145839 2175
rect 145625 2085 145653 2113
rect 145687 2085 145715 2113
rect 145749 2085 145777 2113
rect 145811 2085 145839 2113
rect 145625 2023 145653 2051
rect 145687 2023 145715 2051
rect 145749 2023 145777 2051
rect 145811 2023 145839 2051
rect 145625 1961 145653 1989
rect 145687 1961 145715 1989
rect 145749 1961 145777 1989
rect 145811 1961 145839 1989
rect 145625 -108 145653 -80
rect 145687 -108 145715 -80
rect 145749 -108 145777 -80
rect 145811 -108 145839 -80
rect 145625 -170 145653 -142
rect 145687 -170 145715 -142
rect 145749 -170 145777 -142
rect 145811 -170 145839 -142
rect 145625 -232 145653 -204
rect 145687 -232 145715 -204
rect 145749 -232 145777 -204
rect 145811 -232 145839 -204
rect 145625 -294 145653 -266
rect 145687 -294 145715 -266
rect 145749 -294 145777 -266
rect 145811 -294 145839 -266
rect 147485 122147 147513 122175
rect 147547 122147 147575 122175
rect 147609 122147 147637 122175
rect 147671 122147 147699 122175
rect 147485 122085 147513 122113
rect 147547 122085 147575 122113
rect 147609 122085 147637 122113
rect 147671 122085 147699 122113
rect 147485 122023 147513 122051
rect 147547 122023 147575 122051
rect 147609 122023 147637 122051
rect 147671 122023 147699 122051
rect 147485 121961 147513 121989
rect 147547 121961 147575 121989
rect 147609 121961 147637 121989
rect 147671 121961 147699 121989
rect 147485 113147 147513 113175
rect 147547 113147 147575 113175
rect 147609 113147 147637 113175
rect 147671 113147 147699 113175
rect 147485 113085 147513 113113
rect 147547 113085 147575 113113
rect 147609 113085 147637 113113
rect 147671 113085 147699 113113
rect 147485 113023 147513 113051
rect 147547 113023 147575 113051
rect 147609 113023 147637 113051
rect 147671 113023 147699 113051
rect 147485 112961 147513 112989
rect 147547 112961 147575 112989
rect 147609 112961 147637 112989
rect 147671 112961 147699 112989
rect 147485 104147 147513 104175
rect 147547 104147 147575 104175
rect 147609 104147 147637 104175
rect 147671 104147 147699 104175
rect 147485 104085 147513 104113
rect 147547 104085 147575 104113
rect 147609 104085 147637 104113
rect 147671 104085 147699 104113
rect 147485 104023 147513 104051
rect 147547 104023 147575 104051
rect 147609 104023 147637 104051
rect 147671 104023 147699 104051
rect 147485 103961 147513 103989
rect 147547 103961 147575 103989
rect 147609 103961 147637 103989
rect 147671 103961 147699 103989
rect 147485 95147 147513 95175
rect 147547 95147 147575 95175
rect 147609 95147 147637 95175
rect 147671 95147 147699 95175
rect 147485 95085 147513 95113
rect 147547 95085 147575 95113
rect 147609 95085 147637 95113
rect 147671 95085 147699 95113
rect 147485 95023 147513 95051
rect 147547 95023 147575 95051
rect 147609 95023 147637 95051
rect 147671 95023 147699 95051
rect 147485 94961 147513 94989
rect 147547 94961 147575 94989
rect 147609 94961 147637 94989
rect 147671 94961 147699 94989
rect 147485 86147 147513 86175
rect 147547 86147 147575 86175
rect 147609 86147 147637 86175
rect 147671 86147 147699 86175
rect 147485 86085 147513 86113
rect 147547 86085 147575 86113
rect 147609 86085 147637 86113
rect 147671 86085 147699 86113
rect 147485 86023 147513 86051
rect 147547 86023 147575 86051
rect 147609 86023 147637 86051
rect 147671 86023 147699 86051
rect 147485 85961 147513 85989
rect 147547 85961 147575 85989
rect 147609 85961 147637 85989
rect 147671 85961 147699 85989
rect 147485 77147 147513 77175
rect 147547 77147 147575 77175
rect 147609 77147 147637 77175
rect 147671 77147 147699 77175
rect 147485 77085 147513 77113
rect 147547 77085 147575 77113
rect 147609 77085 147637 77113
rect 147671 77085 147699 77113
rect 147485 77023 147513 77051
rect 147547 77023 147575 77051
rect 147609 77023 147637 77051
rect 147671 77023 147699 77051
rect 147485 76961 147513 76989
rect 147547 76961 147575 76989
rect 147609 76961 147637 76989
rect 147671 76961 147699 76989
rect 147485 68147 147513 68175
rect 147547 68147 147575 68175
rect 147609 68147 147637 68175
rect 147671 68147 147699 68175
rect 147485 68085 147513 68113
rect 147547 68085 147575 68113
rect 147609 68085 147637 68113
rect 147671 68085 147699 68113
rect 147485 68023 147513 68051
rect 147547 68023 147575 68051
rect 147609 68023 147637 68051
rect 147671 68023 147699 68051
rect 147485 67961 147513 67989
rect 147547 67961 147575 67989
rect 147609 67961 147637 67989
rect 147671 67961 147699 67989
rect 147485 59147 147513 59175
rect 147547 59147 147575 59175
rect 147609 59147 147637 59175
rect 147671 59147 147699 59175
rect 147485 59085 147513 59113
rect 147547 59085 147575 59113
rect 147609 59085 147637 59113
rect 147671 59085 147699 59113
rect 147485 59023 147513 59051
rect 147547 59023 147575 59051
rect 147609 59023 147637 59051
rect 147671 59023 147699 59051
rect 147485 58961 147513 58989
rect 147547 58961 147575 58989
rect 147609 58961 147637 58989
rect 147671 58961 147699 58989
rect 147485 50147 147513 50175
rect 147547 50147 147575 50175
rect 147609 50147 147637 50175
rect 147671 50147 147699 50175
rect 147485 50085 147513 50113
rect 147547 50085 147575 50113
rect 147609 50085 147637 50113
rect 147671 50085 147699 50113
rect 147485 50023 147513 50051
rect 147547 50023 147575 50051
rect 147609 50023 147637 50051
rect 147671 50023 147699 50051
rect 147485 49961 147513 49989
rect 147547 49961 147575 49989
rect 147609 49961 147637 49989
rect 147671 49961 147699 49989
rect 147485 41147 147513 41175
rect 147547 41147 147575 41175
rect 147609 41147 147637 41175
rect 147671 41147 147699 41175
rect 147485 41085 147513 41113
rect 147547 41085 147575 41113
rect 147609 41085 147637 41113
rect 147671 41085 147699 41113
rect 147485 41023 147513 41051
rect 147547 41023 147575 41051
rect 147609 41023 147637 41051
rect 147671 41023 147699 41051
rect 147485 40961 147513 40989
rect 147547 40961 147575 40989
rect 147609 40961 147637 40989
rect 147671 40961 147699 40989
rect 147485 32147 147513 32175
rect 147547 32147 147575 32175
rect 147609 32147 147637 32175
rect 147671 32147 147699 32175
rect 147485 32085 147513 32113
rect 147547 32085 147575 32113
rect 147609 32085 147637 32113
rect 147671 32085 147699 32113
rect 147485 32023 147513 32051
rect 147547 32023 147575 32051
rect 147609 32023 147637 32051
rect 147671 32023 147699 32051
rect 147485 31961 147513 31989
rect 147547 31961 147575 31989
rect 147609 31961 147637 31989
rect 147671 31961 147699 31989
rect 147485 23147 147513 23175
rect 147547 23147 147575 23175
rect 147609 23147 147637 23175
rect 147671 23147 147699 23175
rect 147485 23085 147513 23113
rect 147547 23085 147575 23113
rect 147609 23085 147637 23113
rect 147671 23085 147699 23113
rect 147485 23023 147513 23051
rect 147547 23023 147575 23051
rect 147609 23023 147637 23051
rect 147671 23023 147699 23051
rect 147485 22961 147513 22989
rect 147547 22961 147575 22989
rect 147609 22961 147637 22989
rect 147671 22961 147699 22989
rect 147485 14147 147513 14175
rect 147547 14147 147575 14175
rect 147609 14147 147637 14175
rect 147671 14147 147699 14175
rect 147485 14085 147513 14113
rect 147547 14085 147575 14113
rect 147609 14085 147637 14113
rect 147671 14085 147699 14113
rect 147485 14023 147513 14051
rect 147547 14023 147575 14051
rect 147609 14023 147637 14051
rect 147671 14023 147699 14051
rect 147485 13961 147513 13989
rect 147547 13961 147575 13989
rect 147609 13961 147637 13989
rect 147671 13961 147699 13989
rect 147485 5147 147513 5175
rect 147547 5147 147575 5175
rect 147609 5147 147637 5175
rect 147671 5147 147699 5175
rect 147485 5085 147513 5113
rect 147547 5085 147575 5113
rect 147609 5085 147637 5113
rect 147671 5085 147699 5113
rect 147485 5023 147513 5051
rect 147547 5023 147575 5051
rect 147609 5023 147637 5051
rect 147671 5023 147699 5051
rect 147485 4961 147513 4989
rect 147547 4961 147575 4989
rect 147609 4961 147637 4989
rect 147671 4961 147699 4989
rect 147485 -588 147513 -560
rect 147547 -588 147575 -560
rect 147609 -588 147637 -560
rect 147671 -588 147699 -560
rect 147485 -650 147513 -622
rect 147547 -650 147575 -622
rect 147609 -650 147637 -622
rect 147671 -650 147699 -622
rect 147485 -712 147513 -684
rect 147547 -712 147575 -684
rect 147609 -712 147637 -684
rect 147671 -712 147699 -684
rect 147485 -774 147513 -746
rect 147547 -774 147575 -746
rect 147609 -774 147637 -746
rect 147671 -774 147699 -746
rect 154625 119147 154653 119175
rect 154687 119147 154715 119175
rect 154749 119147 154777 119175
rect 154811 119147 154839 119175
rect 154625 119085 154653 119113
rect 154687 119085 154715 119113
rect 154749 119085 154777 119113
rect 154811 119085 154839 119113
rect 154625 119023 154653 119051
rect 154687 119023 154715 119051
rect 154749 119023 154777 119051
rect 154811 119023 154839 119051
rect 154625 118961 154653 118989
rect 154687 118961 154715 118989
rect 154749 118961 154777 118989
rect 154811 118961 154839 118989
rect 154625 110147 154653 110175
rect 154687 110147 154715 110175
rect 154749 110147 154777 110175
rect 154811 110147 154839 110175
rect 154625 110085 154653 110113
rect 154687 110085 154715 110113
rect 154749 110085 154777 110113
rect 154811 110085 154839 110113
rect 154625 110023 154653 110051
rect 154687 110023 154715 110051
rect 154749 110023 154777 110051
rect 154811 110023 154839 110051
rect 154625 109961 154653 109989
rect 154687 109961 154715 109989
rect 154749 109961 154777 109989
rect 154811 109961 154839 109989
rect 154625 101147 154653 101175
rect 154687 101147 154715 101175
rect 154749 101147 154777 101175
rect 154811 101147 154839 101175
rect 154625 101085 154653 101113
rect 154687 101085 154715 101113
rect 154749 101085 154777 101113
rect 154811 101085 154839 101113
rect 154625 101023 154653 101051
rect 154687 101023 154715 101051
rect 154749 101023 154777 101051
rect 154811 101023 154839 101051
rect 154625 100961 154653 100989
rect 154687 100961 154715 100989
rect 154749 100961 154777 100989
rect 154811 100961 154839 100989
rect 154625 92147 154653 92175
rect 154687 92147 154715 92175
rect 154749 92147 154777 92175
rect 154811 92147 154839 92175
rect 154625 92085 154653 92113
rect 154687 92085 154715 92113
rect 154749 92085 154777 92113
rect 154811 92085 154839 92113
rect 154625 92023 154653 92051
rect 154687 92023 154715 92051
rect 154749 92023 154777 92051
rect 154811 92023 154839 92051
rect 154625 91961 154653 91989
rect 154687 91961 154715 91989
rect 154749 91961 154777 91989
rect 154811 91961 154839 91989
rect 154625 83147 154653 83175
rect 154687 83147 154715 83175
rect 154749 83147 154777 83175
rect 154811 83147 154839 83175
rect 154625 83085 154653 83113
rect 154687 83085 154715 83113
rect 154749 83085 154777 83113
rect 154811 83085 154839 83113
rect 154625 83023 154653 83051
rect 154687 83023 154715 83051
rect 154749 83023 154777 83051
rect 154811 83023 154839 83051
rect 154625 82961 154653 82989
rect 154687 82961 154715 82989
rect 154749 82961 154777 82989
rect 154811 82961 154839 82989
rect 154625 74147 154653 74175
rect 154687 74147 154715 74175
rect 154749 74147 154777 74175
rect 154811 74147 154839 74175
rect 154625 74085 154653 74113
rect 154687 74085 154715 74113
rect 154749 74085 154777 74113
rect 154811 74085 154839 74113
rect 154625 74023 154653 74051
rect 154687 74023 154715 74051
rect 154749 74023 154777 74051
rect 154811 74023 154839 74051
rect 154625 73961 154653 73989
rect 154687 73961 154715 73989
rect 154749 73961 154777 73989
rect 154811 73961 154839 73989
rect 154625 65147 154653 65175
rect 154687 65147 154715 65175
rect 154749 65147 154777 65175
rect 154811 65147 154839 65175
rect 154625 65085 154653 65113
rect 154687 65085 154715 65113
rect 154749 65085 154777 65113
rect 154811 65085 154839 65113
rect 154625 65023 154653 65051
rect 154687 65023 154715 65051
rect 154749 65023 154777 65051
rect 154811 65023 154839 65051
rect 154625 64961 154653 64989
rect 154687 64961 154715 64989
rect 154749 64961 154777 64989
rect 154811 64961 154839 64989
rect 154625 56147 154653 56175
rect 154687 56147 154715 56175
rect 154749 56147 154777 56175
rect 154811 56147 154839 56175
rect 154625 56085 154653 56113
rect 154687 56085 154715 56113
rect 154749 56085 154777 56113
rect 154811 56085 154839 56113
rect 154625 56023 154653 56051
rect 154687 56023 154715 56051
rect 154749 56023 154777 56051
rect 154811 56023 154839 56051
rect 154625 55961 154653 55989
rect 154687 55961 154715 55989
rect 154749 55961 154777 55989
rect 154811 55961 154839 55989
rect 154625 47147 154653 47175
rect 154687 47147 154715 47175
rect 154749 47147 154777 47175
rect 154811 47147 154839 47175
rect 154625 47085 154653 47113
rect 154687 47085 154715 47113
rect 154749 47085 154777 47113
rect 154811 47085 154839 47113
rect 154625 47023 154653 47051
rect 154687 47023 154715 47051
rect 154749 47023 154777 47051
rect 154811 47023 154839 47051
rect 154625 46961 154653 46989
rect 154687 46961 154715 46989
rect 154749 46961 154777 46989
rect 154811 46961 154839 46989
rect 154625 38147 154653 38175
rect 154687 38147 154715 38175
rect 154749 38147 154777 38175
rect 154811 38147 154839 38175
rect 154625 38085 154653 38113
rect 154687 38085 154715 38113
rect 154749 38085 154777 38113
rect 154811 38085 154839 38113
rect 154625 38023 154653 38051
rect 154687 38023 154715 38051
rect 154749 38023 154777 38051
rect 154811 38023 154839 38051
rect 154625 37961 154653 37989
rect 154687 37961 154715 37989
rect 154749 37961 154777 37989
rect 154811 37961 154839 37989
rect 154625 29147 154653 29175
rect 154687 29147 154715 29175
rect 154749 29147 154777 29175
rect 154811 29147 154839 29175
rect 154625 29085 154653 29113
rect 154687 29085 154715 29113
rect 154749 29085 154777 29113
rect 154811 29085 154839 29113
rect 154625 29023 154653 29051
rect 154687 29023 154715 29051
rect 154749 29023 154777 29051
rect 154811 29023 154839 29051
rect 154625 28961 154653 28989
rect 154687 28961 154715 28989
rect 154749 28961 154777 28989
rect 154811 28961 154839 28989
rect 154625 20147 154653 20175
rect 154687 20147 154715 20175
rect 154749 20147 154777 20175
rect 154811 20147 154839 20175
rect 154625 20085 154653 20113
rect 154687 20085 154715 20113
rect 154749 20085 154777 20113
rect 154811 20085 154839 20113
rect 154625 20023 154653 20051
rect 154687 20023 154715 20051
rect 154749 20023 154777 20051
rect 154811 20023 154839 20051
rect 154625 19961 154653 19989
rect 154687 19961 154715 19989
rect 154749 19961 154777 19989
rect 154811 19961 154839 19989
rect 154625 11147 154653 11175
rect 154687 11147 154715 11175
rect 154749 11147 154777 11175
rect 154811 11147 154839 11175
rect 154625 11085 154653 11113
rect 154687 11085 154715 11113
rect 154749 11085 154777 11113
rect 154811 11085 154839 11113
rect 154625 11023 154653 11051
rect 154687 11023 154715 11051
rect 154749 11023 154777 11051
rect 154811 11023 154839 11051
rect 154625 10961 154653 10989
rect 154687 10961 154715 10989
rect 154749 10961 154777 10989
rect 154811 10961 154839 10989
rect 154625 2147 154653 2175
rect 154687 2147 154715 2175
rect 154749 2147 154777 2175
rect 154811 2147 154839 2175
rect 154625 2085 154653 2113
rect 154687 2085 154715 2113
rect 154749 2085 154777 2113
rect 154811 2085 154839 2113
rect 154625 2023 154653 2051
rect 154687 2023 154715 2051
rect 154749 2023 154777 2051
rect 154811 2023 154839 2051
rect 154625 1961 154653 1989
rect 154687 1961 154715 1989
rect 154749 1961 154777 1989
rect 154811 1961 154839 1989
rect 154625 -108 154653 -80
rect 154687 -108 154715 -80
rect 154749 -108 154777 -80
rect 154811 -108 154839 -80
rect 154625 -170 154653 -142
rect 154687 -170 154715 -142
rect 154749 -170 154777 -142
rect 154811 -170 154839 -142
rect 154625 -232 154653 -204
rect 154687 -232 154715 -204
rect 154749 -232 154777 -204
rect 154811 -232 154839 -204
rect 154625 -294 154653 -266
rect 154687 -294 154715 -266
rect 154749 -294 154777 -266
rect 154811 -294 154839 -266
rect 156485 299058 156513 299086
rect 156547 299058 156575 299086
rect 156609 299058 156637 299086
rect 156671 299058 156699 299086
rect 156485 298996 156513 299024
rect 156547 298996 156575 299024
rect 156609 298996 156637 299024
rect 156671 298996 156699 299024
rect 156485 298934 156513 298962
rect 156547 298934 156575 298962
rect 156609 298934 156637 298962
rect 156671 298934 156699 298962
rect 156485 298872 156513 298900
rect 156547 298872 156575 298900
rect 156609 298872 156637 298900
rect 156671 298872 156699 298900
rect 156485 293147 156513 293175
rect 156547 293147 156575 293175
rect 156609 293147 156637 293175
rect 156671 293147 156699 293175
rect 156485 293085 156513 293113
rect 156547 293085 156575 293113
rect 156609 293085 156637 293113
rect 156671 293085 156699 293113
rect 156485 293023 156513 293051
rect 156547 293023 156575 293051
rect 156609 293023 156637 293051
rect 156671 293023 156699 293051
rect 156485 292961 156513 292989
rect 156547 292961 156575 292989
rect 156609 292961 156637 292989
rect 156671 292961 156699 292989
rect 156485 284147 156513 284175
rect 156547 284147 156575 284175
rect 156609 284147 156637 284175
rect 156671 284147 156699 284175
rect 156485 284085 156513 284113
rect 156547 284085 156575 284113
rect 156609 284085 156637 284113
rect 156671 284085 156699 284113
rect 156485 284023 156513 284051
rect 156547 284023 156575 284051
rect 156609 284023 156637 284051
rect 156671 284023 156699 284051
rect 156485 283961 156513 283989
rect 156547 283961 156575 283989
rect 156609 283961 156637 283989
rect 156671 283961 156699 283989
rect 156485 275147 156513 275175
rect 156547 275147 156575 275175
rect 156609 275147 156637 275175
rect 156671 275147 156699 275175
rect 156485 275085 156513 275113
rect 156547 275085 156575 275113
rect 156609 275085 156637 275113
rect 156671 275085 156699 275113
rect 156485 275023 156513 275051
rect 156547 275023 156575 275051
rect 156609 275023 156637 275051
rect 156671 275023 156699 275051
rect 156485 274961 156513 274989
rect 156547 274961 156575 274989
rect 156609 274961 156637 274989
rect 156671 274961 156699 274989
rect 156485 266147 156513 266175
rect 156547 266147 156575 266175
rect 156609 266147 156637 266175
rect 156671 266147 156699 266175
rect 156485 266085 156513 266113
rect 156547 266085 156575 266113
rect 156609 266085 156637 266113
rect 156671 266085 156699 266113
rect 156485 266023 156513 266051
rect 156547 266023 156575 266051
rect 156609 266023 156637 266051
rect 156671 266023 156699 266051
rect 156485 265961 156513 265989
rect 156547 265961 156575 265989
rect 156609 265961 156637 265989
rect 156671 265961 156699 265989
rect 156485 257147 156513 257175
rect 156547 257147 156575 257175
rect 156609 257147 156637 257175
rect 156671 257147 156699 257175
rect 156485 257085 156513 257113
rect 156547 257085 156575 257113
rect 156609 257085 156637 257113
rect 156671 257085 156699 257113
rect 156485 257023 156513 257051
rect 156547 257023 156575 257051
rect 156609 257023 156637 257051
rect 156671 257023 156699 257051
rect 156485 256961 156513 256989
rect 156547 256961 156575 256989
rect 156609 256961 156637 256989
rect 156671 256961 156699 256989
rect 156485 248147 156513 248175
rect 156547 248147 156575 248175
rect 156609 248147 156637 248175
rect 156671 248147 156699 248175
rect 156485 248085 156513 248113
rect 156547 248085 156575 248113
rect 156609 248085 156637 248113
rect 156671 248085 156699 248113
rect 156485 248023 156513 248051
rect 156547 248023 156575 248051
rect 156609 248023 156637 248051
rect 156671 248023 156699 248051
rect 156485 247961 156513 247989
rect 156547 247961 156575 247989
rect 156609 247961 156637 247989
rect 156671 247961 156699 247989
rect 156485 239147 156513 239175
rect 156547 239147 156575 239175
rect 156609 239147 156637 239175
rect 156671 239147 156699 239175
rect 156485 239085 156513 239113
rect 156547 239085 156575 239113
rect 156609 239085 156637 239113
rect 156671 239085 156699 239113
rect 156485 239023 156513 239051
rect 156547 239023 156575 239051
rect 156609 239023 156637 239051
rect 156671 239023 156699 239051
rect 156485 238961 156513 238989
rect 156547 238961 156575 238989
rect 156609 238961 156637 238989
rect 156671 238961 156699 238989
rect 156485 230147 156513 230175
rect 156547 230147 156575 230175
rect 156609 230147 156637 230175
rect 156671 230147 156699 230175
rect 156485 230085 156513 230113
rect 156547 230085 156575 230113
rect 156609 230085 156637 230113
rect 156671 230085 156699 230113
rect 156485 230023 156513 230051
rect 156547 230023 156575 230051
rect 156609 230023 156637 230051
rect 156671 230023 156699 230051
rect 156485 229961 156513 229989
rect 156547 229961 156575 229989
rect 156609 229961 156637 229989
rect 156671 229961 156699 229989
rect 156485 221147 156513 221175
rect 156547 221147 156575 221175
rect 156609 221147 156637 221175
rect 156671 221147 156699 221175
rect 156485 221085 156513 221113
rect 156547 221085 156575 221113
rect 156609 221085 156637 221113
rect 156671 221085 156699 221113
rect 156485 221023 156513 221051
rect 156547 221023 156575 221051
rect 156609 221023 156637 221051
rect 156671 221023 156699 221051
rect 156485 220961 156513 220989
rect 156547 220961 156575 220989
rect 156609 220961 156637 220989
rect 156671 220961 156699 220989
rect 156485 212147 156513 212175
rect 156547 212147 156575 212175
rect 156609 212147 156637 212175
rect 156671 212147 156699 212175
rect 156485 212085 156513 212113
rect 156547 212085 156575 212113
rect 156609 212085 156637 212113
rect 156671 212085 156699 212113
rect 156485 212023 156513 212051
rect 156547 212023 156575 212051
rect 156609 212023 156637 212051
rect 156671 212023 156699 212051
rect 156485 211961 156513 211989
rect 156547 211961 156575 211989
rect 156609 211961 156637 211989
rect 156671 211961 156699 211989
rect 156485 203147 156513 203175
rect 156547 203147 156575 203175
rect 156609 203147 156637 203175
rect 156671 203147 156699 203175
rect 156485 203085 156513 203113
rect 156547 203085 156575 203113
rect 156609 203085 156637 203113
rect 156671 203085 156699 203113
rect 156485 203023 156513 203051
rect 156547 203023 156575 203051
rect 156609 203023 156637 203051
rect 156671 203023 156699 203051
rect 156485 202961 156513 202989
rect 156547 202961 156575 202989
rect 156609 202961 156637 202989
rect 156671 202961 156699 202989
rect 156485 194147 156513 194175
rect 156547 194147 156575 194175
rect 156609 194147 156637 194175
rect 156671 194147 156699 194175
rect 156485 194085 156513 194113
rect 156547 194085 156575 194113
rect 156609 194085 156637 194113
rect 156671 194085 156699 194113
rect 156485 194023 156513 194051
rect 156547 194023 156575 194051
rect 156609 194023 156637 194051
rect 156671 194023 156699 194051
rect 156485 193961 156513 193989
rect 156547 193961 156575 193989
rect 156609 193961 156637 193989
rect 156671 193961 156699 193989
rect 156485 185147 156513 185175
rect 156547 185147 156575 185175
rect 156609 185147 156637 185175
rect 156671 185147 156699 185175
rect 156485 185085 156513 185113
rect 156547 185085 156575 185113
rect 156609 185085 156637 185113
rect 156671 185085 156699 185113
rect 156485 185023 156513 185051
rect 156547 185023 156575 185051
rect 156609 185023 156637 185051
rect 156671 185023 156699 185051
rect 156485 184961 156513 184989
rect 156547 184961 156575 184989
rect 156609 184961 156637 184989
rect 156671 184961 156699 184989
rect 156485 176147 156513 176175
rect 156547 176147 156575 176175
rect 156609 176147 156637 176175
rect 156671 176147 156699 176175
rect 156485 176085 156513 176113
rect 156547 176085 156575 176113
rect 156609 176085 156637 176113
rect 156671 176085 156699 176113
rect 156485 176023 156513 176051
rect 156547 176023 156575 176051
rect 156609 176023 156637 176051
rect 156671 176023 156699 176051
rect 156485 175961 156513 175989
rect 156547 175961 156575 175989
rect 156609 175961 156637 175989
rect 156671 175961 156699 175989
rect 156485 167147 156513 167175
rect 156547 167147 156575 167175
rect 156609 167147 156637 167175
rect 156671 167147 156699 167175
rect 156485 167085 156513 167113
rect 156547 167085 156575 167113
rect 156609 167085 156637 167113
rect 156671 167085 156699 167113
rect 156485 167023 156513 167051
rect 156547 167023 156575 167051
rect 156609 167023 156637 167051
rect 156671 167023 156699 167051
rect 156485 166961 156513 166989
rect 156547 166961 156575 166989
rect 156609 166961 156637 166989
rect 156671 166961 156699 166989
rect 156485 158147 156513 158175
rect 156547 158147 156575 158175
rect 156609 158147 156637 158175
rect 156671 158147 156699 158175
rect 156485 158085 156513 158113
rect 156547 158085 156575 158113
rect 156609 158085 156637 158113
rect 156671 158085 156699 158113
rect 156485 158023 156513 158051
rect 156547 158023 156575 158051
rect 156609 158023 156637 158051
rect 156671 158023 156699 158051
rect 156485 157961 156513 157989
rect 156547 157961 156575 157989
rect 156609 157961 156637 157989
rect 156671 157961 156699 157989
rect 156485 149147 156513 149175
rect 156547 149147 156575 149175
rect 156609 149147 156637 149175
rect 156671 149147 156699 149175
rect 156485 149085 156513 149113
rect 156547 149085 156575 149113
rect 156609 149085 156637 149113
rect 156671 149085 156699 149113
rect 156485 149023 156513 149051
rect 156547 149023 156575 149051
rect 156609 149023 156637 149051
rect 156671 149023 156699 149051
rect 156485 148961 156513 148989
rect 156547 148961 156575 148989
rect 156609 148961 156637 148989
rect 156671 148961 156699 148989
rect 156485 140147 156513 140175
rect 156547 140147 156575 140175
rect 156609 140147 156637 140175
rect 156671 140147 156699 140175
rect 156485 140085 156513 140113
rect 156547 140085 156575 140113
rect 156609 140085 156637 140113
rect 156671 140085 156699 140113
rect 156485 140023 156513 140051
rect 156547 140023 156575 140051
rect 156609 140023 156637 140051
rect 156671 140023 156699 140051
rect 156485 139961 156513 139989
rect 156547 139961 156575 139989
rect 156609 139961 156637 139989
rect 156671 139961 156699 139989
rect 156485 131147 156513 131175
rect 156547 131147 156575 131175
rect 156609 131147 156637 131175
rect 156671 131147 156699 131175
rect 156485 131085 156513 131113
rect 156547 131085 156575 131113
rect 156609 131085 156637 131113
rect 156671 131085 156699 131113
rect 156485 131023 156513 131051
rect 156547 131023 156575 131051
rect 156609 131023 156637 131051
rect 156671 131023 156699 131051
rect 156485 130961 156513 130989
rect 156547 130961 156575 130989
rect 156609 130961 156637 130989
rect 156671 130961 156699 130989
rect 156485 122147 156513 122175
rect 156547 122147 156575 122175
rect 156609 122147 156637 122175
rect 156671 122147 156699 122175
rect 156485 122085 156513 122113
rect 156547 122085 156575 122113
rect 156609 122085 156637 122113
rect 156671 122085 156699 122113
rect 156485 122023 156513 122051
rect 156547 122023 156575 122051
rect 156609 122023 156637 122051
rect 156671 122023 156699 122051
rect 156485 121961 156513 121989
rect 156547 121961 156575 121989
rect 156609 121961 156637 121989
rect 156671 121961 156699 121989
rect 156485 113147 156513 113175
rect 156547 113147 156575 113175
rect 156609 113147 156637 113175
rect 156671 113147 156699 113175
rect 156485 113085 156513 113113
rect 156547 113085 156575 113113
rect 156609 113085 156637 113113
rect 156671 113085 156699 113113
rect 156485 113023 156513 113051
rect 156547 113023 156575 113051
rect 156609 113023 156637 113051
rect 156671 113023 156699 113051
rect 156485 112961 156513 112989
rect 156547 112961 156575 112989
rect 156609 112961 156637 112989
rect 156671 112961 156699 112989
rect 156485 104147 156513 104175
rect 156547 104147 156575 104175
rect 156609 104147 156637 104175
rect 156671 104147 156699 104175
rect 156485 104085 156513 104113
rect 156547 104085 156575 104113
rect 156609 104085 156637 104113
rect 156671 104085 156699 104113
rect 156485 104023 156513 104051
rect 156547 104023 156575 104051
rect 156609 104023 156637 104051
rect 156671 104023 156699 104051
rect 156485 103961 156513 103989
rect 156547 103961 156575 103989
rect 156609 103961 156637 103989
rect 156671 103961 156699 103989
rect 156485 95147 156513 95175
rect 156547 95147 156575 95175
rect 156609 95147 156637 95175
rect 156671 95147 156699 95175
rect 156485 95085 156513 95113
rect 156547 95085 156575 95113
rect 156609 95085 156637 95113
rect 156671 95085 156699 95113
rect 156485 95023 156513 95051
rect 156547 95023 156575 95051
rect 156609 95023 156637 95051
rect 156671 95023 156699 95051
rect 156485 94961 156513 94989
rect 156547 94961 156575 94989
rect 156609 94961 156637 94989
rect 156671 94961 156699 94989
rect 156485 86147 156513 86175
rect 156547 86147 156575 86175
rect 156609 86147 156637 86175
rect 156671 86147 156699 86175
rect 156485 86085 156513 86113
rect 156547 86085 156575 86113
rect 156609 86085 156637 86113
rect 156671 86085 156699 86113
rect 156485 86023 156513 86051
rect 156547 86023 156575 86051
rect 156609 86023 156637 86051
rect 156671 86023 156699 86051
rect 156485 85961 156513 85989
rect 156547 85961 156575 85989
rect 156609 85961 156637 85989
rect 156671 85961 156699 85989
rect 156485 77147 156513 77175
rect 156547 77147 156575 77175
rect 156609 77147 156637 77175
rect 156671 77147 156699 77175
rect 156485 77085 156513 77113
rect 156547 77085 156575 77113
rect 156609 77085 156637 77113
rect 156671 77085 156699 77113
rect 156485 77023 156513 77051
rect 156547 77023 156575 77051
rect 156609 77023 156637 77051
rect 156671 77023 156699 77051
rect 156485 76961 156513 76989
rect 156547 76961 156575 76989
rect 156609 76961 156637 76989
rect 156671 76961 156699 76989
rect 156485 68147 156513 68175
rect 156547 68147 156575 68175
rect 156609 68147 156637 68175
rect 156671 68147 156699 68175
rect 156485 68085 156513 68113
rect 156547 68085 156575 68113
rect 156609 68085 156637 68113
rect 156671 68085 156699 68113
rect 156485 68023 156513 68051
rect 156547 68023 156575 68051
rect 156609 68023 156637 68051
rect 156671 68023 156699 68051
rect 156485 67961 156513 67989
rect 156547 67961 156575 67989
rect 156609 67961 156637 67989
rect 156671 67961 156699 67989
rect 156485 59147 156513 59175
rect 156547 59147 156575 59175
rect 156609 59147 156637 59175
rect 156671 59147 156699 59175
rect 156485 59085 156513 59113
rect 156547 59085 156575 59113
rect 156609 59085 156637 59113
rect 156671 59085 156699 59113
rect 156485 59023 156513 59051
rect 156547 59023 156575 59051
rect 156609 59023 156637 59051
rect 156671 59023 156699 59051
rect 156485 58961 156513 58989
rect 156547 58961 156575 58989
rect 156609 58961 156637 58989
rect 156671 58961 156699 58989
rect 156485 50147 156513 50175
rect 156547 50147 156575 50175
rect 156609 50147 156637 50175
rect 156671 50147 156699 50175
rect 156485 50085 156513 50113
rect 156547 50085 156575 50113
rect 156609 50085 156637 50113
rect 156671 50085 156699 50113
rect 156485 50023 156513 50051
rect 156547 50023 156575 50051
rect 156609 50023 156637 50051
rect 156671 50023 156699 50051
rect 156485 49961 156513 49989
rect 156547 49961 156575 49989
rect 156609 49961 156637 49989
rect 156671 49961 156699 49989
rect 156485 41147 156513 41175
rect 156547 41147 156575 41175
rect 156609 41147 156637 41175
rect 156671 41147 156699 41175
rect 156485 41085 156513 41113
rect 156547 41085 156575 41113
rect 156609 41085 156637 41113
rect 156671 41085 156699 41113
rect 156485 41023 156513 41051
rect 156547 41023 156575 41051
rect 156609 41023 156637 41051
rect 156671 41023 156699 41051
rect 156485 40961 156513 40989
rect 156547 40961 156575 40989
rect 156609 40961 156637 40989
rect 156671 40961 156699 40989
rect 156485 32147 156513 32175
rect 156547 32147 156575 32175
rect 156609 32147 156637 32175
rect 156671 32147 156699 32175
rect 156485 32085 156513 32113
rect 156547 32085 156575 32113
rect 156609 32085 156637 32113
rect 156671 32085 156699 32113
rect 156485 32023 156513 32051
rect 156547 32023 156575 32051
rect 156609 32023 156637 32051
rect 156671 32023 156699 32051
rect 156485 31961 156513 31989
rect 156547 31961 156575 31989
rect 156609 31961 156637 31989
rect 156671 31961 156699 31989
rect 156485 23147 156513 23175
rect 156547 23147 156575 23175
rect 156609 23147 156637 23175
rect 156671 23147 156699 23175
rect 156485 23085 156513 23113
rect 156547 23085 156575 23113
rect 156609 23085 156637 23113
rect 156671 23085 156699 23113
rect 156485 23023 156513 23051
rect 156547 23023 156575 23051
rect 156609 23023 156637 23051
rect 156671 23023 156699 23051
rect 156485 22961 156513 22989
rect 156547 22961 156575 22989
rect 156609 22961 156637 22989
rect 156671 22961 156699 22989
rect 156485 14147 156513 14175
rect 156547 14147 156575 14175
rect 156609 14147 156637 14175
rect 156671 14147 156699 14175
rect 156485 14085 156513 14113
rect 156547 14085 156575 14113
rect 156609 14085 156637 14113
rect 156671 14085 156699 14113
rect 156485 14023 156513 14051
rect 156547 14023 156575 14051
rect 156609 14023 156637 14051
rect 156671 14023 156699 14051
rect 156485 13961 156513 13989
rect 156547 13961 156575 13989
rect 156609 13961 156637 13989
rect 156671 13961 156699 13989
rect 156485 5147 156513 5175
rect 156547 5147 156575 5175
rect 156609 5147 156637 5175
rect 156671 5147 156699 5175
rect 156485 5085 156513 5113
rect 156547 5085 156575 5113
rect 156609 5085 156637 5113
rect 156671 5085 156699 5113
rect 156485 5023 156513 5051
rect 156547 5023 156575 5051
rect 156609 5023 156637 5051
rect 156671 5023 156699 5051
rect 156485 4961 156513 4989
rect 156547 4961 156575 4989
rect 156609 4961 156637 4989
rect 156671 4961 156699 4989
rect 156485 -588 156513 -560
rect 156547 -588 156575 -560
rect 156609 -588 156637 -560
rect 156671 -588 156699 -560
rect 156485 -650 156513 -622
rect 156547 -650 156575 -622
rect 156609 -650 156637 -622
rect 156671 -650 156699 -622
rect 156485 -712 156513 -684
rect 156547 -712 156575 -684
rect 156609 -712 156637 -684
rect 156671 -712 156699 -684
rect 156485 -774 156513 -746
rect 156547 -774 156575 -746
rect 156609 -774 156637 -746
rect 156671 -774 156699 -746
rect 163625 298578 163653 298606
rect 163687 298578 163715 298606
rect 163749 298578 163777 298606
rect 163811 298578 163839 298606
rect 163625 298516 163653 298544
rect 163687 298516 163715 298544
rect 163749 298516 163777 298544
rect 163811 298516 163839 298544
rect 163625 298454 163653 298482
rect 163687 298454 163715 298482
rect 163749 298454 163777 298482
rect 163811 298454 163839 298482
rect 163625 298392 163653 298420
rect 163687 298392 163715 298420
rect 163749 298392 163777 298420
rect 163811 298392 163839 298420
rect 163625 290147 163653 290175
rect 163687 290147 163715 290175
rect 163749 290147 163777 290175
rect 163811 290147 163839 290175
rect 163625 290085 163653 290113
rect 163687 290085 163715 290113
rect 163749 290085 163777 290113
rect 163811 290085 163839 290113
rect 163625 290023 163653 290051
rect 163687 290023 163715 290051
rect 163749 290023 163777 290051
rect 163811 290023 163839 290051
rect 163625 289961 163653 289989
rect 163687 289961 163715 289989
rect 163749 289961 163777 289989
rect 163811 289961 163839 289989
rect 163625 281147 163653 281175
rect 163687 281147 163715 281175
rect 163749 281147 163777 281175
rect 163811 281147 163839 281175
rect 163625 281085 163653 281113
rect 163687 281085 163715 281113
rect 163749 281085 163777 281113
rect 163811 281085 163839 281113
rect 163625 281023 163653 281051
rect 163687 281023 163715 281051
rect 163749 281023 163777 281051
rect 163811 281023 163839 281051
rect 163625 280961 163653 280989
rect 163687 280961 163715 280989
rect 163749 280961 163777 280989
rect 163811 280961 163839 280989
rect 163625 272147 163653 272175
rect 163687 272147 163715 272175
rect 163749 272147 163777 272175
rect 163811 272147 163839 272175
rect 163625 272085 163653 272113
rect 163687 272085 163715 272113
rect 163749 272085 163777 272113
rect 163811 272085 163839 272113
rect 163625 272023 163653 272051
rect 163687 272023 163715 272051
rect 163749 272023 163777 272051
rect 163811 272023 163839 272051
rect 163625 271961 163653 271989
rect 163687 271961 163715 271989
rect 163749 271961 163777 271989
rect 163811 271961 163839 271989
rect 163625 263147 163653 263175
rect 163687 263147 163715 263175
rect 163749 263147 163777 263175
rect 163811 263147 163839 263175
rect 163625 263085 163653 263113
rect 163687 263085 163715 263113
rect 163749 263085 163777 263113
rect 163811 263085 163839 263113
rect 163625 263023 163653 263051
rect 163687 263023 163715 263051
rect 163749 263023 163777 263051
rect 163811 263023 163839 263051
rect 163625 262961 163653 262989
rect 163687 262961 163715 262989
rect 163749 262961 163777 262989
rect 163811 262961 163839 262989
rect 163625 254147 163653 254175
rect 163687 254147 163715 254175
rect 163749 254147 163777 254175
rect 163811 254147 163839 254175
rect 163625 254085 163653 254113
rect 163687 254085 163715 254113
rect 163749 254085 163777 254113
rect 163811 254085 163839 254113
rect 163625 254023 163653 254051
rect 163687 254023 163715 254051
rect 163749 254023 163777 254051
rect 163811 254023 163839 254051
rect 163625 253961 163653 253989
rect 163687 253961 163715 253989
rect 163749 253961 163777 253989
rect 163811 253961 163839 253989
rect 163625 245147 163653 245175
rect 163687 245147 163715 245175
rect 163749 245147 163777 245175
rect 163811 245147 163839 245175
rect 163625 245085 163653 245113
rect 163687 245085 163715 245113
rect 163749 245085 163777 245113
rect 163811 245085 163839 245113
rect 163625 245023 163653 245051
rect 163687 245023 163715 245051
rect 163749 245023 163777 245051
rect 163811 245023 163839 245051
rect 163625 244961 163653 244989
rect 163687 244961 163715 244989
rect 163749 244961 163777 244989
rect 163811 244961 163839 244989
rect 163625 236147 163653 236175
rect 163687 236147 163715 236175
rect 163749 236147 163777 236175
rect 163811 236147 163839 236175
rect 163625 236085 163653 236113
rect 163687 236085 163715 236113
rect 163749 236085 163777 236113
rect 163811 236085 163839 236113
rect 163625 236023 163653 236051
rect 163687 236023 163715 236051
rect 163749 236023 163777 236051
rect 163811 236023 163839 236051
rect 163625 235961 163653 235989
rect 163687 235961 163715 235989
rect 163749 235961 163777 235989
rect 163811 235961 163839 235989
rect 163625 227147 163653 227175
rect 163687 227147 163715 227175
rect 163749 227147 163777 227175
rect 163811 227147 163839 227175
rect 163625 227085 163653 227113
rect 163687 227085 163715 227113
rect 163749 227085 163777 227113
rect 163811 227085 163839 227113
rect 163625 227023 163653 227051
rect 163687 227023 163715 227051
rect 163749 227023 163777 227051
rect 163811 227023 163839 227051
rect 163625 226961 163653 226989
rect 163687 226961 163715 226989
rect 163749 226961 163777 226989
rect 163811 226961 163839 226989
rect 163625 218147 163653 218175
rect 163687 218147 163715 218175
rect 163749 218147 163777 218175
rect 163811 218147 163839 218175
rect 163625 218085 163653 218113
rect 163687 218085 163715 218113
rect 163749 218085 163777 218113
rect 163811 218085 163839 218113
rect 163625 218023 163653 218051
rect 163687 218023 163715 218051
rect 163749 218023 163777 218051
rect 163811 218023 163839 218051
rect 163625 217961 163653 217989
rect 163687 217961 163715 217989
rect 163749 217961 163777 217989
rect 163811 217961 163839 217989
rect 163625 209147 163653 209175
rect 163687 209147 163715 209175
rect 163749 209147 163777 209175
rect 163811 209147 163839 209175
rect 163625 209085 163653 209113
rect 163687 209085 163715 209113
rect 163749 209085 163777 209113
rect 163811 209085 163839 209113
rect 163625 209023 163653 209051
rect 163687 209023 163715 209051
rect 163749 209023 163777 209051
rect 163811 209023 163839 209051
rect 163625 208961 163653 208989
rect 163687 208961 163715 208989
rect 163749 208961 163777 208989
rect 163811 208961 163839 208989
rect 163625 200147 163653 200175
rect 163687 200147 163715 200175
rect 163749 200147 163777 200175
rect 163811 200147 163839 200175
rect 163625 200085 163653 200113
rect 163687 200085 163715 200113
rect 163749 200085 163777 200113
rect 163811 200085 163839 200113
rect 163625 200023 163653 200051
rect 163687 200023 163715 200051
rect 163749 200023 163777 200051
rect 163811 200023 163839 200051
rect 163625 199961 163653 199989
rect 163687 199961 163715 199989
rect 163749 199961 163777 199989
rect 163811 199961 163839 199989
rect 163625 191147 163653 191175
rect 163687 191147 163715 191175
rect 163749 191147 163777 191175
rect 163811 191147 163839 191175
rect 163625 191085 163653 191113
rect 163687 191085 163715 191113
rect 163749 191085 163777 191113
rect 163811 191085 163839 191113
rect 163625 191023 163653 191051
rect 163687 191023 163715 191051
rect 163749 191023 163777 191051
rect 163811 191023 163839 191051
rect 163625 190961 163653 190989
rect 163687 190961 163715 190989
rect 163749 190961 163777 190989
rect 163811 190961 163839 190989
rect 163625 182147 163653 182175
rect 163687 182147 163715 182175
rect 163749 182147 163777 182175
rect 163811 182147 163839 182175
rect 163625 182085 163653 182113
rect 163687 182085 163715 182113
rect 163749 182085 163777 182113
rect 163811 182085 163839 182113
rect 163625 182023 163653 182051
rect 163687 182023 163715 182051
rect 163749 182023 163777 182051
rect 163811 182023 163839 182051
rect 163625 181961 163653 181989
rect 163687 181961 163715 181989
rect 163749 181961 163777 181989
rect 163811 181961 163839 181989
rect 163625 173147 163653 173175
rect 163687 173147 163715 173175
rect 163749 173147 163777 173175
rect 163811 173147 163839 173175
rect 163625 173085 163653 173113
rect 163687 173085 163715 173113
rect 163749 173085 163777 173113
rect 163811 173085 163839 173113
rect 163625 173023 163653 173051
rect 163687 173023 163715 173051
rect 163749 173023 163777 173051
rect 163811 173023 163839 173051
rect 163625 172961 163653 172989
rect 163687 172961 163715 172989
rect 163749 172961 163777 172989
rect 163811 172961 163839 172989
rect 163625 164147 163653 164175
rect 163687 164147 163715 164175
rect 163749 164147 163777 164175
rect 163811 164147 163839 164175
rect 163625 164085 163653 164113
rect 163687 164085 163715 164113
rect 163749 164085 163777 164113
rect 163811 164085 163839 164113
rect 163625 164023 163653 164051
rect 163687 164023 163715 164051
rect 163749 164023 163777 164051
rect 163811 164023 163839 164051
rect 163625 163961 163653 163989
rect 163687 163961 163715 163989
rect 163749 163961 163777 163989
rect 163811 163961 163839 163989
rect 163625 155147 163653 155175
rect 163687 155147 163715 155175
rect 163749 155147 163777 155175
rect 163811 155147 163839 155175
rect 163625 155085 163653 155113
rect 163687 155085 163715 155113
rect 163749 155085 163777 155113
rect 163811 155085 163839 155113
rect 163625 155023 163653 155051
rect 163687 155023 163715 155051
rect 163749 155023 163777 155051
rect 163811 155023 163839 155051
rect 163625 154961 163653 154989
rect 163687 154961 163715 154989
rect 163749 154961 163777 154989
rect 163811 154961 163839 154989
rect 163625 146147 163653 146175
rect 163687 146147 163715 146175
rect 163749 146147 163777 146175
rect 163811 146147 163839 146175
rect 163625 146085 163653 146113
rect 163687 146085 163715 146113
rect 163749 146085 163777 146113
rect 163811 146085 163839 146113
rect 163625 146023 163653 146051
rect 163687 146023 163715 146051
rect 163749 146023 163777 146051
rect 163811 146023 163839 146051
rect 163625 145961 163653 145989
rect 163687 145961 163715 145989
rect 163749 145961 163777 145989
rect 163811 145961 163839 145989
rect 163625 137147 163653 137175
rect 163687 137147 163715 137175
rect 163749 137147 163777 137175
rect 163811 137147 163839 137175
rect 163625 137085 163653 137113
rect 163687 137085 163715 137113
rect 163749 137085 163777 137113
rect 163811 137085 163839 137113
rect 163625 137023 163653 137051
rect 163687 137023 163715 137051
rect 163749 137023 163777 137051
rect 163811 137023 163839 137051
rect 163625 136961 163653 136989
rect 163687 136961 163715 136989
rect 163749 136961 163777 136989
rect 163811 136961 163839 136989
rect 163625 128147 163653 128175
rect 163687 128147 163715 128175
rect 163749 128147 163777 128175
rect 163811 128147 163839 128175
rect 163625 128085 163653 128113
rect 163687 128085 163715 128113
rect 163749 128085 163777 128113
rect 163811 128085 163839 128113
rect 163625 128023 163653 128051
rect 163687 128023 163715 128051
rect 163749 128023 163777 128051
rect 163811 128023 163839 128051
rect 163625 127961 163653 127989
rect 163687 127961 163715 127989
rect 163749 127961 163777 127989
rect 163811 127961 163839 127989
rect 163625 119147 163653 119175
rect 163687 119147 163715 119175
rect 163749 119147 163777 119175
rect 163811 119147 163839 119175
rect 163625 119085 163653 119113
rect 163687 119085 163715 119113
rect 163749 119085 163777 119113
rect 163811 119085 163839 119113
rect 163625 119023 163653 119051
rect 163687 119023 163715 119051
rect 163749 119023 163777 119051
rect 163811 119023 163839 119051
rect 163625 118961 163653 118989
rect 163687 118961 163715 118989
rect 163749 118961 163777 118989
rect 163811 118961 163839 118989
rect 163625 110147 163653 110175
rect 163687 110147 163715 110175
rect 163749 110147 163777 110175
rect 163811 110147 163839 110175
rect 163625 110085 163653 110113
rect 163687 110085 163715 110113
rect 163749 110085 163777 110113
rect 163811 110085 163839 110113
rect 163625 110023 163653 110051
rect 163687 110023 163715 110051
rect 163749 110023 163777 110051
rect 163811 110023 163839 110051
rect 163625 109961 163653 109989
rect 163687 109961 163715 109989
rect 163749 109961 163777 109989
rect 163811 109961 163839 109989
rect 163625 101147 163653 101175
rect 163687 101147 163715 101175
rect 163749 101147 163777 101175
rect 163811 101147 163839 101175
rect 163625 101085 163653 101113
rect 163687 101085 163715 101113
rect 163749 101085 163777 101113
rect 163811 101085 163839 101113
rect 163625 101023 163653 101051
rect 163687 101023 163715 101051
rect 163749 101023 163777 101051
rect 163811 101023 163839 101051
rect 163625 100961 163653 100989
rect 163687 100961 163715 100989
rect 163749 100961 163777 100989
rect 163811 100961 163839 100989
rect 163625 92147 163653 92175
rect 163687 92147 163715 92175
rect 163749 92147 163777 92175
rect 163811 92147 163839 92175
rect 163625 92085 163653 92113
rect 163687 92085 163715 92113
rect 163749 92085 163777 92113
rect 163811 92085 163839 92113
rect 163625 92023 163653 92051
rect 163687 92023 163715 92051
rect 163749 92023 163777 92051
rect 163811 92023 163839 92051
rect 163625 91961 163653 91989
rect 163687 91961 163715 91989
rect 163749 91961 163777 91989
rect 163811 91961 163839 91989
rect 163625 83147 163653 83175
rect 163687 83147 163715 83175
rect 163749 83147 163777 83175
rect 163811 83147 163839 83175
rect 163625 83085 163653 83113
rect 163687 83085 163715 83113
rect 163749 83085 163777 83113
rect 163811 83085 163839 83113
rect 163625 83023 163653 83051
rect 163687 83023 163715 83051
rect 163749 83023 163777 83051
rect 163811 83023 163839 83051
rect 163625 82961 163653 82989
rect 163687 82961 163715 82989
rect 163749 82961 163777 82989
rect 163811 82961 163839 82989
rect 163625 74147 163653 74175
rect 163687 74147 163715 74175
rect 163749 74147 163777 74175
rect 163811 74147 163839 74175
rect 163625 74085 163653 74113
rect 163687 74085 163715 74113
rect 163749 74085 163777 74113
rect 163811 74085 163839 74113
rect 163625 74023 163653 74051
rect 163687 74023 163715 74051
rect 163749 74023 163777 74051
rect 163811 74023 163839 74051
rect 163625 73961 163653 73989
rect 163687 73961 163715 73989
rect 163749 73961 163777 73989
rect 163811 73961 163839 73989
rect 163625 65147 163653 65175
rect 163687 65147 163715 65175
rect 163749 65147 163777 65175
rect 163811 65147 163839 65175
rect 163625 65085 163653 65113
rect 163687 65085 163715 65113
rect 163749 65085 163777 65113
rect 163811 65085 163839 65113
rect 163625 65023 163653 65051
rect 163687 65023 163715 65051
rect 163749 65023 163777 65051
rect 163811 65023 163839 65051
rect 163625 64961 163653 64989
rect 163687 64961 163715 64989
rect 163749 64961 163777 64989
rect 163811 64961 163839 64989
rect 163625 56147 163653 56175
rect 163687 56147 163715 56175
rect 163749 56147 163777 56175
rect 163811 56147 163839 56175
rect 163625 56085 163653 56113
rect 163687 56085 163715 56113
rect 163749 56085 163777 56113
rect 163811 56085 163839 56113
rect 163625 56023 163653 56051
rect 163687 56023 163715 56051
rect 163749 56023 163777 56051
rect 163811 56023 163839 56051
rect 163625 55961 163653 55989
rect 163687 55961 163715 55989
rect 163749 55961 163777 55989
rect 163811 55961 163839 55989
rect 163625 47147 163653 47175
rect 163687 47147 163715 47175
rect 163749 47147 163777 47175
rect 163811 47147 163839 47175
rect 163625 47085 163653 47113
rect 163687 47085 163715 47113
rect 163749 47085 163777 47113
rect 163811 47085 163839 47113
rect 163625 47023 163653 47051
rect 163687 47023 163715 47051
rect 163749 47023 163777 47051
rect 163811 47023 163839 47051
rect 163625 46961 163653 46989
rect 163687 46961 163715 46989
rect 163749 46961 163777 46989
rect 163811 46961 163839 46989
rect 163625 38147 163653 38175
rect 163687 38147 163715 38175
rect 163749 38147 163777 38175
rect 163811 38147 163839 38175
rect 163625 38085 163653 38113
rect 163687 38085 163715 38113
rect 163749 38085 163777 38113
rect 163811 38085 163839 38113
rect 163625 38023 163653 38051
rect 163687 38023 163715 38051
rect 163749 38023 163777 38051
rect 163811 38023 163839 38051
rect 163625 37961 163653 37989
rect 163687 37961 163715 37989
rect 163749 37961 163777 37989
rect 163811 37961 163839 37989
rect 163625 29147 163653 29175
rect 163687 29147 163715 29175
rect 163749 29147 163777 29175
rect 163811 29147 163839 29175
rect 163625 29085 163653 29113
rect 163687 29085 163715 29113
rect 163749 29085 163777 29113
rect 163811 29085 163839 29113
rect 163625 29023 163653 29051
rect 163687 29023 163715 29051
rect 163749 29023 163777 29051
rect 163811 29023 163839 29051
rect 163625 28961 163653 28989
rect 163687 28961 163715 28989
rect 163749 28961 163777 28989
rect 163811 28961 163839 28989
rect 163625 20147 163653 20175
rect 163687 20147 163715 20175
rect 163749 20147 163777 20175
rect 163811 20147 163839 20175
rect 163625 20085 163653 20113
rect 163687 20085 163715 20113
rect 163749 20085 163777 20113
rect 163811 20085 163839 20113
rect 163625 20023 163653 20051
rect 163687 20023 163715 20051
rect 163749 20023 163777 20051
rect 163811 20023 163839 20051
rect 163625 19961 163653 19989
rect 163687 19961 163715 19989
rect 163749 19961 163777 19989
rect 163811 19961 163839 19989
rect 163625 11147 163653 11175
rect 163687 11147 163715 11175
rect 163749 11147 163777 11175
rect 163811 11147 163839 11175
rect 163625 11085 163653 11113
rect 163687 11085 163715 11113
rect 163749 11085 163777 11113
rect 163811 11085 163839 11113
rect 163625 11023 163653 11051
rect 163687 11023 163715 11051
rect 163749 11023 163777 11051
rect 163811 11023 163839 11051
rect 163625 10961 163653 10989
rect 163687 10961 163715 10989
rect 163749 10961 163777 10989
rect 163811 10961 163839 10989
rect 163625 2147 163653 2175
rect 163687 2147 163715 2175
rect 163749 2147 163777 2175
rect 163811 2147 163839 2175
rect 163625 2085 163653 2113
rect 163687 2085 163715 2113
rect 163749 2085 163777 2113
rect 163811 2085 163839 2113
rect 163625 2023 163653 2051
rect 163687 2023 163715 2051
rect 163749 2023 163777 2051
rect 163811 2023 163839 2051
rect 163625 1961 163653 1989
rect 163687 1961 163715 1989
rect 163749 1961 163777 1989
rect 163811 1961 163839 1989
rect 163625 -108 163653 -80
rect 163687 -108 163715 -80
rect 163749 -108 163777 -80
rect 163811 -108 163839 -80
rect 163625 -170 163653 -142
rect 163687 -170 163715 -142
rect 163749 -170 163777 -142
rect 163811 -170 163839 -142
rect 163625 -232 163653 -204
rect 163687 -232 163715 -204
rect 163749 -232 163777 -204
rect 163811 -232 163839 -204
rect 163625 -294 163653 -266
rect 163687 -294 163715 -266
rect 163749 -294 163777 -266
rect 163811 -294 163839 -266
rect 165485 299058 165513 299086
rect 165547 299058 165575 299086
rect 165609 299058 165637 299086
rect 165671 299058 165699 299086
rect 165485 298996 165513 299024
rect 165547 298996 165575 299024
rect 165609 298996 165637 299024
rect 165671 298996 165699 299024
rect 165485 298934 165513 298962
rect 165547 298934 165575 298962
rect 165609 298934 165637 298962
rect 165671 298934 165699 298962
rect 165485 298872 165513 298900
rect 165547 298872 165575 298900
rect 165609 298872 165637 298900
rect 165671 298872 165699 298900
rect 165485 293147 165513 293175
rect 165547 293147 165575 293175
rect 165609 293147 165637 293175
rect 165671 293147 165699 293175
rect 165485 293085 165513 293113
rect 165547 293085 165575 293113
rect 165609 293085 165637 293113
rect 165671 293085 165699 293113
rect 165485 293023 165513 293051
rect 165547 293023 165575 293051
rect 165609 293023 165637 293051
rect 165671 293023 165699 293051
rect 165485 292961 165513 292989
rect 165547 292961 165575 292989
rect 165609 292961 165637 292989
rect 165671 292961 165699 292989
rect 165485 284147 165513 284175
rect 165547 284147 165575 284175
rect 165609 284147 165637 284175
rect 165671 284147 165699 284175
rect 165485 284085 165513 284113
rect 165547 284085 165575 284113
rect 165609 284085 165637 284113
rect 165671 284085 165699 284113
rect 165485 284023 165513 284051
rect 165547 284023 165575 284051
rect 165609 284023 165637 284051
rect 165671 284023 165699 284051
rect 165485 283961 165513 283989
rect 165547 283961 165575 283989
rect 165609 283961 165637 283989
rect 165671 283961 165699 283989
rect 165485 275147 165513 275175
rect 165547 275147 165575 275175
rect 165609 275147 165637 275175
rect 165671 275147 165699 275175
rect 165485 275085 165513 275113
rect 165547 275085 165575 275113
rect 165609 275085 165637 275113
rect 165671 275085 165699 275113
rect 165485 275023 165513 275051
rect 165547 275023 165575 275051
rect 165609 275023 165637 275051
rect 165671 275023 165699 275051
rect 165485 274961 165513 274989
rect 165547 274961 165575 274989
rect 165609 274961 165637 274989
rect 165671 274961 165699 274989
rect 165485 266147 165513 266175
rect 165547 266147 165575 266175
rect 165609 266147 165637 266175
rect 165671 266147 165699 266175
rect 165485 266085 165513 266113
rect 165547 266085 165575 266113
rect 165609 266085 165637 266113
rect 165671 266085 165699 266113
rect 165485 266023 165513 266051
rect 165547 266023 165575 266051
rect 165609 266023 165637 266051
rect 165671 266023 165699 266051
rect 165485 265961 165513 265989
rect 165547 265961 165575 265989
rect 165609 265961 165637 265989
rect 165671 265961 165699 265989
rect 165485 257147 165513 257175
rect 165547 257147 165575 257175
rect 165609 257147 165637 257175
rect 165671 257147 165699 257175
rect 165485 257085 165513 257113
rect 165547 257085 165575 257113
rect 165609 257085 165637 257113
rect 165671 257085 165699 257113
rect 165485 257023 165513 257051
rect 165547 257023 165575 257051
rect 165609 257023 165637 257051
rect 165671 257023 165699 257051
rect 165485 256961 165513 256989
rect 165547 256961 165575 256989
rect 165609 256961 165637 256989
rect 165671 256961 165699 256989
rect 165485 248147 165513 248175
rect 165547 248147 165575 248175
rect 165609 248147 165637 248175
rect 165671 248147 165699 248175
rect 165485 248085 165513 248113
rect 165547 248085 165575 248113
rect 165609 248085 165637 248113
rect 165671 248085 165699 248113
rect 165485 248023 165513 248051
rect 165547 248023 165575 248051
rect 165609 248023 165637 248051
rect 165671 248023 165699 248051
rect 165485 247961 165513 247989
rect 165547 247961 165575 247989
rect 165609 247961 165637 247989
rect 165671 247961 165699 247989
rect 165485 239147 165513 239175
rect 165547 239147 165575 239175
rect 165609 239147 165637 239175
rect 165671 239147 165699 239175
rect 165485 239085 165513 239113
rect 165547 239085 165575 239113
rect 165609 239085 165637 239113
rect 165671 239085 165699 239113
rect 165485 239023 165513 239051
rect 165547 239023 165575 239051
rect 165609 239023 165637 239051
rect 165671 239023 165699 239051
rect 165485 238961 165513 238989
rect 165547 238961 165575 238989
rect 165609 238961 165637 238989
rect 165671 238961 165699 238989
rect 165485 230147 165513 230175
rect 165547 230147 165575 230175
rect 165609 230147 165637 230175
rect 165671 230147 165699 230175
rect 165485 230085 165513 230113
rect 165547 230085 165575 230113
rect 165609 230085 165637 230113
rect 165671 230085 165699 230113
rect 165485 230023 165513 230051
rect 165547 230023 165575 230051
rect 165609 230023 165637 230051
rect 165671 230023 165699 230051
rect 165485 229961 165513 229989
rect 165547 229961 165575 229989
rect 165609 229961 165637 229989
rect 165671 229961 165699 229989
rect 165485 221147 165513 221175
rect 165547 221147 165575 221175
rect 165609 221147 165637 221175
rect 165671 221147 165699 221175
rect 165485 221085 165513 221113
rect 165547 221085 165575 221113
rect 165609 221085 165637 221113
rect 165671 221085 165699 221113
rect 165485 221023 165513 221051
rect 165547 221023 165575 221051
rect 165609 221023 165637 221051
rect 165671 221023 165699 221051
rect 165485 220961 165513 220989
rect 165547 220961 165575 220989
rect 165609 220961 165637 220989
rect 165671 220961 165699 220989
rect 165485 212147 165513 212175
rect 165547 212147 165575 212175
rect 165609 212147 165637 212175
rect 165671 212147 165699 212175
rect 165485 212085 165513 212113
rect 165547 212085 165575 212113
rect 165609 212085 165637 212113
rect 165671 212085 165699 212113
rect 165485 212023 165513 212051
rect 165547 212023 165575 212051
rect 165609 212023 165637 212051
rect 165671 212023 165699 212051
rect 165485 211961 165513 211989
rect 165547 211961 165575 211989
rect 165609 211961 165637 211989
rect 165671 211961 165699 211989
rect 165485 203147 165513 203175
rect 165547 203147 165575 203175
rect 165609 203147 165637 203175
rect 165671 203147 165699 203175
rect 165485 203085 165513 203113
rect 165547 203085 165575 203113
rect 165609 203085 165637 203113
rect 165671 203085 165699 203113
rect 165485 203023 165513 203051
rect 165547 203023 165575 203051
rect 165609 203023 165637 203051
rect 165671 203023 165699 203051
rect 165485 202961 165513 202989
rect 165547 202961 165575 202989
rect 165609 202961 165637 202989
rect 165671 202961 165699 202989
rect 165485 194147 165513 194175
rect 165547 194147 165575 194175
rect 165609 194147 165637 194175
rect 165671 194147 165699 194175
rect 165485 194085 165513 194113
rect 165547 194085 165575 194113
rect 165609 194085 165637 194113
rect 165671 194085 165699 194113
rect 165485 194023 165513 194051
rect 165547 194023 165575 194051
rect 165609 194023 165637 194051
rect 165671 194023 165699 194051
rect 165485 193961 165513 193989
rect 165547 193961 165575 193989
rect 165609 193961 165637 193989
rect 165671 193961 165699 193989
rect 165485 185147 165513 185175
rect 165547 185147 165575 185175
rect 165609 185147 165637 185175
rect 165671 185147 165699 185175
rect 165485 185085 165513 185113
rect 165547 185085 165575 185113
rect 165609 185085 165637 185113
rect 165671 185085 165699 185113
rect 165485 185023 165513 185051
rect 165547 185023 165575 185051
rect 165609 185023 165637 185051
rect 165671 185023 165699 185051
rect 165485 184961 165513 184989
rect 165547 184961 165575 184989
rect 165609 184961 165637 184989
rect 165671 184961 165699 184989
rect 165485 176147 165513 176175
rect 165547 176147 165575 176175
rect 165609 176147 165637 176175
rect 165671 176147 165699 176175
rect 165485 176085 165513 176113
rect 165547 176085 165575 176113
rect 165609 176085 165637 176113
rect 165671 176085 165699 176113
rect 165485 176023 165513 176051
rect 165547 176023 165575 176051
rect 165609 176023 165637 176051
rect 165671 176023 165699 176051
rect 165485 175961 165513 175989
rect 165547 175961 165575 175989
rect 165609 175961 165637 175989
rect 165671 175961 165699 175989
rect 165485 167147 165513 167175
rect 165547 167147 165575 167175
rect 165609 167147 165637 167175
rect 165671 167147 165699 167175
rect 165485 167085 165513 167113
rect 165547 167085 165575 167113
rect 165609 167085 165637 167113
rect 165671 167085 165699 167113
rect 165485 167023 165513 167051
rect 165547 167023 165575 167051
rect 165609 167023 165637 167051
rect 165671 167023 165699 167051
rect 165485 166961 165513 166989
rect 165547 166961 165575 166989
rect 165609 166961 165637 166989
rect 165671 166961 165699 166989
rect 165485 158147 165513 158175
rect 165547 158147 165575 158175
rect 165609 158147 165637 158175
rect 165671 158147 165699 158175
rect 165485 158085 165513 158113
rect 165547 158085 165575 158113
rect 165609 158085 165637 158113
rect 165671 158085 165699 158113
rect 165485 158023 165513 158051
rect 165547 158023 165575 158051
rect 165609 158023 165637 158051
rect 165671 158023 165699 158051
rect 165485 157961 165513 157989
rect 165547 157961 165575 157989
rect 165609 157961 165637 157989
rect 165671 157961 165699 157989
rect 165485 149147 165513 149175
rect 165547 149147 165575 149175
rect 165609 149147 165637 149175
rect 165671 149147 165699 149175
rect 165485 149085 165513 149113
rect 165547 149085 165575 149113
rect 165609 149085 165637 149113
rect 165671 149085 165699 149113
rect 165485 149023 165513 149051
rect 165547 149023 165575 149051
rect 165609 149023 165637 149051
rect 165671 149023 165699 149051
rect 165485 148961 165513 148989
rect 165547 148961 165575 148989
rect 165609 148961 165637 148989
rect 165671 148961 165699 148989
rect 165485 140147 165513 140175
rect 165547 140147 165575 140175
rect 165609 140147 165637 140175
rect 165671 140147 165699 140175
rect 165485 140085 165513 140113
rect 165547 140085 165575 140113
rect 165609 140085 165637 140113
rect 165671 140085 165699 140113
rect 165485 140023 165513 140051
rect 165547 140023 165575 140051
rect 165609 140023 165637 140051
rect 165671 140023 165699 140051
rect 165485 139961 165513 139989
rect 165547 139961 165575 139989
rect 165609 139961 165637 139989
rect 165671 139961 165699 139989
rect 165485 131147 165513 131175
rect 165547 131147 165575 131175
rect 165609 131147 165637 131175
rect 165671 131147 165699 131175
rect 165485 131085 165513 131113
rect 165547 131085 165575 131113
rect 165609 131085 165637 131113
rect 165671 131085 165699 131113
rect 165485 131023 165513 131051
rect 165547 131023 165575 131051
rect 165609 131023 165637 131051
rect 165671 131023 165699 131051
rect 165485 130961 165513 130989
rect 165547 130961 165575 130989
rect 165609 130961 165637 130989
rect 165671 130961 165699 130989
rect 165485 122147 165513 122175
rect 165547 122147 165575 122175
rect 165609 122147 165637 122175
rect 165671 122147 165699 122175
rect 165485 122085 165513 122113
rect 165547 122085 165575 122113
rect 165609 122085 165637 122113
rect 165671 122085 165699 122113
rect 165485 122023 165513 122051
rect 165547 122023 165575 122051
rect 165609 122023 165637 122051
rect 165671 122023 165699 122051
rect 165485 121961 165513 121989
rect 165547 121961 165575 121989
rect 165609 121961 165637 121989
rect 165671 121961 165699 121989
rect 165485 113147 165513 113175
rect 165547 113147 165575 113175
rect 165609 113147 165637 113175
rect 165671 113147 165699 113175
rect 165485 113085 165513 113113
rect 165547 113085 165575 113113
rect 165609 113085 165637 113113
rect 165671 113085 165699 113113
rect 165485 113023 165513 113051
rect 165547 113023 165575 113051
rect 165609 113023 165637 113051
rect 165671 113023 165699 113051
rect 165485 112961 165513 112989
rect 165547 112961 165575 112989
rect 165609 112961 165637 112989
rect 165671 112961 165699 112989
rect 165485 104147 165513 104175
rect 165547 104147 165575 104175
rect 165609 104147 165637 104175
rect 165671 104147 165699 104175
rect 165485 104085 165513 104113
rect 165547 104085 165575 104113
rect 165609 104085 165637 104113
rect 165671 104085 165699 104113
rect 165485 104023 165513 104051
rect 165547 104023 165575 104051
rect 165609 104023 165637 104051
rect 165671 104023 165699 104051
rect 165485 103961 165513 103989
rect 165547 103961 165575 103989
rect 165609 103961 165637 103989
rect 165671 103961 165699 103989
rect 165485 95147 165513 95175
rect 165547 95147 165575 95175
rect 165609 95147 165637 95175
rect 165671 95147 165699 95175
rect 165485 95085 165513 95113
rect 165547 95085 165575 95113
rect 165609 95085 165637 95113
rect 165671 95085 165699 95113
rect 165485 95023 165513 95051
rect 165547 95023 165575 95051
rect 165609 95023 165637 95051
rect 165671 95023 165699 95051
rect 165485 94961 165513 94989
rect 165547 94961 165575 94989
rect 165609 94961 165637 94989
rect 165671 94961 165699 94989
rect 165485 86147 165513 86175
rect 165547 86147 165575 86175
rect 165609 86147 165637 86175
rect 165671 86147 165699 86175
rect 165485 86085 165513 86113
rect 165547 86085 165575 86113
rect 165609 86085 165637 86113
rect 165671 86085 165699 86113
rect 165485 86023 165513 86051
rect 165547 86023 165575 86051
rect 165609 86023 165637 86051
rect 165671 86023 165699 86051
rect 165485 85961 165513 85989
rect 165547 85961 165575 85989
rect 165609 85961 165637 85989
rect 165671 85961 165699 85989
rect 165485 77147 165513 77175
rect 165547 77147 165575 77175
rect 165609 77147 165637 77175
rect 165671 77147 165699 77175
rect 165485 77085 165513 77113
rect 165547 77085 165575 77113
rect 165609 77085 165637 77113
rect 165671 77085 165699 77113
rect 165485 77023 165513 77051
rect 165547 77023 165575 77051
rect 165609 77023 165637 77051
rect 165671 77023 165699 77051
rect 165485 76961 165513 76989
rect 165547 76961 165575 76989
rect 165609 76961 165637 76989
rect 165671 76961 165699 76989
rect 165485 68147 165513 68175
rect 165547 68147 165575 68175
rect 165609 68147 165637 68175
rect 165671 68147 165699 68175
rect 165485 68085 165513 68113
rect 165547 68085 165575 68113
rect 165609 68085 165637 68113
rect 165671 68085 165699 68113
rect 165485 68023 165513 68051
rect 165547 68023 165575 68051
rect 165609 68023 165637 68051
rect 165671 68023 165699 68051
rect 165485 67961 165513 67989
rect 165547 67961 165575 67989
rect 165609 67961 165637 67989
rect 165671 67961 165699 67989
rect 165485 59147 165513 59175
rect 165547 59147 165575 59175
rect 165609 59147 165637 59175
rect 165671 59147 165699 59175
rect 165485 59085 165513 59113
rect 165547 59085 165575 59113
rect 165609 59085 165637 59113
rect 165671 59085 165699 59113
rect 165485 59023 165513 59051
rect 165547 59023 165575 59051
rect 165609 59023 165637 59051
rect 165671 59023 165699 59051
rect 165485 58961 165513 58989
rect 165547 58961 165575 58989
rect 165609 58961 165637 58989
rect 165671 58961 165699 58989
rect 165485 50147 165513 50175
rect 165547 50147 165575 50175
rect 165609 50147 165637 50175
rect 165671 50147 165699 50175
rect 165485 50085 165513 50113
rect 165547 50085 165575 50113
rect 165609 50085 165637 50113
rect 165671 50085 165699 50113
rect 165485 50023 165513 50051
rect 165547 50023 165575 50051
rect 165609 50023 165637 50051
rect 165671 50023 165699 50051
rect 165485 49961 165513 49989
rect 165547 49961 165575 49989
rect 165609 49961 165637 49989
rect 165671 49961 165699 49989
rect 165485 41147 165513 41175
rect 165547 41147 165575 41175
rect 165609 41147 165637 41175
rect 165671 41147 165699 41175
rect 165485 41085 165513 41113
rect 165547 41085 165575 41113
rect 165609 41085 165637 41113
rect 165671 41085 165699 41113
rect 165485 41023 165513 41051
rect 165547 41023 165575 41051
rect 165609 41023 165637 41051
rect 165671 41023 165699 41051
rect 165485 40961 165513 40989
rect 165547 40961 165575 40989
rect 165609 40961 165637 40989
rect 165671 40961 165699 40989
rect 165485 32147 165513 32175
rect 165547 32147 165575 32175
rect 165609 32147 165637 32175
rect 165671 32147 165699 32175
rect 165485 32085 165513 32113
rect 165547 32085 165575 32113
rect 165609 32085 165637 32113
rect 165671 32085 165699 32113
rect 165485 32023 165513 32051
rect 165547 32023 165575 32051
rect 165609 32023 165637 32051
rect 165671 32023 165699 32051
rect 165485 31961 165513 31989
rect 165547 31961 165575 31989
rect 165609 31961 165637 31989
rect 165671 31961 165699 31989
rect 165485 23147 165513 23175
rect 165547 23147 165575 23175
rect 165609 23147 165637 23175
rect 165671 23147 165699 23175
rect 165485 23085 165513 23113
rect 165547 23085 165575 23113
rect 165609 23085 165637 23113
rect 165671 23085 165699 23113
rect 165485 23023 165513 23051
rect 165547 23023 165575 23051
rect 165609 23023 165637 23051
rect 165671 23023 165699 23051
rect 165485 22961 165513 22989
rect 165547 22961 165575 22989
rect 165609 22961 165637 22989
rect 165671 22961 165699 22989
rect 165485 14147 165513 14175
rect 165547 14147 165575 14175
rect 165609 14147 165637 14175
rect 165671 14147 165699 14175
rect 165485 14085 165513 14113
rect 165547 14085 165575 14113
rect 165609 14085 165637 14113
rect 165671 14085 165699 14113
rect 165485 14023 165513 14051
rect 165547 14023 165575 14051
rect 165609 14023 165637 14051
rect 165671 14023 165699 14051
rect 165485 13961 165513 13989
rect 165547 13961 165575 13989
rect 165609 13961 165637 13989
rect 165671 13961 165699 13989
rect 165485 5147 165513 5175
rect 165547 5147 165575 5175
rect 165609 5147 165637 5175
rect 165671 5147 165699 5175
rect 165485 5085 165513 5113
rect 165547 5085 165575 5113
rect 165609 5085 165637 5113
rect 165671 5085 165699 5113
rect 165485 5023 165513 5051
rect 165547 5023 165575 5051
rect 165609 5023 165637 5051
rect 165671 5023 165699 5051
rect 165485 4961 165513 4989
rect 165547 4961 165575 4989
rect 165609 4961 165637 4989
rect 165671 4961 165699 4989
rect 165485 -588 165513 -560
rect 165547 -588 165575 -560
rect 165609 -588 165637 -560
rect 165671 -588 165699 -560
rect 165485 -650 165513 -622
rect 165547 -650 165575 -622
rect 165609 -650 165637 -622
rect 165671 -650 165699 -622
rect 165485 -712 165513 -684
rect 165547 -712 165575 -684
rect 165609 -712 165637 -684
rect 165671 -712 165699 -684
rect 165485 -774 165513 -746
rect 165547 -774 165575 -746
rect 165609 -774 165637 -746
rect 165671 -774 165699 -746
rect 172625 298578 172653 298606
rect 172687 298578 172715 298606
rect 172749 298578 172777 298606
rect 172811 298578 172839 298606
rect 172625 298516 172653 298544
rect 172687 298516 172715 298544
rect 172749 298516 172777 298544
rect 172811 298516 172839 298544
rect 172625 298454 172653 298482
rect 172687 298454 172715 298482
rect 172749 298454 172777 298482
rect 172811 298454 172839 298482
rect 172625 298392 172653 298420
rect 172687 298392 172715 298420
rect 172749 298392 172777 298420
rect 172811 298392 172839 298420
rect 172625 290147 172653 290175
rect 172687 290147 172715 290175
rect 172749 290147 172777 290175
rect 172811 290147 172839 290175
rect 172625 290085 172653 290113
rect 172687 290085 172715 290113
rect 172749 290085 172777 290113
rect 172811 290085 172839 290113
rect 172625 290023 172653 290051
rect 172687 290023 172715 290051
rect 172749 290023 172777 290051
rect 172811 290023 172839 290051
rect 172625 289961 172653 289989
rect 172687 289961 172715 289989
rect 172749 289961 172777 289989
rect 172811 289961 172839 289989
rect 172625 281147 172653 281175
rect 172687 281147 172715 281175
rect 172749 281147 172777 281175
rect 172811 281147 172839 281175
rect 172625 281085 172653 281113
rect 172687 281085 172715 281113
rect 172749 281085 172777 281113
rect 172811 281085 172839 281113
rect 172625 281023 172653 281051
rect 172687 281023 172715 281051
rect 172749 281023 172777 281051
rect 172811 281023 172839 281051
rect 172625 280961 172653 280989
rect 172687 280961 172715 280989
rect 172749 280961 172777 280989
rect 172811 280961 172839 280989
rect 172625 272147 172653 272175
rect 172687 272147 172715 272175
rect 172749 272147 172777 272175
rect 172811 272147 172839 272175
rect 172625 272085 172653 272113
rect 172687 272085 172715 272113
rect 172749 272085 172777 272113
rect 172811 272085 172839 272113
rect 172625 272023 172653 272051
rect 172687 272023 172715 272051
rect 172749 272023 172777 272051
rect 172811 272023 172839 272051
rect 172625 271961 172653 271989
rect 172687 271961 172715 271989
rect 172749 271961 172777 271989
rect 172811 271961 172839 271989
rect 172625 263147 172653 263175
rect 172687 263147 172715 263175
rect 172749 263147 172777 263175
rect 172811 263147 172839 263175
rect 172625 263085 172653 263113
rect 172687 263085 172715 263113
rect 172749 263085 172777 263113
rect 172811 263085 172839 263113
rect 172625 263023 172653 263051
rect 172687 263023 172715 263051
rect 172749 263023 172777 263051
rect 172811 263023 172839 263051
rect 172625 262961 172653 262989
rect 172687 262961 172715 262989
rect 172749 262961 172777 262989
rect 172811 262961 172839 262989
rect 172625 254147 172653 254175
rect 172687 254147 172715 254175
rect 172749 254147 172777 254175
rect 172811 254147 172839 254175
rect 172625 254085 172653 254113
rect 172687 254085 172715 254113
rect 172749 254085 172777 254113
rect 172811 254085 172839 254113
rect 172625 254023 172653 254051
rect 172687 254023 172715 254051
rect 172749 254023 172777 254051
rect 172811 254023 172839 254051
rect 172625 253961 172653 253989
rect 172687 253961 172715 253989
rect 172749 253961 172777 253989
rect 172811 253961 172839 253989
rect 172625 245147 172653 245175
rect 172687 245147 172715 245175
rect 172749 245147 172777 245175
rect 172811 245147 172839 245175
rect 172625 245085 172653 245113
rect 172687 245085 172715 245113
rect 172749 245085 172777 245113
rect 172811 245085 172839 245113
rect 172625 245023 172653 245051
rect 172687 245023 172715 245051
rect 172749 245023 172777 245051
rect 172811 245023 172839 245051
rect 172625 244961 172653 244989
rect 172687 244961 172715 244989
rect 172749 244961 172777 244989
rect 172811 244961 172839 244989
rect 172625 236147 172653 236175
rect 172687 236147 172715 236175
rect 172749 236147 172777 236175
rect 172811 236147 172839 236175
rect 172625 236085 172653 236113
rect 172687 236085 172715 236113
rect 172749 236085 172777 236113
rect 172811 236085 172839 236113
rect 172625 236023 172653 236051
rect 172687 236023 172715 236051
rect 172749 236023 172777 236051
rect 172811 236023 172839 236051
rect 172625 235961 172653 235989
rect 172687 235961 172715 235989
rect 172749 235961 172777 235989
rect 172811 235961 172839 235989
rect 172625 227147 172653 227175
rect 172687 227147 172715 227175
rect 172749 227147 172777 227175
rect 172811 227147 172839 227175
rect 172625 227085 172653 227113
rect 172687 227085 172715 227113
rect 172749 227085 172777 227113
rect 172811 227085 172839 227113
rect 172625 227023 172653 227051
rect 172687 227023 172715 227051
rect 172749 227023 172777 227051
rect 172811 227023 172839 227051
rect 172625 226961 172653 226989
rect 172687 226961 172715 226989
rect 172749 226961 172777 226989
rect 172811 226961 172839 226989
rect 172625 218147 172653 218175
rect 172687 218147 172715 218175
rect 172749 218147 172777 218175
rect 172811 218147 172839 218175
rect 172625 218085 172653 218113
rect 172687 218085 172715 218113
rect 172749 218085 172777 218113
rect 172811 218085 172839 218113
rect 172625 218023 172653 218051
rect 172687 218023 172715 218051
rect 172749 218023 172777 218051
rect 172811 218023 172839 218051
rect 172625 217961 172653 217989
rect 172687 217961 172715 217989
rect 172749 217961 172777 217989
rect 172811 217961 172839 217989
rect 172625 209147 172653 209175
rect 172687 209147 172715 209175
rect 172749 209147 172777 209175
rect 172811 209147 172839 209175
rect 172625 209085 172653 209113
rect 172687 209085 172715 209113
rect 172749 209085 172777 209113
rect 172811 209085 172839 209113
rect 172625 209023 172653 209051
rect 172687 209023 172715 209051
rect 172749 209023 172777 209051
rect 172811 209023 172839 209051
rect 172625 208961 172653 208989
rect 172687 208961 172715 208989
rect 172749 208961 172777 208989
rect 172811 208961 172839 208989
rect 172625 200147 172653 200175
rect 172687 200147 172715 200175
rect 172749 200147 172777 200175
rect 172811 200147 172839 200175
rect 172625 200085 172653 200113
rect 172687 200085 172715 200113
rect 172749 200085 172777 200113
rect 172811 200085 172839 200113
rect 172625 200023 172653 200051
rect 172687 200023 172715 200051
rect 172749 200023 172777 200051
rect 172811 200023 172839 200051
rect 172625 199961 172653 199989
rect 172687 199961 172715 199989
rect 172749 199961 172777 199989
rect 172811 199961 172839 199989
rect 172625 191147 172653 191175
rect 172687 191147 172715 191175
rect 172749 191147 172777 191175
rect 172811 191147 172839 191175
rect 172625 191085 172653 191113
rect 172687 191085 172715 191113
rect 172749 191085 172777 191113
rect 172811 191085 172839 191113
rect 172625 191023 172653 191051
rect 172687 191023 172715 191051
rect 172749 191023 172777 191051
rect 172811 191023 172839 191051
rect 172625 190961 172653 190989
rect 172687 190961 172715 190989
rect 172749 190961 172777 190989
rect 172811 190961 172839 190989
rect 172625 182147 172653 182175
rect 172687 182147 172715 182175
rect 172749 182147 172777 182175
rect 172811 182147 172839 182175
rect 172625 182085 172653 182113
rect 172687 182085 172715 182113
rect 172749 182085 172777 182113
rect 172811 182085 172839 182113
rect 172625 182023 172653 182051
rect 172687 182023 172715 182051
rect 172749 182023 172777 182051
rect 172811 182023 172839 182051
rect 172625 181961 172653 181989
rect 172687 181961 172715 181989
rect 172749 181961 172777 181989
rect 172811 181961 172839 181989
rect 172625 173147 172653 173175
rect 172687 173147 172715 173175
rect 172749 173147 172777 173175
rect 172811 173147 172839 173175
rect 172625 173085 172653 173113
rect 172687 173085 172715 173113
rect 172749 173085 172777 173113
rect 172811 173085 172839 173113
rect 172625 173023 172653 173051
rect 172687 173023 172715 173051
rect 172749 173023 172777 173051
rect 172811 173023 172839 173051
rect 172625 172961 172653 172989
rect 172687 172961 172715 172989
rect 172749 172961 172777 172989
rect 172811 172961 172839 172989
rect 172625 164147 172653 164175
rect 172687 164147 172715 164175
rect 172749 164147 172777 164175
rect 172811 164147 172839 164175
rect 172625 164085 172653 164113
rect 172687 164085 172715 164113
rect 172749 164085 172777 164113
rect 172811 164085 172839 164113
rect 172625 164023 172653 164051
rect 172687 164023 172715 164051
rect 172749 164023 172777 164051
rect 172811 164023 172839 164051
rect 172625 163961 172653 163989
rect 172687 163961 172715 163989
rect 172749 163961 172777 163989
rect 172811 163961 172839 163989
rect 172625 155147 172653 155175
rect 172687 155147 172715 155175
rect 172749 155147 172777 155175
rect 172811 155147 172839 155175
rect 172625 155085 172653 155113
rect 172687 155085 172715 155113
rect 172749 155085 172777 155113
rect 172811 155085 172839 155113
rect 172625 155023 172653 155051
rect 172687 155023 172715 155051
rect 172749 155023 172777 155051
rect 172811 155023 172839 155051
rect 172625 154961 172653 154989
rect 172687 154961 172715 154989
rect 172749 154961 172777 154989
rect 172811 154961 172839 154989
rect 172625 146147 172653 146175
rect 172687 146147 172715 146175
rect 172749 146147 172777 146175
rect 172811 146147 172839 146175
rect 172625 146085 172653 146113
rect 172687 146085 172715 146113
rect 172749 146085 172777 146113
rect 172811 146085 172839 146113
rect 172625 146023 172653 146051
rect 172687 146023 172715 146051
rect 172749 146023 172777 146051
rect 172811 146023 172839 146051
rect 172625 145961 172653 145989
rect 172687 145961 172715 145989
rect 172749 145961 172777 145989
rect 172811 145961 172839 145989
rect 172625 137147 172653 137175
rect 172687 137147 172715 137175
rect 172749 137147 172777 137175
rect 172811 137147 172839 137175
rect 172625 137085 172653 137113
rect 172687 137085 172715 137113
rect 172749 137085 172777 137113
rect 172811 137085 172839 137113
rect 172625 137023 172653 137051
rect 172687 137023 172715 137051
rect 172749 137023 172777 137051
rect 172811 137023 172839 137051
rect 172625 136961 172653 136989
rect 172687 136961 172715 136989
rect 172749 136961 172777 136989
rect 172811 136961 172839 136989
rect 172625 128147 172653 128175
rect 172687 128147 172715 128175
rect 172749 128147 172777 128175
rect 172811 128147 172839 128175
rect 172625 128085 172653 128113
rect 172687 128085 172715 128113
rect 172749 128085 172777 128113
rect 172811 128085 172839 128113
rect 172625 128023 172653 128051
rect 172687 128023 172715 128051
rect 172749 128023 172777 128051
rect 172811 128023 172839 128051
rect 172625 127961 172653 127989
rect 172687 127961 172715 127989
rect 172749 127961 172777 127989
rect 172811 127961 172839 127989
rect 172625 119147 172653 119175
rect 172687 119147 172715 119175
rect 172749 119147 172777 119175
rect 172811 119147 172839 119175
rect 172625 119085 172653 119113
rect 172687 119085 172715 119113
rect 172749 119085 172777 119113
rect 172811 119085 172839 119113
rect 172625 119023 172653 119051
rect 172687 119023 172715 119051
rect 172749 119023 172777 119051
rect 172811 119023 172839 119051
rect 172625 118961 172653 118989
rect 172687 118961 172715 118989
rect 172749 118961 172777 118989
rect 172811 118961 172839 118989
rect 172625 110147 172653 110175
rect 172687 110147 172715 110175
rect 172749 110147 172777 110175
rect 172811 110147 172839 110175
rect 172625 110085 172653 110113
rect 172687 110085 172715 110113
rect 172749 110085 172777 110113
rect 172811 110085 172839 110113
rect 172625 110023 172653 110051
rect 172687 110023 172715 110051
rect 172749 110023 172777 110051
rect 172811 110023 172839 110051
rect 172625 109961 172653 109989
rect 172687 109961 172715 109989
rect 172749 109961 172777 109989
rect 172811 109961 172839 109989
rect 172625 101147 172653 101175
rect 172687 101147 172715 101175
rect 172749 101147 172777 101175
rect 172811 101147 172839 101175
rect 172625 101085 172653 101113
rect 172687 101085 172715 101113
rect 172749 101085 172777 101113
rect 172811 101085 172839 101113
rect 172625 101023 172653 101051
rect 172687 101023 172715 101051
rect 172749 101023 172777 101051
rect 172811 101023 172839 101051
rect 172625 100961 172653 100989
rect 172687 100961 172715 100989
rect 172749 100961 172777 100989
rect 172811 100961 172839 100989
rect 172625 92147 172653 92175
rect 172687 92147 172715 92175
rect 172749 92147 172777 92175
rect 172811 92147 172839 92175
rect 172625 92085 172653 92113
rect 172687 92085 172715 92113
rect 172749 92085 172777 92113
rect 172811 92085 172839 92113
rect 172625 92023 172653 92051
rect 172687 92023 172715 92051
rect 172749 92023 172777 92051
rect 172811 92023 172839 92051
rect 172625 91961 172653 91989
rect 172687 91961 172715 91989
rect 172749 91961 172777 91989
rect 172811 91961 172839 91989
rect 172625 83147 172653 83175
rect 172687 83147 172715 83175
rect 172749 83147 172777 83175
rect 172811 83147 172839 83175
rect 172625 83085 172653 83113
rect 172687 83085 172715 83113
rect 172749 83085 172777 83113
rect 172811 83085 172839 83113
rect 172625 83023 172653 83051
rect 172687 83023 172715 83051
rect 172749 83023 172777 83051
rect 172811 83023 172839 83051
rect 172625 82961 172653 82989
rect 172687 82961 172715 82989
rect 172749 82961 172777 82989
rect 172811 82961 172839 82989
rect 172625 74147 172653 74175
rect 172687 74147 172715 74175
rect 172749 74147 172777 74175
rect 172811 74147 172839 74175
rect 172625 74085 172653 74113
rect 172687 74085 172715 74113
rect 172749 74085 172777 74113
rect 172811 74085 172839 74113
rect 172625 74023 172653 74051
rect 172687 74023 172715 74051
rect 172749 74023 172777 74051
rect 172811 74023 172839 74051
rect 172625 73961 172653 73989
rect 172687 73961 172715 73989
rect 172749 73961 172777 73989
rect 172811 73961 172839 73989
rect 172625 65147 172653 65175
rect 172687 65147 172715 65175
rect 172749 65147 172777 65175
rect 172811 65147 172839 65175
rect 172625 65085 172653 65113
rect 172687 65085 172715 65113
rect 172749 65085 172777 65113
rect 172811 65085 172839 65113
rect 172625 65023 172653 65051
rect 172687 65023 172715 65051
rect 172749 65023 172777 65051
rect 172811 65023 172839 65051
rect 172625 64961 172653 64989
rect 172687 64961 172715 64989
rect 172749 64961 172777 64989
rect 172811 64961 172839 64989
rect 172625 56147 172653 56175
rect 172687 56147 172715 56175
rect 172749 56147 172777 56175
rect 172811 56147 172839 56175
rect 172625 56085 172653 56113
rect 172687 56085 172715 56113
rect 172749 56085 172777 56113
rect 172811 56085 172839 56113
rect 172625 56023 172653 56051
rect 172687 56023 172715 56051
rect 172749 56023 172777 56051
rect 172811 56023 172839 56051
rect 172625 55961 172653 55989
rect 172687 55961 172715 55989
rect 172749 55961 172777 55989
rect 172811 55961 172839 55989
rect 172625 47147 172653 47175
rect 172687 47147 172715 47175
rect 172749 47147 172777 47175
rect 172811 47147 172839 47175
rect 172625 47085 172653 47113
rect 172687 47085 172715 47113
rect 172749 47085 172777 47113
rect 172811 47085 172839 47113
rect 172625 47023 172653 47051
rect 172687 47023 172715 47051
rect 172749 47023 172777 47051
rect 172811 47023 172839 47051
rect 172625 46961 172653 46989
rect 172687 46961 172715 46989
rect 172749 46961 172777 46989
rect 172811 46961 172839 46989
rect 172625 38147 172653 38175
rect 172687 38147 172715 38175
rect 172749 38147 172777 38175
rect 172811 38147 172839 38175
rect 172625 38085 172653 38113
rect 172687 38085 172715 38113
rect 172749 38085 172777 38113
rect 172811 38085 172839 38113
rect 172625 38023 172653 38051
rect 172687 38023 172715 38051
rect 172749 38023 172777 38051
rect 172811 38023 172839 38051
rect 172625 37961 172653 37989
rect 172687 37961 172715 37989
rect 172749 37961 172777 37989
rect 172811 37961 172839 37989
rect 172625 29147 172653 29175
rect 172687 29147 172715 29175
rect 172749 29147 172777 29175
rect 172811 29147 172839 29175
rect 172625 29085 172653 29113
rect 172687 29085 172715 29113
rect 172749 29085 172777 29113
rect 172811 29085 172839 29113
rect 172625 29023 172653 29051
rect 172687 29023 172715 29051
rect 172749 29023 172777 29051
rect 172811 29023 172839 29051
rect 172625 28961 172653 28989
rect 172687 28961 172715 28989
rect 172749 28961 172777 28989
rect 172811 28961 172839 28989
rect 172625 20147 172653 20175
rect 172687 20147 172715 20175
rect 172749 20147 172777 20175
rect 172811 20147 172839 20175
rect 172625 20085 172653 20113
rect 172687 20085 172715 20113
rect 172749 20085 172777 20113
rect 172811 20085 172839 20113
rect 172625 20023 172653 20051
rect 172687 20023 172715 20051
rect 172749 20023 172777 20051
rect 172811 20023 172839 20051
rect 172625 19961 172653 19989
rect 172687 19961 172715 19989
rect 172749 19961 172777 19989
rect 172811 19961 172839 19989
rect 172625 11147 172653 11175
rect 172687 11147 172715 11175
rect 172749 11147 172777 11175
rect 172811 11147 172839 11175
rect 172625 11085 172653 11113
rect 172687 11085 172715 11113
rect 172749 11085 172777 11113
rect 172811 11085 172839 11113
rect 172625 11023 172653 11051
rect 172687 11023 172715 11051
rect 172749 11023 172777 11051
rect 172811 11023 172839 11051
rect 172625 10961 172653 10989
rect 172687 10961 172715 10989
rect 172749 10961 172777 10989
rect 172811 10961 172839 10989
rect 172625 2147 172653 2175
rect 172687 2147 172715 2175
rect 172749 2147 172777 2175
rect 172811 2147 172839 2175
rect 172625 2085 172653 2113
rect 172687 2085 172715 2113
rect 172749 2085 172777 2113
rect 172811 2085 172839 2113
rect 172625 2023 172653 2051
rect 172687 2023 172715 2051
rect 172749 2023 172777 2051
rect 172811 2023 172839 2051
rect 172625 1961 172653 1989
rect 172687 1961 172715 1989
rect 172749 1961 172777 1989
rect 172811 1961 172839 1989
rect 172625 -108 172653 -80
rect 172687 -108 172715 -80
rect 172749 -108 172777 -80
rect 172811 -108 172839 -80
rect 172625 -170 172653 -142
rect 172687 -170 172715 -142
rect 172749 -170 172777 -142
rect 172811 -170 172839 -142
rect 172625 -232 172653 -204
rect 172687 -232 172715 -204
rect 172749 -232 172777 -204
rect 172811 -232 172839 -204
rect 172625 -294 172653 -266
rect 172687 -294 172715 -266
rect 172749 -294 172777 -266
rect 172811 -294 172839 -266
rect 174485 299058 174513 299086
rect 174547 299058 174575 299086
rect 174609 299058 174637 299086
rect 174671 299058 174699 299086
rect 174485 298996 174513 299024
rect 174547 298996 174575 299024
rect 174609 298996 174637 299024
rect 174671 298996 174699 299024
rect 174485 298934 174513 298962
rect 174547 298934 174575 298962
rect 174609 298934 174637 298962
rect 174671 298934 174699 298962
rect 174485 298872 174513 298900
rect 174547 298872 174575 298900
rect 174609 298872 174637 298900
rect 174671 298872 174699 298900
rect 174485 293147 174513 293175
rect 174547 293147 174575 293175
rect 174609 293147 174637 293175
rect 174671 293147 174699 293175
rect 174485 293085 174513 293113
rect 174547 293085 174575 293113
rect 174609 293085 174637 293113
rect 174671 293085 174699 293113
rect 174485 293023 174513 293051
rect 174547 293023 174575 293051
rect 174609 293023 174637 293051
rect 174671 293023 174699 293051
rect 174485 292961 174513 292989
rect 174547 292961 174575 292989
rect 174609 292961 174637 292989
rect 174671 292961 174699 292989
rect 174485 284147 174513 284175
rect 174547 284147 174575 284175
rect 174609 284147 174637 284175
rect 174671 284147 174699 284175
rect 174485 284085 174513 284113
rect 174547 284085 174575 284113
rect 174609 284085 174637 284113
rect 174671 284085 174699 284113
rect 174485 284023 174513 284051
rect 174547 284023 174575 284051
rect 174609 284023 174637 284051
rect 174671 284023 174699 284051
rect 174485 283961 174513 283989
rect 174547 283961 174575 283989
rect 174609 283961 174637 283989
rect 174671 283961 174699 283989
rect 174485 275147 174513 275175
rect 174547 275147 174575 275175
rect 174609 275147 174637 275175
rect 174671 275147 174699 275175
rect 174485 275085 174513 275113
rect 174547 275085 174575 275113
rect 174609 275085 174637 275113
rect 174671 275085 174699 275113
rect 174485 275023 174513 275051
rect 174547 275023 174575 275051
rect 174609 275023 174637 275051
rect 174671 275023 174699 275051
rect 174485 274961 174513 274989
rect 174547 274961 174575 274989
rect 174609 274961 174637 274989
rect 174671 274961 174699 274989
rect 174485 266147 174513 266175
rect 174547 266147 174575 266175
rect 174609 266147 174637 266175
rect 174671 266147 174699 266175
rect 174485 266085 174513 266113
rect 174547 266085 174575 266113
rect 174609 266085 174637 266113
rect 174671 266085 174699 266113
rect 174485 266023 174513 266051
rect 174547 266023 174575 266051
rect 174609 266023 174637 266051
rect 174671 266023 174699 266051
rect 174485 265961 174513 265989
rect 174547 265961 174575 265989
rect 174609 265961 174637 265989
rect 174671 265961 174699 265989
rect 174485 257147 174513 257175
rect 174547 257147 174575 257175
rect 174609 257147 174637 257175
rect 174671 257147 174699 257175
rect 174485 257085 174513 257113
rect 174547 257085 174575 257113
rect 174609 257085 174637 257113
rect 174671 257085 174699 257113
rect 174485 257023 174513 257051
rect 174547 257023 174575 257051
rect 174609 257023 174637 257051
rect 174671 257023 174699 257051
rect 174485 256961 174513 256989
rect 174547 256961 174575 256989
rect 174609 256961 174637 256989
rect 174671 256961 174699 256989
rect 174485 248147 174513 248175
rect 174547 248147 174575 248175
rect 174609 248147 174637 248175
rect 174671 248147 174699 248175
rect 174485 248085 174513 248113
rect 174547 248085 174575 248113
rect 174609 248085 174637 248113
rect 174671 248085 174699 248113
rect 174485 248023 174513 248051
rect 174547 248023 174575 248051
rect 174609 248023 174637 248051
rect 174671 248023 174699 248051
rect 174485 247961 174513 247989
rect 174547 247961 174575 247989
rect 174609 247961 174637 247989
rect 174671 247961 174699 247989
rect 174485 239147 174513 239175
rect 174547 239147 174575 239175
rect 174609 239147 174637 239175
rect 174671 239147 174699 239175
rect 174485 239085 174513 239113
rect 174547 239085 174575 239113
rect 174609 239085 174637 239113
rect 174671 239085 174699 239113
rect 174485 239023 174513 239051
rect 174547 239023 174575 239051
rect 174609 239023 174637 239051
rect 174671 239023 174699 239051
rect 174485 238961 174513 238989
rect 174547 238961 174575 238989
rect 174609 238961 174637 238989
rect 174671 238961 174699 238989
rect 174485 230147 174513 230175
rect 174547 230147 174575 230175
rect 174609 230147 174637 230175
rect 174671 230147 174699 230175
rect 174485 230085 174513 230113
rect 174547 230085 174575 230113
rect 174609 230085 174637 230113
rect 174671 230085 174699 230113
rect 174485 230023 174513 230051
rect 174547 230023 174575 230051
rect 174609 230023 174637 230051
rect 174671 230023 174699 230051
rect 174485 229961 174513 229989
rect 174547 229961 174575 229989
rect 174609 229961 174637 229989
rect 174671 229961 174699 229989
rect 174485 221147 174513 221175
rect 174547 221147 174575 221175
rect 174609 221147 174637 221175
rect 174671 221147 174699 221175
rect 174485 221085 174513 221113
rect 174547 221085 174575 221113
rect 174609 221085 174637 221113
rect 174671 221085 174699 221113
rect 174485 221023 174513 221051
rect 174547 221023 174575 221051
rect 174609 221023 174637 221051
rect 174671 221023 174699 221051
rect 174485 220961 174513 220989
rect 174547 220961 174575 220989
rect 174609 220961 174637 220989
rect 174671 220961 174699 220989
rect 174485 212147 174513 212175
rect 174547 212147 174575 212175
rect 174609 212147 174637 212175
rect 174671 212147 174699 212175
rect 174485 212085 174513 212113
rect 174547 212085 174575 212113
rect 174609 212085 174637 212113
rect 174671 212085 174699 212113
rect 174485 212023 174513 212051
rect 174547 212023 174575 212051
rect 174609 212023 174637 212051
rect 174671 212023 174699 212051
rect 174485 211961 174513 211989
rect 174547 211961 174575 211989
rect 174609 211961 174637 211989
rect 174671 211961 174699 211989
rect 174485 203147 174513 203175
rect 174547 203147 174575 203175
rect 174609 203147 174637 203175
rect 174671 203147 174699 203175
rect 174485 203085 174513 203113
rect 174547 203085 174575 203113
rect 174609 203085 174637 203113
rect 174671 203085 174699 203113
rect 174485 203023 174513 203051
rect 174547 203023 174575 203051
rect 174609 203023 174637 203051
rect 174671 203023 174699 203051
rect 174485 202961 174513 202989
rect 174547 202961 174575 202989
rect 174609 202961 174637 202989
rect 174671 202961 174699 202989
rect 174485 194147 174513 194175
rect 174547 194147 174575 194175
rect 174609 194147 174637 194175
rect 174671 194147 174699 194175
rect 174485 194085 174513 194113
rect 174547 194085 174575 194113
rect 174609 194085 174637 194113
rect 174671 194085 174699 194113
rect 174485 194023 174513 194051
rect 174547 194023 174575 194051
rect 174609 194023 174637 194051
rect 174671 194023 174699 194051
rect 174485 193961 174513 193989
rect 174547 193961 174575 193989
rect 174609 193961 174637 193989
rect 174671 193961 174699 193989
rect 174485 185147 174513 185175
rect 174547 185147 174575 185175
rect 174609 185147 174637 185175
rect 174671 185147 174699 185175
rect 174485 185085 174513 185113
rect 174547 185085 174575 185113
rect 174609 185085 174637 185113
rect 174671 185085 174699 185113
rect 174485 185023 174513 185051
rect 174547 185023 174575 185051
rect 174609 185023 174637 185051
rect 174671 185023 174699 185051
rect 174485 184961 174513 184989
rect 174547 184961 174575 184989
rect 174609 184961 174637 184989
rect 174671 184961 174699 184989
rect 174485 176147 174513 176175
rect 174547 176147 174575 176175
rect 174609 176147 174637 176175
rect 174671 176147 174699 176175
rect 174485 176085 174513 176113
rect 174547 176085 174575 176113
rect 174609 176085 174637 176113
rect 174671 176085 174699 176113
rect 174485 176023 174513 176051
rect 174547 176023 174575 176051
rect 174609 176023 174637 176051
rect 174671 176023 174699 176051
rect 174485 175961 174513 175989
rect 174547 175961 174575 175989
rect 174609 175961 174637 175989
rect 174671 175961 174699 175989
rect 174485 167147 174513 167175
rect 174547 167147 174575 167175
rect 174609 167147 174637 167175
rect 174671 167147 174699 167175
rect 174485 167085 174513 167113
rect 174547 167085 174575 167113
rect 174609 167085 174637 167113
rect 174671 167085 174699 167113
rect 174485 167023 174513 167051
rect 174547 167023 174575 167051
rect 174609 167023 174637 167051
rect 174671 167023 174699 167051
rect 174485 166961 174513 166989
rect 174547 166961 174575 166989
rect 174609 166961 174637 166989
rect 174671 166961 174699 166989
rect 174485 158147 174513 158175
rect 174547 158147 174575 158175
rect 174609 158147 174637 158175
rect 174671 158147 174699 158175
rect 174485 158085 174513 158113
rect 174547 158085 174575 158113
rect 174609 158085 174637 158113
rect 174671 158085 174699 158113
rect 174485 158023 174513 158051
rect 174547 158023 174575 158051
rect 174609 158023 174637 158051
rect 174671 158023 174699 158051
rect 174485 157961 174513 157989
rect 174547 157961 174575 157989
rect 174609 157961 174637 157989
rect 174671 157961 174699 157989
rect 174485 149147 174513 149175
rect 174547 149147 174575 149175
rect 174609 149147 174637 149175
rect 174671 149147 174699 149175
rect 174485 149085 174513 149113
rect 174547 149085 174575 149113
rect 174609 149085 174637 149113
rect 174671 149085 174699 149113
rect 174485 149023 174513 149051
rect 174547 149023 174575 149051
rect 174609 149023 174637 149051
rect 174671 149023 174699 149051
rect 174485 148961 174513 148989
rect 174547 148961 174575 148989
rect 174609 148961 174637 148989
rect 174671 148961 174699 148989
rect 174485 140147 174513 140175
rect 174547 140147 174575 140175
rect 174609 140147 174637 140175
rect 174671 140147 174699 140175
rect 174485 140085 174513 140113
rect 174547 140085 174575 140113
rect 174609 140085 174637 140113
rect 174671 140085 174699 140113
rect 174485 140023 174513 140051
rect 174547 140023 174575 140051
rect 174609 140023 174637 140051
rect 174671 140023 174699 140051
rect 174485 139961 174513 139989
rect 174547 139961 174575 139989
rect 174609 139961 174637 139989
rect 174671 139961 174699 139989
rect 174485 131147 174513 131175
rect 174547 131147 174575 131175
rect 174609 131147 174637 131175
rect 174671 131147 174699 131175
rect 174485 131085 174513 131113
rect 174547 131085 174575 131113
rect 174609 131085 174637 131113
rect 174671 131085 174699 131113
rect 174485 131023 174513 131051
rect 174547 131023 174575 131051
rect 174609 131023 174637 131051
rect 174671 131023 174699 131051
rect 174485 130961 174513 130989
rect 174547 130961 174575 130989
rect 174609 130961 174637 130989
rect 174671 130961 174699 130989
rect 174485 122147 174513 122175
rect 174547 122147 174575 122175
rect 174609 122147 174637 122175
rect 174671 122147 174699 122175
rect 174485 122085 174513 122113
rect 174547 122085 174575 122113
rect 174609 122085 174637 122113
rect 174671 122085 174699 122113
rect 174485 122023 174513 122051
rect 174547 122023 174575 122051
rect 174609 122023 174637 122051
rect 174671 122023 174699 122051
rect 174485 121961 174513 121989
rect 174547 121961 174575 121989
rect 174609 121961 174637 121989
rect 174671 121961 174699 121989
rect 174485 113147 174513 113175
rect 174547 113147 174575 113175
rect 174609 113147 174637 113175
rect 174671 113147 174699 113175
rect 174485 113085 174513 113113
rect 174547 113085 174575 113113
rect 174609 113085 174637 113113
rect 174671 113085 174699 113113
rect 174485 113023 174513 113051
rect 174547 113023 174575 113051
rect 174609 113023 174637 113051
rect 174671 113023 174699 113051
rect 174485 112961 174513 112989
rect 174547 112961 174575 112989
rect 174609 112961 174637 112989
rect 174671 112961 174699 112989
rect 174485 104147 174513 104175
rect 174547 104147 174575 104175
rect 174609 104147 174637 104175
rect 174671 104147 174699 104175
rect 174485 104085 174513 104113
rect 174547 104085 174575 104113
rect 174609 104085 174637 104113
rect 174671 104085 174699 104113
rect 174485 104023 174513 104051
rect 174547 104023 174575 104051
rect 174609 104023 174637 104051
rect 174671 104023 174699 104051
rect 174485 103961 174513 103989
rect 174547 103961 174575 103989
rect 174609 103961 174637 103989
rect 174671 103961 174699 103989
rect 174485 95147 174513 95175
rect 174547 95147 174575 95175
rect 174609 95147 174637 95175
rect 174671 95147 174699 95175
rect 174485 95085 174513 95113
rect 174547 95085 174575 95113
rect 174609 95085 174637 95113
rect 174671 95085 174699 95113
rect 174485 95023 174513 95051
rect 174547 95023 174575 95051
rect 174609 95023 174637 95051
rect 174671 95023 174699 95051
rect 174485 94961 174513 94989
rect 174547 94961 174575 94989
rect 174609 94961 174637 94989
rect 174671 94961 174699 94989
rect 174485 86147 174513 86175
rect 174547 86147 174575 86175
rect 174609 86147 174637 86175
rect 174671 86147 174699 86175
rect 174485 86085 174513 86113
rect 174547 86085 174575 86113
rect 174609 86085 174637 86113
rect 174671 86085 174699 86113
rect 174485 86023 174513 86051
rect 174547 86023 174575 86051
rect 174609 86023 174637 86051
rect 174671 86023 174699 86051
rect 174485 85961 174513 85989
rect 174547 85961 174575 85989
rect 174609 85961 174637 85989
rect 174671 85961 174699 85989
rect 174485 77147 174513 77175
rect 174547 77147 174575 77175
rect 174609 77147 174637 77175
rect 174671 77147 174699 77175
rect 174485 77085 174513 77113
rect 174547 77085 174575 77113
rect 174609 77085 174637 77113
rect 174671 77085 174699 77113
rect 174485 77023 174513 77051
rect 174547 77023 174575 77051
rect 174609 77023 174637 77051
rect 174671 77023 174699 77051
rect 174485 76961 174513 76989
rect 174547 76961 174575 76989
rect 174609 76961 174637 76989
rect 174671 76961 174699 76989
rect 174485 68147 174513 68175
rect 174547 68147 174575 68175
rect 174609 68147 174637 68175
rect 174671 68147 174699 68175
rect 174485 68085 174513 68113
rect 174547 68085 174575 68113
rect 174609 68085 174637 68113
rect 174671 68085 174699 68113
rect 174485 68023 174513 68051
rect 174547 68023 174575 68051
rect 174609 68023 174637 68051
rect 174671 68023 174699 68051
rect 174485 67961 174513 67989
rect 174547 67961 174575 67989
rect 174609 67961 174637 67989
rect 174671 67961 174699 67989
rect 174485 59147 174513 59175
rect 174547 59147 174575 59175
rect 174609 59147 174637 59175
rect 174671 59147 174699 59175
rect 174485 59085 174513 59113
rect 174547 59085 174575 59113
rect 174609 59085 174637 59113
rect 174671 59085 174699 59113
rect 174485 59023 174513 59051
rect 174547 59023 174575 59051
rect 174609 59023 174637 59051
rect 174671 59023 174699 59051
rect 174485 58961 174513 58989
rect 174547 58961 174575 58989
rect 174609 58961 174637 58989
rect 174671 58961 174699 58989
rect 174485 50147 174513 50175
rect 174547 50147 174575 50175
rect 174609 50147 174637 50175
rect 174671 50147 174699 50175
rect 174485 50085 174513 50113
rect 174547 50085 174575 50113
rect 174609 50085 174637 50113
rect 174671 50085 174699 50113
rect 174485 50023 174513 50051
rect 174547 50023 174575 50051
rect 174609 50023 174637 50051
rect 174671 50023 174699 50051
rect 174485 49961 174513 49989
rect 174547 49961 174575 49989
rect 174609 49961 174637 49989
rect 174671 49961 174699 49989
rect 174485 41147 174513 41175
rect 174547 41147 174575 41175
rect 174609 41147 174637 41175
rect 174671 41147 174699 41175
rect 174485 41085 174513 41113
rect 174547 41085 174575 41113
rect 174609 41085 174637 41113
rect 174671 41085 174699 41113
rect 174485 41023 174513 41051
rect 174547 41023 174575 41051
rect 174609 41023 174637 41051
rect 174671 41023 174699 41051
rect 174485 40961 174513 40989
rect 174547 40961 174575 40989
rect 174609 40961 174637 40989
rect 174671 40961 174699 40989
rect 174485 32147 174513 32175
rect 174547 32147 174575 32175
rect 174609 32147 174637 32175
rect 174671 32147 174699 32175
rect 174485 32085 174513 32113
rect 174547 32085 174575 32113
rect 174609 32085 174637 32113
rect 174671 32085 174699 32113
rect 174485 32023 174513 32051
rect 174547 32023 174575 32051
rect 174609 32023 174637 32051
rect 174671 32023 174699 32051
rect 174485 31961 174513 31989
rect 174547 31961 174575 31989
rect 174609 31961 174637 31989
rect 174671 31961 174699 31989
rect 174485 23147 174513 23175
rect 174547 23147 174575 23175
rect 174609 23147 174637 23175
rect 174671 23147 174699 23175
rect 174485 23085 174513 23113
rect 174547 23085 174575 23113
rect 174609 23085 174637 23113
rect 174671 23085 174699 23113
rect 174485 23023 174513 23051
rect 174547 23023 174575 23051
rect 174609 23023 174637 23051
rect 174671 23023 174699 23051
rect 174485 22961 174513 22989
rect 174547 22961 174575 22989
rect 174609 22961 174637 22989
rect 174671 22961 174699 22989
rect 174485 14147 174513 14175
rect 174547 14147 174575 14175
rect 174609 14147 174637 14175
rect 174671 14147 174699 14175
rect 174485 14085 174513 14113
rect 174547 14085 174575 14113
rect 174609 14085 174637 14113
rect 174671 14085 174699 14113
rect 174485 14023 174513 14051
rect 174547 14023 174575 14051
rect 174609 14023 174637 14051
rect 174671 14023 174699 14051
rect 174485 13961 174513 13989
rect 174547 13961 174575 13989
rect 174609 13961 174637 13989
rect 174671 13961 174699 13989
rect 174485 5147 174513 5175
rect 174547 5147 174575 5175
rect 174609 5147 174637 5175
rect 174671 5147 174699 5175
rect 174485 5085 174513 5113
rect 174547 5085 174575 5113
rect 174609 5085 174637 5113
rect 174671 5085 174699 5113
rect 174485 5023 174513 5051
rect 174547 5023 174575 5051
rect 174609 5023 174637 5051
rect 174671 5023 174699 5051
rect 174485 4961 174513 4989
rect 174547 4961 174575 4989
rect 174609 4961 174637 4989
rect 174671 4961 174699 4989
rect 174485 -588 174513 -560
rect 174547 -588 174575 -560
rect 174609 -588 174637 -560
rect 174671 -588 174699 -560
rect 174485 -650 174513 -622
rect 174547 -650 174575 -622
rect 174609 -650 174637 -622
rect 174671 -650 174699 -622
rect 174485 -712 174513 -684
rect 174547 -712 174575 -684
rect 174609 -712 174637 -684
rect 174671 -712 174699 -684
rect 174485 -774 174513 -746
rect 174547 -774 174575 -746
rect 174609 -774 174637 -746
rect 174671 -774 174699 -746
rect 181625 298578 181653 298606
rect 181687 298578 181715 298606
rect 181749 298578 181777 298606
rect 181811 298578 181839 298606
rect 181625 298516 181653 298544
rect 181687 298516 181715 298544
rect 181749 298516 181777 298544
rect 181811 298516 181839 298544
rect 181625 298454 181653 298482
rect 181687 298454 181715 298482
rect 181749 298454 181777 298482
rect 181811 298454 181839 298482
rect 181625 298392 181653 298420
rect 181687 298392 181715 298420
rect 181749 298392 181777 298420
rect 181811 298392 181839 298420
rect 181625 290147 181653 290175
rect 181687 290147 181715 290175
rect 181749 290147 181777 290175
rect 181811 290147 181839 290175
rect 181625 290085 181653 290113
rect 181687 290085 181715 290113
rect 181749 290085 181777 290113
rect 181811 290085 181839 290113
rect 181625 290023 181653 290051
rect 181687 290023 181715 290051
rect 181749 290023 181777 290051
rect 181811 290023 181839 290051
rect 181625 289961 181653 289989
rect 181687 289961 181715 289989
rect 181749 289961 181777 289989
rect 181811 289961 181839 289989
rect 181625 281147 181653 281175
rect 181687 281147 181715 281175
rect 181749 281147 181777 281175
rect 181811 281147 181839 281175
rect 181625 281085 181653 281113
rect 181687 281085 181715 281113
rect 181749 281085 181777 281113
rect 181811 281085 181839 281113
rect 181625 281023 181653 281051
rect 181687 281023 181715 281051
rect 181749 281023 181777 281051
rect 181811 281023 181839 281051
rect 181625 280961 181653 280989
rect 181687 280961 181715 280989
rect 181749 280961 181777 280989
rect 181811 280961 181839 280989
rect 181625 272147 181653 272175
rect 181687 272147 181715 272175
rect 181749 272147 181777 272175
rect 181811 272147 181839 272175
rect 181625 272085 181653 272113
rect 181687 272085 181715 272113
rect 181749 272085 181777 272113
rect 181811 272085 181839 272113
rect 181625 272023 181653 272051
rect 181687 272023 181715 272051
rect 181749 272023 181777 272051
rect 181811 272023 181839 272051
rect 181625 271961 181653 271989
rect 181687 271961 181715 271989
rect 181749 271961 181777 271989
rect 181811 271961 181839 271989
rect 181625 263147 181653 263175
rect 181687 263147 181715 263175
rect 181749 263147 181777 263175
rect 181811 263147 181839 263175
rect 181625 263085 181653 263113
rect 181687 263085 181715 263113
rect 181749 263085 181777 263113
rect 181811 263085 181839 263113
rect 181625 263023 181653 263051
rect 181687 263023 181715 263051
rect 181749 263023 181777 263051
rect 181811 263023 181839 263051
rect 181625 262961 181653 262989
rect 181687 262961 181715 262989
rect 181749 262961 181777 262989
rect 181811 262961 181839 262989
rect 181625 254147 181653 254175
rect 181687 254147 181715 254175
rect 181749 254147 181777 254175
rect 181811 254147 181839 254175
rect 181625 254085 181653 254113
rect 181687 254085 181715 254113
rect 181749 254085 181777 254113
rect 181811 254085 181839 254113
rect 181625 254023 181653 254051
rect 181687 254023 181715 254051
rect 181749 254023 181777 254051
rect 181811 254023 181839 254051
rect 181625 253961 181653 253989
rect 181687 253961 181715 253989
rect 181749 253961 181777 253989
rect 181811 253961 181839 253989
rect 181625 245147 181653 245175
rect 181687 245147 181715 245175
rect 181749 245147 181777 245175
rect 181811 245147 181839 245175
rect 181625 245085 181653 245113
rect 181687 245085 181715 245113
rect 181749 245085 181777 245113
rect 181811 245085 181839 245113
rect 181625 245023 181653 245051
rect 181687 245023 181715 245051
rect 181749 245023 181777 245051
rect 181811 245023 181839 245051
rect 181625 244961 181653 244989
rect 181687 244961 181715 244989
rect 181749 244961 181777 244989
rect 181811 244961 181839 244989
rect 181625 236147 181653 236175
rect 181687 236147 181715 236175
rect 181749 236147 181777 236175
rect 181811 236147 181839 236175
rect 181625 236085 181653 236113
rect 181687 236085 181715 236113
rect 181749 236085 181777 236113
rect 181811 236085 181839 236113
rect 181625 236023 181653 236051
rect 181687 236023 181715 236051
rect 181749 236023 181777 236051
rect 181811 236023 181839 236051
rect 181625 235961 181653 235989
rect 181687 235961 181715 235989
rect 181749 235961 181777 235989
rect 181811 235961 181839 235989
rect 181625 227147 181653 227175
rect 181687 227147 181715 227175
rect 181749 227147 181777 227175
rect 181811 227147 181839 227175
rect 181625 227085 181653 227113
rect 181687 227085 181715 227113
rect 181749 227085 181777 227113
rect 181811 227085 181839 227113
rect 181625 227023 181653 227051
rect 181687 227023 181715 227051
rect 181749 227023 181777 227051
rect 181811 227023 181839 227051
rect 181625 226961 181653 226989
rect 181687 226961 181715 226989
rect 181749 226961 181777 226989
rect 181811 226961 181839 226989
rect 181625 218147 181653 218175
rect 181687 218147 181715 218175
rect 181749 218147 181777 218175
rect 181811 218147 181839 218175
rect 181625 218085 181653 218113
rect 181687 218085 181715 218113
rect 181749 218085 181777 218113
rect 181811 218085 181839 218113
rect 181625 218023 181653 218051
rect 181687 218023 181715 218051
rect 181749 218023 181777 218051
rect 181811 218023 181839 218051
rect 181625 217961 181653 217989
rect 181687 217961 181715 217989
rect 181749 217961 181777 217989
rect 181811 217961 181839 217989
rect 181625 209147 181653 209175
rect 181687 209147 181715 209175
rect 181749 209147 181777 209175
rect 181811 209147 181839 209175
rect 181625 209085 181653 209113
rect 181687 209085 181715 209113
rect 181749 209085 181777 209113
rect 181811 209085 181839 209113
rect 181625 209023 181653 209051
rect 181687 209023 181715 209051
rect 181749 209023 181777 209051
rect 181811 209023 181839 209051
rect 181625 208961 181653 208989
rect 181687 208961 181715 208989
rect 181749 208961 181777 208989
rect 181811 208961 181839 208989
rect 181625 200147 181653 200175
rect 181687 200147 181715 200175
rect 181749 200147 181777 200175
rect 181811 200147 181839 200175
rect 181625 200085 181653 200113
rect 181687 200085 181715 200113
rect 181749 200085 181777 200113
rect 181811 200085 181839 200113
rect 181625 200023 181653 200051
rect 181687 200023 181715 200051
rect 181749 200023 181777 200051
rect 181811 200023 181839 200051
rect 181625 199961 181653 199989
rect 181687 199961 181715 199989
rect 181749 199961 181777 199989
rect 181811 199961 181839 199989
rect 181625 191147 181653 191175
rect 181687 191147 181715 191175
rect 181749 191147 181777 191175
rect 181811 191147 181839 191175
rect 181625 191085 181653 191113
rect 181687 191085 181715 191113
rect 181749 191085 181777 191113
rect 181811 191085 181839 191113
rect 181625 191023 181653 191051
rect 181687 191023 181715 191051
rect 181749 191023 181777 191051
rect 181811 191023 181839 191051
rect 181625 190961 181653 190989
rect 181687 190961 181715 190989
rect 181749 190961 181777 190989
rect 181811 190961 181839 190989
rect 181625 182147 181653 182175
rect 181687 182147 181715 182175
rect 181749 182147 181777 182175
rect 181811 182147 181839 182175
rect 181625 182085 181653 182113
rect 181687 182085 181715 182113
rect 181749 182085 181777 182113
rect 181811 182085 181839 182113
rect 181625 182023 181653 182051
rect 181687 182023 181715 182051
rect 181749 182023 181777 182051
rect 181811 182023 181839 182051
rect 181625 181961 181653 181989
rect 181687 181961 181715 181989
rect 181749 181961 181777 181989
rect 181811 181961 181839 181989
rect 181625 173147 181653 173175
rect 181687 173147 181715 173175
rect 181749 173147 181777 173175
rect 181811 173147 181839 173175
rect 181625 173085 181653 173113
rect 181687 173085 181715 173113
rect 181749 173085 181777 173113
rect 181811 173085 181839 173113
rect 181625 173023 181653 173051
rect 181687 173023 181715 173051
rect 181749 173023 181777 173051
rect 181811 173023 181839 173051
rect 181625 172961 181653 172989
rect 181687 172961 181715 172989
rect 181749 172961 181777 172989
rect 181811 172961 181839 172989
rect 181625 164147 181653 164175
rect 181687 164147 181715 164175
rect 181749 164147 181777 164175
rect 181811 164147 181839 164175
rect 181625 164085 181653 164113
rect 181687 164085 181715 164113
rect 181749 164085 181777 164113
rect 181811 164085 181839 164113
rect 181625 164023 181653 164051
rect 181687 164023 181715 164051
rect 181749 164023 181777 164051
rect 181811 164023 181839 164051
rect 181625 163961 181653 163989
rect 181687 163961 181715 163989
rect 181749 163961 181777 163989
rect 181811 163961 181839 163989
rect 181625 155147 181653 155175
rect 181687 155147 181715 155175
rect 181749 155147 181777 155175
rect 181811 155147 181839 155175
rect 181625 155085 181653 155113
rect 181687 155085 181715 155113
rect 181749 155085 181777 155113
rect 181811 155085 181839 155113
rect 181625 155023 181653 155051
rect 181687 155023 181715 155051
rect 181749 155023 181777 155051
rect 181811 155023 181839 155051
rect 181625 154961 181653 154989
rect 181687 154961 181715 154989
rect 181749 154961 181777 154989
rect 181811 154961 181839 154989
rect 181625 146147 181653 146175
rect 181687 146147 181715 146175
rect 181749 146147 181777 146175
rect 181811 146147 181839 146175
rect 181625 146085 181653 146113
rect 181687 146085 181715 146113
rect 181749 146085 181777 146113
rect 181811 146085 181839 146113
rect 181625 146023 181653 146051
rect 181687 146023 181715 146051
rect 181749 146023 181777 146051
rect 181811 146023 181839 146051
rect 181625 145961 181653 145989
rect 181687 145961 181715 145989
rect 181749 145961 181777 145989
rect 181811 145961 181839 145989
rect 181625 137147 181653 137175
rect 181687 137147 181715 137175
rect 181749 137147 181777 137175
rect 181811 137147 181839 137175
rect 181625 137085 181653 137113
rect 181687 137085 181715 137113
rect 181749 137085 181777 137113
rect 181811 137085 181839 137113
rect 181625 137023 181653 137051
rect 181687 137023 181715 137051
rect 181749 137023 181777 137051
rect 181811 137023 181839 137051
rect 181625 136961 181653 136989
rect 181687 136961 181715 136989
rect 181749 136961 181777 136989
rect 181811 136961 181839 136989
rect 181625 128147 181653 128175
rect 181687 128147 181715 128175
rect 181749 128147 181777 128175
rect 181811 128147 181839 128175
rect 181625 128085 181653 128113
rect 181687 128085 181715 128113
rect 181749 128085 181777 128113
rect 181811 128085 181839 128113
rect 181625 128023 181653 128051
rect 181687 128023 181715 128051
rect 181749 128023 181777 128051
rect 181811 128023 181839 128051
rect 181625 127961 181653 127989
rect 181687 127961 181715 127989
rect 181749 127961 181777 127989
rect 181811 127961 181839 127989
rect 181625 119147 181653 119175
rect 181687 119147 181715 119175
rect 181749 119147 181777 119175
rect 181811 119147 181839 119175
rect 181625 119085 181653 119113
rect 181687 119085 181715 119113
rect 181749 119085 181777 119113
rect 181811 119085 181839 119113
rect 181625 119023 181653 119051
rect 181687 119023 181715 119051
rect 181749 119023 181777 119051
rect 181811 119023 181839 119051
rect 181625 118961 181653 118989
rect 181687 118961 181715 118989
rect 181749 118961 181777 118989
rect 181811 118961 181839 118989
rect 181625 110147 181653 110175
rect 181687 110147 181715 110175
rect 181749 110147 181777 110175
rect 181811 110147 181839 110175
rect 181625 110085 181653 110113
rect 181687 110085 181715 110113
rect 181749 110085 181777 110113
rect 181811 110085 181839 110113
rect 181625 110023 181653 110051
rect 181687 110023 181715 110051
rect 181749 110023 181777 110051
rect 181811 110023 181839 110051
rect 181625 109961 181653 109989
rect 181687 109961 181715 109989
rect 181749 109961 181777 109989
rect 181811 109961 181839 109989
rect 181625 101147 181653 101175
rect 181687 101147 181715 101175
rect 181749 101147 181777 101175
rect 181811 101147 181839 101175
rect 181625 101085 181653 101113
rect 181687 101085 181715 101113
rect 181749 101085 181777 101113
rect 181811 101085 181839 101113
rect 181625 101023 181653 101051
rect 181687 101023 181715 101051
rect 181749 101023 181777 101051
rect 181811 101023 181839 101051
rect 181625 100961 181653 100989
rect 181687 100961 181715 100989
rect 181749 100961 181777 100989
rect 181811 100961 181839 100989
rect 181625 92147 181653 92175
rect 181687 92147 181715 92175
rect 181749 92147 181777 92175
rect 181811 92147 181839 92175
rect 181625 92085 181653 92113
rect 181687 92085 181715 92113
rect 181749 92085 181777 92113
rect 181811 92085 181839 92113
rect 181625 92023 181653 92051
rect 181687 92023 181715 92051
rect 181749 92023 181777 92051
rect 181811 92023 181839 92051
rect 181625 91961 181653 91989
rect 181687 91961 181715 91989
rect 181749 91961 181777 91989
rect 181811 91961 181839 91989
rect 181625 83147 181653 83175
rect 181687 83147 181715 83175
rect 181749 83147 181777 83175
rect 181811 83147 181839 83175
rect 181625 83085 181653 83113
rect 181687 83085 181715 83113
rect 181749 83085 181777 83113
rect 181811 83085 181839 83113
rect 181625 83023 181653 83051
rect 181687 83023 181715 83051
rect 181749 83023 181777 83051
rect 181811 83023 181839 83051
rect 181625 82961 181653 82989
rect 181687 82961 181715 82989
rect 181749 82961 181777 82989
rect 181811 82961 181839 82989
rect 181625 74147 181653 74175
rect 181687 74147 181715 74175
rect 181749 74147 181777 74175
rect 181811 74147 181839 74175
rect 181625 74085 181653 74113
rect 181687 74085 181715 74113
rect 181749 74085 181777 74113
rect 181811 74085 181839 74113
rect 181625 74023 181653 74051
rect 181687 74023 181715 74051
rect 181749 74023 181777 74051
rect 181811 74023 181839 74051
rect 181625 73961 181653 73989
rect 181687 73961 181715 73989
rect 181749 73961 181777 73989
rect 181811 73961 181839 73989
rect 181625 65147 181653 65175
rect 181687 65147 181715 65175
rect 181749 65147 181777 65175
rect 181811 65147 181839 65175
rect 181625 65085 181653 65113
rect 181687 65085 181715 65113
rect 181749 65085 181777 65113
rect 181811 65085 181839 65113
rect 181625 65023 181653 65051
rect 181687 65023 181715 65051
rect 181749 65023 181777 65051
rect 181811 65023 181839 65051
rect 181625 64961 181653 64989
rect 181687 64961 181715 64989
rect 181749 64961 181777 64989
rect 181811 64961 181839 64989
rect 181625 56147 181653 56175
rect 181687 56147 181715 56175
rect 181749 56147 181777 56175
rect 181811 56147 181839 56175
rect 181625 56085 181653 56113
rect 181687 56085 181715 56113
rect 181749 56085 181777 56113
rect 181811 56085 181839 56113
rect 181625 56023 181653 56051
rect 181687 56023 181715 56051
rect 181749 56023 181777 56051
rect 181811 56023 181839 56051
rect 181625 55961 181653 55989
rect 181687 55961 181715 55989
rect 181749 55961 181777 55989
rect 181811 55961 181839 55989
rect 181625 47147 181653 47175
rect 181687 47147 181715 47175
rect 181749 47147 181777 47175
rect 181811 47147 181839 47175
rect 181625 47085 181653 47113
rect 181687 47085 181715 47113
rect 181749 47085 181777 47113
rect 181811 47085 181839 47113
rect 181625 47023 181653 47051
rect 181687 47023 181715 47051
rect 181749 47023 181777 47051
rect 181811 47023 181839 47051
rect 181625 46961 181653 46989
rect 181687 46961 181715 46989
rect 181749 46961 181777 46989
rect 181811 46961 181839 46989
rect 181625 38147 181653 38175
rect 181687 38147 181715 38175
rect 181749 38147 181777 38175
rect 181811 38147 181839 38175
rect 181625 38085 181653 38113
rect 181687 38085 181715 38113
rect 181749 38085 181777 38113
rect 181811 38085 181839 38113
rect 181625 38023 181653 38051
rect 181687 38023 181715 38051
rect 181749 38023 181777 38051
rect 181811 38023 181839 38051
rect 181625 37961 181653 37989
rect 181687 37961 181715 37989
rect 181749 37961 181777 37989
rect 181811 37961 181839 37989
rect 181625 29147 181653 29175
rect 181687 29147 181715 29175
rect 181749 29147 181777 29175
rect 181811 29147 181839 29175
rect 181625 29085 181653 29113
rect 181687 29085 181715 29113
rect 181749 29085 181777 29113
rect 181811 29085 181839 29113
rect 181625 29023 181653 29051
rect 181687 29023 181715 29051
rect 181749 29023 181777 29051
rect 181811 29023 181839 29051
rect 181625 28961 181653 28989
rect 181687 28961 181715 28989
rect 181749 28961 181777 28989
rect 181811 28961 181839 28989
rect 181625 20147 181653 20175
rect 181687 20147 181715 20175
rect 181749 20147 181777 20175
rect 181811 20147 181839 20175
rect 181625 20085 181653 20113
rect 181687 20085 181715 20113
rect 181749 20085 181777 20113
rect 181811 20085 181839 20113
rect 181625 20023 181653 20051
rect 181687 20023 181715 20051
rect 181749 20023 181777 20051
rect 181811 20023 181839 20051
rect 181625 19961 181653 19989
rect 181687 19961 181715 19989
rect 181749 19961 181777 19989
rect 181811 19961 181839 19989
rect 181625 11147 181653 11175
rect 181687 11147 181715 11175
rect 181749 11147 181777 11175
rect 181811 11147 181839 11175
rect 181625 11085 181653 11113
rect 181687 11085 181715 11113
rect 181749 11085 181777 11113
rect 181811 11085 181839 11113
rect 181625 11023 181653 11051
rect 181687 11023 181715 11051
rect 181749 11023 181777 11051
rect 181811 11023 181839 11051
rect 181625 10961 181653 10989
rect 181687 10961 181715 10989
rect 181749 10961 181777 10989
rect 181811 10961 181839 10989
rect 181625 2147 181653 2175
rect 181687 2147 181715 2175
rect 181749 2147 181777 2175
rect 181811 2147 181839 2175
rect 181625 2085 181653 2113
rect 181687 2085 181715 2113
rect 181749 2085 181777 2113
rect 181811 2085 181839 2113
rect 181625 2023 181653 2051
rect 181687 2023 181715 2051
rect 181749 2023 181777 2051
rect 181811 2023 181839 2051
rect 181625 1961 181653 1989
rect 181687 1961 181715 1989
rect 181749 1961 181777 1989
rect 181811 1961 181839 1989
rect 181625 -108 181653 -80
rect 181687 -108 181715 -80
rect 181749 -108 181777 -80
rect 181811 -108 181839 -80
rect 181625 -170 181653 -142
rect 181687 -170 181715 -142
rect 181749 -170 181777 -142
rect 181811 -170 181839 -142
rect 181625 -232 181653 -204
rect 181687 -232 181715 -204
rect 181749 -232 181777 -204
rect 181811 -232 181839 -204
rect 181625 -294 181653 -266
rect 181687 -294 181715 -266
rect 181749 -294 181777 -266
rect 181811 -294 181839 -266
rect 183485 299058 183513 299086
rect 183547 299058 183575 299086
rect 183609 299058 183637 299086
rect 183671 299058 183699 299086
rect 183485 298996 183513 299024
rect 183547 298996 183575 299024
rect 183609 298996 183637 299024
rect 183671 298996 183699 299024
rect 183485 298934 183513 298962
rect 183547 298934 183575 298962
rect 183609 298934 183637 298962
rect 183671 298934 183699 298962
rect 183485 298872 183513 298900
rect 183547 298872 183575 298900
rect 183609 298872 183637 298900
rect 183671 298872 183699 298900
rect 183485 293147 183513 293175
rect 183547 293147 183575 293175
rect 183609 293147 183637 293175
rect 183671 293147 183699 293175
rect 183485 293085 183513 293113
rect 183547 293085 183575 293113
rect 183609 293085 183637 293113
rect 183671 293085 183699 293113
rect 183485 293023 183513 293051
rect 183547 293023 183575 293051
rect 183609 293023 183637 293051
rect 183671 293023 183699 293051
rect 183485 292961 183513 292989
rect 183547 292961 183575 292989
rect 183609 292961 183637 292989
rect 183671 292961 183699 292989
rect 183485 284147 183513 284175
rect 183547 284147 183575 284175
rect 183609 284147 183637 284175
rect 183671 284147 183699 284175
rect 183485 284085 183513 284113
rect 183547 284085 183575 284113
rect 183609 284085 183637 284113
rect 183671 284085 183699 284113
rect 183485 284023 183513 284051
rect 183547 284023 183575 284051
rect 183609 284023 183637 284051
rect 183671 284023 183699 284051
rect 183485 283961 183513 283989
rect 183547 283961 183575 283989
rect 183609 283961 183637 283989
rect 183671 283961 183699 283989
rect 183485 275147 183513 275175
rect 183547 275147 183575 275175
rect 183609 275147 183637 275175
rect 183671 275147 183699 275175
rect 183485 275085 183513 275113
rect 183547 275085 183575 275113
rect 183609 275085 183637 275113
rect 183671 275085 183699 275113
rect 183485 275023 183513 275051
rect 183547 275023 183575 275051
rect 183609 275023 183637 275051
rect 183671 275023 183699 275051
rect 183485 274961 183513 274989
rect 183547 274961 183575 274989
rect 183609 274961 183637 274989
rect 183671 274961 183699 274989
rect 183485 266147 183513 266175
rect 183547 266147 183575 266175
rect 183609 266147 183637 266175
rect 183671 266147 183699 266175
rect 183485 266085 183513 266113
rect 183547 266085 183575 266113
rect 183609 266085 183637 266113
rect 183671 266085 183699 266113
rect 183485 266023 183513 266051
rect 183547 266023 183575 266051
rect 183609 266023 183637 266051
rect 183671 266023 183699 266051
rect 183485 265961 183513 265989
rect 183547 265961 183575 265989
rect 183609 265961 183637 265989
rect 183671 265961 183699 265989
rect 183485 257147 183513 257175
rect 183547 257147 183575 257175
rect 183609 257147 183637 257175
rect 183671 257147 183699 257175
rect 183485 257085 183513 257113
rect 183547 257085 183575 257113
rect 183609 257085 183637 257113
rect 183671 257085 183699 257113
rect 183485 257023 183513 257051
rect 183547 257023 183575 257051
rect 183609 257023 183637 257051
rect 183671 257023 183699 257051
rect 183485 256961 183513 256989
rect 183547 256961 183575 256989
rect 183609 256961 183637 256989
rect 183671 256961 183699 256989
rect 183485 248147 183513 248175
rect 183547 248147 183575 248175
rect 183609 248147 183637 248175
rect 183671 248147 183699 248175
rect 183485 248085 183513 248113
rect 183547 248085 183575 248113
rect 183609 248085 183637 248113
rect 183671 248085 183699 248113
rect 183485 248023 183513 248051
rect 183547 248023 183575 248051
rect 183609 248023 183637 248051
rect 183671 248023 183699 248051
rect 183485 247961 183513 247989
rect 183547 247961 183575 247989
rect 183609 247961 183637 247989
rect 183671 247961 183699 247989
rect 183485 239147 183513 239175
rect 183547 239147 183575 239175
rect 183609 239147 183637 239175
rect 183671 239147 183699 239175
rect 183485 239085 183513 239113
rect 183547 239085 183575 239113
rect 183609 239085 183637 239113
rect 183671 239085 183699 239113
rect 183485 239023 183513 239051
rect 183547 239023 183575 239051
rect 183609 239023 183637 239051
rect 183671 239023 183699 239051
rect 183485 238961 183513 238989
rect 183547 238961 183575 238989
rect 183609 238961 183637 238989
rect 183671 238961 183699 238989
rect 183485 230147 183513 230175
rect 183547 230147 183575 230175
rect 183609 230147 183637 230175
rect 183671 230147 183699 230175
rect 183485 230085 183513 230113
rect 183547 230085 183575 230113
rect 183609 230085 183637 230113
rect 183671 230085 183699 230113
rect 183485 230023 183513 230051
rect 183547 230023 183575 230051
rect 183609 230023 183637 230051
rect 183671 230023 183699 230051
rect 183485 229961 183513 229989
rect 183547 229961 183575 229989
rect 183609 229961 183637 229989
rect 183671 229961 183699 229989
rect 183485 221147 183513 221175
rect 183547 221147 183575 221175
rect 183609 221147 183637 221175
rect 183671 221147 183699 221175
rect 183485 221085 183513 221113
rect 183547 221085 183575 221113
rect 183609 221085 183637 221113
rect 183671 221085 183699 221113
rect 183485 221023 183513 221051
rect 183547 221023 183575 221051
rect 183609 221023 183637 221051
rect 183671 221023 183699 221051
rect 183485 220961 183513 220989
rect 183547 220961 183575 220989
rect 183609 220961 183637 220989
rect 183671 220961 183699 220989
rect 183485 212147 183513 212175
rect 183547 212147 183575 212175
rect 183609 212147 183637 212175
rect 183671 212147 183699 212175
rect 183485 212085 183513 212113
rect 183547 212085 183575 212113
rect 183609 212085 183637 212113
rect 183671 212085 183699 212113
rect 183485 212023 183513 212051
rect 183547 212023 183575 212051
rect 183609 212023 183637 212051
rect 183671 212023 183699 212051
rect 183485 211961 183513 211989
rect 183547 211961 183575 211989
rect 183609 211961 183637 211989
rect 183671 211961 183699 211989
rect 183485 203147 183513 203175
rect 183547 203147 183575 203175
rect 183609 203147 183637 203175
rect 183671 203147 183699 203175
rect 183485 203085 183513 203113
rect 183547 203085 183575 203113
rect 183609 203085 183637 203113
rect 183671 203085 183699 203113
rect 183485 203023 183513 203051
rect 183547 203023 183575 203051
rect 183609 203023 183637 203051
rect 183671 203023 183699 203051
rect 183485 202961 183513 202989
rect 183547 202961 183575 202989
rect 183609 202961 183637 202989
rect 183671 202961 183699 202989
rect 183485 194147 183513 194175
rect 183547 194147 183575 194175
rect 183609 194147 183637 194175
rect 183671 194147 183699 194175
rect 183485 194085 183513 194113
rect 183547 194085 183575 194113
rect 183609 194085 183637 194113
rect 183671 194085 183699 194113
rect 183485 194023 183513 194051
rect 183547 194023 183575 194051
rect 183609 194023 183637 194051
rect 183671 194023 183699 194051
rect 183485 193961 183513 193989
rect 183547 193961 183575 193989
rect 183609 193961 183637 193989
rect 183671 193961 183699 193989
rect 183485 185147 183513 185175
rect 183547 185147 183575 185175
rect 183609 185147 183637 185175
rect 183671 185147 183699 185175
rect 183485 185085 183513 185113
rect 183547 185085 183575 185113
rect 183609 185085 183637 185113
rect 183671 185085 183699 185113
rect 183485 185023 183513 185051
rect 183547 185023 183575 185051
rect 183609 185023 183637 185051
rect 183671 185023 183699 185051
rect 183485 184961 183513 184989
rect 183547 184961 183575 184989
rect 183609 184961 183637 184989
rect 183671 184961 183699 184989
rect 183485 176147 183513 176175
rect 183547 176147 183575 176175
rect 183609 176147 183637 176175
rect 183671 176147 183699 176175
rect 183485 176085 183513 176113
rect 183547 176085 183575 176113
rect 183609 176085 183637 176113
rect 183671 176085 183699 176113
rect 183485 176023 183513 176051
rect 183547 176023 183575 176051
rect 183609 176023 183637 176051
rect 183671 176023 183699 176051
rect 183485 175961 183513 175989
rect 183547 175961 183575 175989
rect 183609 175961 183637 175989
rect 183671 175961 183699 175989
rect 183485 167147 183513 167175
rect 183547 167147 183575 167175
rect 183609 167147 183637 167175
rect 183671 167147 183699 167175
rect 183485 167085 183513 167113
rect 183547 167085 183575 167113
rect 183609 167085 183637 167113
rect 183671 167085 183699 167113
rect 183485 167023 183513 167051
rect 183547 167023 183575 167051
rect 183609 167023 183637 167051
rect 183671 167023 183699 167051
rect 183485 166961 183513 166989
rect 183547 166961 183575 166989
rect 183609 166961 183637 166989
rect 183671 166961 183699 166989
rect 183485 158147 183513 158175
rect 183547 158147 183575 158175
rect 183609 158147 183637 158175
rect 183671 158147 183699 158175
rect 183485 158085 183513 158113
rect 183547 158085 183575 158113
rect 183609 158085 183637 158113
rect 183671 158085 183699 158113
rect 183485 158023 183513 158051
rect 183547 158023 183575 158051
rect 183609 158023 183637 158051
rect 183671 158023 183699 158051
rect 183485 157961 183513 157989
rect 183547 157961 183575 157989
rect 183609 157961 183637 157989
rect 183671 157961 183699 157989
rect 183485 149147 183513 149175
rect 183547 149147 183575 149175
rect 183609 149147 183637 149175
rect 183671 149147 183699 149175
rect 183485 149085 183513 149113
rect 183547 149085 183575 149113
rect 183609 149085 183637 149113
rect 183671 149085 183699 149113
rect 183485 149023 183513 149051
rect 183547 149023 183575 149051
rect 183609 149023 183637 149051
rect 183671 149023 183699 149051
rect 183485 148961 183513 148989
rect 183547 148961 183575 148989
rect 183609 148961 183637 148989
rect 183671 148961 183699 148989
rect 183485 140147 183513 140175
rect 183547 140147 183575 140175
rect 183609 140147 183637 140175
rect 183671 140147 183699 140175
rect 183485 140085 183513 140113
rect 183547 140085 183575 140113
rect 183609 140085 183637 140113
rect 183671 140085 183699 140113
rect 183485 140023 183513 140051
rect 183547 140023 183575 140051
rect 183609 140023 183637 140051
rect 183671 140023 183699 140051
rect 183485 139961 183513 139989
rect 183547 139961 183575 139989
rect 183609 139961 183637 139989
rect 183671 139961 183699 139989
rect 183485 131147 183513 131175
rect 183547 131147 183575 131175
rect 183609 131147 183637 131175
rect 183671 131147 183699 131175
rect 183485 131085 183513 131113
rect 183547 131085 183575 131113
rect 183609 131085 183637 131113
rect 183671 131085 183699 131113
rect 183485 131023 183513 131051
rect 183547 131023 183575 131051
rect 183609 131023 183637 131051
rect 183671 131023 183699 131051
rect 183485 130961 183513 130989
rect 183547 130961 183575 130989
rect 183609 130961 183637 130989
rect 183671 130961 183699 130989
rect 183485 122147 183513 122175
rect 183547 122147 183575 122175
rect 183609 122147 183637 122175
rect 183671 122147 183699 122175
rect 183485 122085 183513 122113
rect 183547 122085 183575 122113
rect 183609 122085 183637 122113
rect 183671 122085 183699 122113
rect 183485 122023 183513 122051
rect 183547 122023 183575 122051
rect 183609 122023 183637 122051
rect 183671 122023 183699 122051
rect 183485 121961 183513 121989
rect 183547 121961 183575 121989
rect 183609 121961 183637 121989
rect 183671 121961 183699 121989
rect 183485 113147 183513 113175
rect 183547 113147 183575 113175
rect 183609 113147 183637 113175
rect 183671 113147 183699 113175
rect 183485 113085 183513 113113
rect 183547 113085 183575 113113
rect 183609 113085 183637 113113
rect 183671 113085 183699 113113
rect 183485 113023 183513 113051
rect 183547 113023 183575 113051
rect 183609 113023 183637 113051
rect 183671 113023 183699 113051
rect 183485 112961 183513 112989
rect 183547 112961 183575 112989
rect 183609 112961 183637 112989
rect 183671 112961 183699 112989
rect 183485 104147 183513 104175
rect 183547 104147 183575 104175
rect 183609 104147 183637 104175
rect 183671 104147 183699 104175
rect 183485 104085 183513 104113
rect 183547 104085 183575 104113
rect 183609 104085 183637 104113
rect 183671 104085 183699 104113
rect 183485 104023 183513 104051
rect 183547 104023 183575 104051
rect 183609 104023 183637 104051
rect 183671 104023 183699 104051
rect 183485 103961 183513 103989
rect 183547 103961 183575 103989
rect 183609 103961 183637 103989
rect 183671 103961 183699 103989
rect 183485 95147 183513 95175
rect 183547 95147 183575 95175
rect 183609 95147 183637 95175
rect 183671 95147 183699 95175
rect 183485 95085 183513 95113
rect 183547 95085 183575 95113
rect 183609 95085 183637 95113
rect 183671 95085 183699 95113
rect 183485 95023 183513 95051
rect 183547 95023 183575 95051
rect 183609 95023 183637 95051
rect 183671 95023 183699 95051
rect 183485 94961 183513 94989
rect 183547 94961 183575 94989
rect 183609 94961 183637 94989
rect 183671 94961 183699 94989
rect 183485 86147 183513 86175
rect 183547 86147 183575 86175
rect 183609 86147 183637 86175
rect 183671 86147 183699 86175
rect 183485 86085 183513 86113
rect 183547 86085 183575 86113
rect 183609 86085 183637 86113
rect 183671 86085 183699 86113
rect 183485 86023 183513 86051
rect 183547 86023 183575 86051
rect 183609 86023 183637 86051
rect 183671 86023 183699 86051
rect 183485 85961 183513 85989
rect 183547 85961 183575 85989
rect 183609 85961 183637 85989
rect 183671 85961 183699 85989
rect 183485 77147 183513 77175
rect 183547 77147 183575 77175
rect 183609 77147 183637 77175
rect 183671 77147 183699 77175
rect 183485 77085 183513 77113
rect 183547 77085 183575 77113
rect 183609 77085 183637 77113
rect 183671 77085 183699 77113
rect 183485 77023 183513 77051
rect 183547 77023 183575 77051
rect 183609 77023 183637 77051
rect 183671 77023 183699 77051
rect 183485 76961 183513 76989
rect 183547 76961 183575 76989
rect 183609 76961 183637 76989
rect 183671 76961 183699 76989
rect 183485 68147 183513 68175
rect 183547 68147 183575 68175
rect 183609 68147 183637 68175
rect 183671 68147 183699 68175
rect 183485 68085 183513 68113
rect 183547 68085 183575 68113
rect 183609 68085 183637 68113
rect 183671 68085 183699 68113
rect 183485 68023 183513 68051
rect 183547 68023 183575 68051
rect 183609 68023 183637 68051
rect 183671 68023 183699 68051
rect 183485 67961 183513 67989
rect 183547 67961 183575 67989
rect 183609 67961 183637 67989
rect 183671 67961 183699 67989
rect 183485 59147 183513 59175
rect 183547 59147 183575 59175
rect 183609 59147 183637 59175
rect 183671 59147 183699 59175
rect 183485 59085 183513 59113
rect 183547 59085 183575 59113
rect 183609 59085 183637 59113
rect 183671 59085 183699 59113
rect 183485 59023 183513 59051
rect 183547 59023 183575 59051
rect 183609 59023 183637 59051
rect 183671 59023 183699 59051
rect 183485 58961 183513 58989
rect 183547 58961 183575 58989
rect 183609 58961 183637 58989
rect 183671 58961 183699 58989
rect 183485 50147 183513 50175
rect 183547 50147 183575 50175
rect 183609 50147 183637 50175
rect 183671 50147 183699 50175
rect 183485 50085 183513 50113
rect 183547 50085 183575 50113
rect 183609 50085 183637 50113
rect 183671 50085 183699 50113
rect 183485 50023 183513 50051
rect 183547 50023 183575 50051
rect 183609 50023 183637 50051
rect 183671 50023 183699 50051
rect 183485 49961 183513 49989
rect 183547 49961 183575 49989
rect 183609 49961 183637 49989
rect 183671 49961 183699 49989
rect 183485 41147 183513 41175
rect 183547 41147 183575 41175
rect 183609 41147 183637 41175
rect 183671 41147 183699 41175
rect 183485 41085 183513 41113
rect 183547 41085 183575 41113
rect 183609 41085 183637 41113
rect 183671 41085 183699 41113
rect 183485 41023 183513 41051
rect 183547 41023 183575 41051
rect 183609 41023 183637 41051
rect 183671 41023 183699 41051
rect 183485 40961 183513 40989
rect 183547 40961 183575 40989
rect 183609 40961 183637 40989
rect 183671 40961 183699 40989
rect 183485 32147 183513 32175
rect 183547 32147 183575 32175
rect 183609 32147 183637 32175
rect 183671 32147 183699 32175
rect 183485 32085 183513 32113
rect 183547 32085 183575 32113
rect 183609 32085 183637 32113
rect 183671 32085 183699 32113
rect 183485 32023 183513 32051
rect 183547 32023 183575 32051
rect 183609 32023 183637 32051
rect 183671 32023 183699 32051
rect 183485 31961 183513 31989
rect 183547 31961 183575 31989
rect 183609 31961 183637 31989
rect 183671 31961 183699 31989
rect 183485 23147 183513 23175
rect 183547 23147 183575 23175
rect 183609 23147 183637 23175
rect 183671 23147 183699 23175
rect 183485 23085 183513 23113
rect 183547 23085 183575 23113
rect 183609 23085 183637 23113
rect 183671 23085 183699 23113
rect 183485 23023 183513 23051
rect 183547 23023 183575 23051
rect 183609 23023 183637 23051
rect 183671 23023 183699 23051
rect 183485 22961 183513 22989
rect 183547 22961 183575 22989
rect 183609 22961 183637 22989
rect 183671 22961 183699 22989
rect 183485 14147 183513 14175
rect 183547 14147 183575 14175
rect 183609 14147 183637 14175
rect 183671 14147 183699 14175
rect 183485 14085 183513 14113
rect 183547 14085 183575 14113
rect 183609 14085 183637 14113
rect 183671 14085 183699 14113
rect 183485 14023 183513 14051
rect 183547 14023 183575 14051
rect 183609 14023 183637 14051
rect 183671 14023 183699 14051
rect 183485 13961 183513 13989
rect 183547 13961 183575 13989
rect 183609 13961 183637 13989
rect 183671 13961 183699 13989
rect 183485 5147 183513 5175
rect 183547 5147 183575 5175
rect 183609 5147 183637 5175
rect 183671 5147 183699 5175
rect 183485 5085 183513 5113
rect 183547 5085 183575 5113
rect 183609 5085 183637 5113
rect 183671 5085 183699 5113
rect 183485 5023 183513 5051
rect 183547 5023 183575 5051
rect 183609 5023 183637 5051
rect 183671 5023 183699 5051
rect 183485 4961 183513 4989
rect 183547 4961 183575 4989
rect 183609 4961 183637 4989
rect 183671 4961 183699 4989
rect 183485 -588 183513 -560
rect 183547 -588 183575 -560
rect 183609 -588 183637 -560
rect 183671 -588 183699 -560
rect 183485 -650 183513 -622
rect 183547 -650 183575 -622
rect 183609 -650 183637 -622
rect 183671 -650 183699 -622
rect 183485 -712 183513 -684
rect 183547 -712 183575 -684
rect 183609 -712 183637 -684
rect 183671 -712 183699 -684
rect 183485 -774 183513 -746
rect 183547 -774 183575 -746
rect 183609 -774 183637 -746
rect 183671 -774 183699 -746
rect 190625 298578 190653 298606
rect 190687 298578 190715 298606
rect 190749 298578 190777 298606
rect 190811 298578 190839 298606
rect 190625 298516 190653 298544
rect 190687 298516 190715 298544
rect 190749 298516 190777 298544
rect 190811 298516 190839 298544
rect 190625 298454 190653 298482
rect 190687 298454 190715 298482
rect 190749 298454 190777 298482
rect 190811 298454 190839 298482
rect 190625 298392 190653 298420
rect 190687 298392 190715 298420
rect 190749 298392 190777 298420
rect 190811 298392 190839 298420
rect 190625 290147 190653 290175
rect 190687 290147 190715 290175
rect 190749 290147 190777 290175
rect 190811 290147 190839 290175
rect 190625 290085 190653 290113
rect 190687 290085 190715 290113
rect 190749 290085 190777 290113
rect 190811 290085 190839 290113
rect 190625 290023 190653 290051
rect 190687 290023 190715 290051
rect 190749 290023 190777 290051
rect 190811 290023 190839 290051
rect 190625 289961 190653 289989
rect 190687 289961 190715 289989
rect 190749 289961 190777 289989
rect 190811 289961 190839 289989
rect 190625 281147 190653 281175
rect 190687 281147 190715 281175
rect 190749 281147 190777 281175
rect 190811 281147 190839 281175
rect 190625 281085 190653 281113
rect 190687 281085 190715 281113
rect 190749 281085 190777 281113
rect 190811 281085 190839 281113
rect 190625 281023 190653 281051
rect 190687 281023 190715 281051
rect 190749 281023 190777 281051
rect 190811 281023 190839 281051
rect 190625 280961 190653 280989
rect 190687 280961 190715 280989
rect 190749 280961 190777 280989
rect 190811 280961 190839 280989
rect 190625 272147 190653 272175
rect 190687 272147 190715 272175
rect 190749 272147 190777 272175
rect 190811 272147 190839 272175
rect 190625 272085 190653 272113
rect 190687 272085 190715 272113
rect 190749 272085 190777 272113
rect 190811 272085 190839 272113
rect 190625 272023 190653 272051
rect 190687 272023 190715 272051
rect 190749 272023 190777 272051
rect 190811 272023 190839 272051
rect 190625 271961 190653 271989
rect 190687 271961 190715 271989
rect 190749 271961 190777 271989
rect 190811 271961 190839 271989
rect 190625 263147 190653 263175
rect 190687 263147 190715 263175
rect 190749 263147 190777 263175
rect 190811 263147 190839 263175
rect 190625 263085 190653 263113
rect 190687 263085 190715 263113
rect 190749 263085 190777 263113
rect 190811 263085 190839 263113
rect 190625 263023 190653 263051
rect 190687 263023 190715 263051
rect 190749 263023 190777 263051
rect 190811 263023 190839 263051
rect 190625 262961 190653 262989
rect 190687 262961 190715 262989
rect 190749 262961 190777 262989
rect 190811 262961 190839 262989
rect 190625 254147 190653 254175
rect 190687 254147 190715 254175
rect 190749 254147 190777 254175
rect 190811 254147 190839 254175
rect 190625 254085 190653 254113
rect 190687 254085 190715 254113
rect 190749 254085 190777 254113
rect 190811 254085 190839 254113
rect 190625 254023 190653 254051
rect 190687 254023 190715 254051
rect 190749 254023 190777 254051
rect 190811 254023 190839 254051
rect 190625 253961 190653 253989
rect 190687 253961 190715 253989
rect 190749 253961 190777 253989
rect 190811 253961 190839 253989
rect 190625 245147 190653 245175
rect 190687 245147 190715 245175
rect 190749 245147 190777 245175
rect 190811 245147 190839 245175
rect 190625 245085 190653 245113
rect 190687 245085 190715 245113
rect 190749 245085 190777 245113
rect 190811 245085 190839 245113
rect 190625 245023 190653 245051
rect 190687 245023 190715 245051
rect 190749 245023 190777 245051
rect 190811 245023 190839 245051
rect 190625 244961 190653 244989
rect 190687 244961 190715 244989
rect 190749 244961 190777 244989
rect 190811 244961 190839 244989
rect 190625 236147 190653 236175
rect 190687 236147 190715 236175
rect 190749 236147 190777 236175
rect 190811 236147 190839 236175
rect 190625 236085 190653 236113
rect 190687 236085 190715 236113
rect 190749 236085 190777 236113
rect 190811 236085 190839 236113
rect 190625 236023 190653 236051
rect 190687 236023 190715 236051
rect 190749 236023 190777 236051
rect 190811 236023 190839 236051
rect 190625 235961 190653 235989
rect 190687 235961 190715 235989
rect 190749 235961 190777 235989
rect 190811 235961 190839 235989
rect 190625 227147 190653 227175
rect 190687 227147 190715 227175
rect 190749 227147 190777 227175
rect 190811 227147 190839 227175
rect 190625 227085 190653 227113
rect 190687 227085 190715 227113
rect 190749 227085 190777 227113
rect 190811 227085 190839 227113
rect 190625 227023 190653 227051
rect 190687 227023 190715 227051
rect 190749 227023 190777 227051
rect 190811 227023 190839 227051
rect 190625 226961 190653 226989
rect 190687 226961 190715 226989
rect 190749 226961 190777 226989
rect 190811 226961 190839 226989
rect 190625 218147 190653 218175
rect 190687 218147 190715 218175
rect 190749 218147 190777 218175
rect 190811 218147 190839 218175
rect 190625 218085 190653 218113
rect 190687 218085 190715 218113
rect 190749 218085 190777 218113
rect 190811 218085 190839 218113
rect 190625 218023 190653 218051
rect 190687 218023 190715 218051
rect 190749 218023 190777 218051
rect 190811 218023 190839 218051
rect 190625 217961 190653 217989
rect 190687 217961 190715 217989
rect 190749 217961 190777 217989
rect 190811 217961 190839 217989
rect 190625 209147 190653 209175
rect 190687 209147 190715 209175
rect 190749 209147 190777 209175
rect 190811 209147 190839 209175
rect 190625 209085 190653 209113
rect 190687 209085 190715 209113
rect 190749 209085 190777 209113
rect 190811 209085 190839 209113
rect 190625 209023 190653 209051
rect 190687 209023 190715 209051
rect 190749 209023 190777 209051
rect 190811 209023 190839 209051
rect 190625 208961 190653 208989
rect 190687 208961 190715 208989
rect 190749 208961 190777 208989
rect 190811 208961 190839 208989
rect 190625 200147 190653 200175
rect 190687 200147 190715 200175
rect 190749 200147 190777 200175
rect 190811 200147 190839 200175
rect 190625 200085 190653 200113
rect 190687 200085 190715 200113
rect 190749 200085 190777 200113
rect 190811 200085 190839 200113
rect 190625 200023 190653 200051
rect 190687 200023 190715 200051
rect 190749 200023 190777 200051
rect 190811 200023 190839 200051
rect 190625 199961 190653 199989
rect 190687 199961 190715 199989
rect 190749 199961 190777 199989
rect 190811 199961 190839 199989
rect 190625 191147 190653 191175
rect 190687 191147 190715 191175
rect 190749 191147 190777 191175
rect 190811 191147 190839 191175
rect 190625 191085 190653 191113
rect 190687 191085 190715 191113
rect 190749 191085 190777 191113
rect 190811 191085 190839 191113
rect 190625 191023 190653 191051
rect 190687 191023 190715 191051
rect 190749 191023 190777 191051
rect 190811 191023 190839 191051
rect 190625 190961 190653 190989
rect 190687 190961 190715 190989
rect 190749 190961 190777 190989
rect 190811 190961 190839 190989
rect 190625 182147 190653 182175
rect 190687 182147 190715 182175
rect 190749 182147 190777 182175
rect 190811 182147 190839 182175
rect 190625 182085 190653 182113
rect 190687 182085 190715 182113
rect 190749 182085 190777 182113
rect 190811 182085 190839 182113
rect 190625 182023 190653 182051
rect 190687 182023 190715 182051
rect 190749 182023 190777 182051
rect 190811 182023 190839 182051
rect 190625 181961 190653 181989
rect 190687 181961 190715 181989
rect 190749 181961 190777 181989
rect 190811 181961 190839 181989
rect 190625 173147 190653 173175
rect 190687 173147 190715 173175
rect 190749 173147 190777 173175
rect 190811 173147 190839 173175
rect 190625 173085 190653 173113
rect 190687 173085 190715 173113
rect 190749 173085 190777 173113
rect 190811 173085 190839 173113
rect 190625 173023 190653 173051
rect 190687 173023 190715 173051
rect 190749 173023 190777 173051
rect 190811 173023 190839 173051
rect 190625 172961 190653 172989
rect 190687 172961 190715 172989
rect 190749 172961 190777 172989
rect 190811 172961 190839 172989
rect 190625 164147 190653 164175
rect 190687 164147 190715 164175
rect 190749 164147 190777 164175
rect 190811 164147 190839 164175
rect 190625 164085 190653 164113
rect 190687 164085 190715 164113
rect 190749 164085 190777 164113
rect 190811 164085 190839 164113
rect 190625 164023 190653 164051
rect 190687 164023 190715 164051
rect 190749 164023 190777 164051
rect 190811 164023 190839 164051
rect 190625 163961 190653 163989
rect 190687 163961 190715 163989
rect 190749 163961 190777 163989
rect 190811 163961 190839 163989
rect 190625 155147 190653 155175
rect 190687 155147 190715 155175
rect 190749 155147 190777 155175
rect 190811 155147 190839 155175
rect 190625 155085 190653 155113
rect 190687 155085 190715 155113
rect 190749 155085 190777 155113
rect 190811 155085 190839 155113
rect 190625 155023 190653 155051
rect 190687 155023 190715 155051
rect 190749 155023 190777 155051
rect 190811 155023 190839 155051
rect 190625 154961 190653 154989
rect 190687 154961 190715 154989
rect 190749 154961 190777 154989
rect 190811 154961 190839 154989
rect 190625 146147 190653 146175
rect 190687 146147 190715 146175
rect 190749 146147 190777 146175
rect 190811 146147 190839 146175
rect 190625 146085 190653 146113
rect 190687 146085 190715 146113
rect 190749 146085 190777 146113
rect 190811 146085 190839 146113
rect 190625 146023 190653 146051
rect 190687 146023 190715 146051
rect 190749 146023 190777 146051
rect 190811 146023 190839 146051
rect 190625 145961 190653 145989
rect 190687 145961 190715 145989
rect 190749 145961 190777 145989
rect 190811 145961 190839 145989
rect 190625 137147 190653 137175
rect 190687 137147 190715 137175
rect 190749 137147 190777 137175
rect 190811 137147 190839 137175
rect 190625 137085 190653 137113
rect 190687 137085 190715 137113
rect 190749 137085 190777 137113
rect 190811 137085 190839 137113
rect 190625 137023 190653 137051
rect 190687 137023 190715 137051
rect 190749 137023 190777 137051
rect 190811 137023 190839 137051
rect 190625 136961 190653 136989
rect 190687 136961 190715 136989
rect 190749 136961 190777 136989
rect 190811 136961 190839 136989
rect 190625 128147 190653 128175
rect 190687 128147 190715 128175
rect 190749 128147 190777 128175
rect 190811 128147 190839 128175
rect 190625 128085 190653 128113
rect 190687 128085 190715 128113
rect 190749 128085 190777 128113
rect 190811 128085 190839 128113
rect 190625 128023 190653 128051
rect 190687 128023 190715 128051
rect 190749 128023 190777 128051
rect 190811 128023 190839 128051
rect 190625 127961 190653 127989
rect 190687 127961 190715 127989
rect 190749 127961 190777 127989
rect 190811 127961 190839 127989
rect 190625 119147 190653 119175
rect 190687 119147 190715 119175
rect 190749 119147 190777 119175
rect 190811 119147 190839 119175
rect 190625 119085 190653 119113
rect 190687 119085 190715 119113
rect 190749 119085 190777 119113
rect 190811 119085 190839 119113
rect 190625 119023 190653 119051
rect 190687 119023 190715 119051
rect 190749 119023 190777 119051
rect 190811 119023 190839 119051
rect 190625 118961 190653 118989
rect 190687 118961 190715 118989
rect 190749 118961 190777 118989
rect 190811 118961 190839 118989
rect 190625 110147 190653 110175
rect 190687 110147 190715 110175
rect 190749 110147 190777 110175
rect 190811 110147 190839 110175
rect 190625 110085 190653 110113
rect 190687 110085 190715 110113
rect 190749 110085 190777 110113
rect 190811 110085 190839 110113
rect 190625 110023 190653 110051
rect 190687 110023 190715 110051
rect 190749 110023 190777 110051
rect 190811 110023 190839 110051
rect 190625 109961 190653 109989
rect 190687 109961 190715 109989
rect 190749 109961 190777 109989
rect 190811 109961 190839 109989
rect 190625 101147 190653 101175
rect 190687 101147 190715 101175
rect 190749 101147 190777 101175
rect 190811 101147 190839 101175
rect 190625 101085 190653 101113
rect 190687 101085 190715 101113
rect 190749 101085 190777 101113
rect 190811 101085 190839 101113
rect 190625 101023 190653 101051
rect 190687 101023 190715 101051
rect 190749 101023 190777 101051
rect 190811 101023 190839 101051
rect 190625 100961 190653 100989
rect 190687 100961 190715 100989
rect 190749 100961 190777 100989
rect 190811 100961 190839 100989
rect 190625 92147 190653 92175
rect 190687 92147 190715 92175
rect 190749 92147 190777 92175
rect 190811 92147 190839 92175
rect 190625 92085 190653 92113
rect 190687 92085 190715 92113
rect 190749 92085 190777 92113
rect 190811 92085 190839 92113
rect 190625 92023 190653 92051
rect 190687 92023 190715 92051
rect 190749 92023 190777 92051
rect 190811 92023 190839 92051
rect 190625 91961 190653 91989
rect 190687 91961 190715 91989
rect 190749 91961 190777 91989
rect 190811 91961 190839 91989
rect 190625 83147 190653 83175
rect 190687 83147 190715 83175
rect 190749 83147 190777 83175
rect 190811 83147 190839 83175
rect 190625 83085 190653 83113
rect 190687 83085 190715 83113
rect 190749 83085 190777 83113
rect 190811 83085 190839 83113
rect 190625 83023 190653 83051
rect 190687 83023 190715 83051
rect 190749 83023 190777 83051
rect 190811 83023 190839 83051
rect 190625 82961 190653 82989
rect 190687 82961 190715 82989
rect 190749 82961 190777 82989
rect 190811 82961 190839 82989
rect 190625 74147 190653 74175
rect 190687 74147 190715 74175
rect 190749 74147 190777 74175
rect 190811 74147 190839 74175
rect 190625 74085 190653 74113
rect 190687 74085 190715 74113
rect 190749 74085 190777 74113
rect 190811 74085 190839 74113
rect 190625 74023 190653 74051
rect 190687 74023 190715 74051
rect 190749 74023 190777 74051
rect 190811 74023 190839 74051
rect 190625 73961 190653 73989
rect 190687 73961 190715 73989
rect 190749 73961 190777 73989
rect 190811 73961 190839 73989
rect 190625 65147 190653 65175
rect 190687 65147 190715 65175
rect 190749 65147 190777 65175
rect 190811 65147 190839 65175
rect 190625 65085 190653 65113
rect 190687 65085 190715 65113
rect 190749 65085 190777 65113
rect 190811 65085 190839 65113
rect 190625 65023 190653 65051
rect 190687 65023 190715 65051
rect 190749 65023 190777 65051
rect 190811 65023 190839 65051
rect 190625 64961 190653 64989
rect 190687 64961 190715 64989
rect 190749 64961 190777 64989
rect 190811 64961 190839 64989
rect 190625 56147 190653 56175
rect 190687 56147 190715 56175
rect 190749 56147 190777 56175
rect 190811 56147 190839 56175
rect 190625 56085 190653 56113
rect 190687 56085 190715 56113
rect 190749 56085 190777 56113
rect 190811 56085 190839 56113
rect 190625 56023 190653 56051
rect 190687 56023 190715 56051
rect 190749 56023 190777 56051
rect 190811 56023 190839 56051
rect 190625 55961 190653 55989
rect 190687 55961 190715 55989
rect 190749 55961 190777 55989
rect 190811 55961 190839 55989
rect 190625 47147 190653 47175
rect 190687 47147 190715 47175
rect 190749 47147 190777 47175
rect 190811 47147 190839 47175
rect 190625 47085 190653 47113
rect 190687 47085 190715 47113
rect 190749 47085 190777 47113
rect 190811 47085 190839 47113
rect 190625 47023 190653 47051
rect 190687 47023 190715 47051
rect 190749 47023 190777 47051
rect 190811 47023 190839 47051
rect 190625 46961 190653 46989
rect 190687 46961 190715 46989
rect 190749 46961 190777 46989
rect 190811 46961 190839 46989
rect 190625 38147 190653 38175
rect 190687 38147 190715 38175
rect 190749 38147 190777 38175
rect 190811 38147 190839 38175
rect 190625 38085 190653 38113
rect 190687 38085 190715 38113
rect 190749 38085 190777 38113
rect 190811 38085 190839 38113
rect 190625 38023 190653 38051
rect 190687 38023 190715 38051
rect 190749 38023 190777 38051
rect 190811 38023 190839 38051
rect 190625 37961 190653 37989
rect 190687 37961 190715 37989
rect 190749 37961 190777 37989
rect 190811 37961 190839 37989
rect 190625 29147 190653 29175
rect 190687 29147 190715 29175
rect 190749 29147 190777 29175
rect 190811 29147 190839 29175
rect 190625 29085 190653 29113
rect 190687 29085 190715 29113
rect 190749 29085 190777 29113
rect 190811 29085 190839 29113
rect 190625 29023 190653 29051
rect 190687 29023 190715 29051
rect 190749 29023 190777 29051
rect 190811 29023 190839 29051
rect 190625 28961 190653 28989
rect 190687 28961 190715 28989
rect 190749 28961 190777 28989
rect 190811 28961 190839 28989
rect 190625 20147 190653 20175
rect 190687 20147 190715 20175
rect 190749 20147 190777 20175
rect 190811 20147 190839 20175
rect 190625 20085 190653 20113
rect 190687 20085 190715 20113
rect 190749 20085 190777 20113
rect 190811 20085 190839 20113
rect 190625 20023 190653 20051
rect 190687 20023 190715 20051
rect 190749 20023 190777 20051
rect 190811 20023 190839 20051
rect 190625 19961 190653 19989
rect 190687 19961 190715 19989
rect 190749 19961 190777 19989
rect 190811 19961 190839 19989
rect 190625 11147 190653 11175
rect 190687 11147 190715 11175
rect 190749 11147 190777 11175
rect 190811 11147 190839 11175
rect 190625 11085 190653 11113
rect 190687 11085 190715 11113
rect 190749 11085 190777 11113
rect 190811 11085 190839 11113
rect 190625 11023 190653 11051
rect 190687 11023 190715 11051
rect 190749 11023 190777 11051
rect 190811 11023 190839 11051
rect 190625 10961 190653 10989
rect 190687 10961 190715 10989
rect 190749 10961 190777 10989
rect 190811 10961 190839 10989
rect 190625 2147 190653 2175
rect 190687 2147 190715 2175
rect 190749 2147 190777 2175
rect 190811 2147 190839 2175
rect 190625 2085 190653 2113
rect 190687 2085 190715 2113
rect 190749 2085 190777 2113
rect 190811 2085 190839 2113
rect 190625 2023 190653 2051
rect 190687 2023 190715 2051
rect 190749 2023 190777 2051
rect 190811 2023 190839 2051
rect 190625 1961 190653 1989
rect 190687 1961 190715 1989
rect 190749 1961 190777 1989
rect 190811 1961 190839 1989
rect 190625 -108 190653 -80
rect 190687 -108 190715 -80
rect 190749 -108 190777 -80
rect 190811 -108 190839 -80
rect 190625 -170 190653 -142
rect 190687 -170 190715 -142
rect 190749 -170 190777 -142
rect 190811 -170 190839 -142
rect 190625 -232 190653 -204
rect 190687 -232 190715 -204
rect 190749 -232 190777 -204
rect 190811 -232 190839 -204
rect 190625 -294 190653 -266
rect 190687 -294 190715 -266
rect 190749 -294 190777 -266
rect 190811 -294 190839 -266
rect 192485 299058 192513 299086
rect 192547 299058 192575 299086
rect 192609 299058 192637 299086
rect 192671 299058 192699 299086
rect 192485 298996 192513 299024
rect 192547 298996 192575 299024
rect 192609 298996 192637 299024
rect 192671 298996 192699 299024
rect 192485 298934 192513 298962
rect 192547 298934 192575 298962
rect 192609 298934 192637 298962
rect 192671 298934 192699 298962
rect 192485 298872 192513 298900
rect 192547 298872 192575 298900
rect 192609 298872 192637 298900
rect 192671 298872 192699 298900
rect 192485 293147 192513 293175
rect 192547 293147 192575 293175
rect 192609 293147 192637 293175
rect 192671 293147 192699 293175
rect 192485 293085 192513 293113
rect 192547 293085 192575 293113
rect 192609 293085 192637 293113
rect 192671 293085 192699 293113
rect 192485 293023 192513 293051
rect 192547 293023 192575 293051
rect 192609 293023 192637 293051
rect 192671 293023 192699 293051
rect 192485 292961 192513 292989
rect 192547 292961 192575 292989
rect 192609 292961 192637 292989
rect 192671 292961 192699 292989
rect 192485 284147 192513 284175
rect 192547 284147 192575 284175
rect 192609 284147 192637 284175
rect 192671 284147 192699 284175
rect 192485 284085 192513 284113
rect 192547 284085 192575 284113
rect 192609 284085 192637 284113
rect 192671 284085 192699 284113
rect 192485 284023 192513 284051
rect 192547 284023 192575 284051
rect 192609 284023 192637 284051
rect 192671 284023 192699 284051
rect 192485 283961 192513 283989
rect 192547 283961 192575 283989
rect 192609 283961 192637 283989
rect 192671 283961 192699 283989
rect 192485 275147 192513 275175
rect 192547 275147 192575 275175
rect 192609 275147 192637 275175
rect 192671 275147 192699 275175
rect 192485 275085 192513 275113
rect 192547 275085 192575 275113
rect 192609 275085 192637 275113
rect 192671 275085 192699 275113
rect 192485 275023 192513 275051
rect 192547 275023 192575 275051
rect 192609 275023 192637 275051
rect 192671 275023 192699 275051
rect 192485 274961 192513 274989
rect 192547 274961 192575 274989
rect 192609 274961 192637 274989
rect 192671 274961 192699 274989
rect 192485 266147 192513 266175
rect 192547 266147 192575 266175
rect 192609 266147 192637 266175
rect 192671 266147 192699 266175
rect 192485 266085 192513 266113
rect 192547 266085 192575 266113
rect 192609 266085 192637 266113
rect 192671 266085 192699 266113
rect 192485 266023 192513 266051
rect 192547 266023 192575 266051
rect 192609 266023 192637 266051
rect 192671 266023 192699 266051
rect 192485 265961 192513 265989
rect 192547 265961 192575 265989
rect 192609 265961 192637 265989
rect 192671 265961 192699 265989
rect 192485 257147 192513 257175
rect 192547 257147 192575 257175
rect 192609 257147 192637 257175
rect 192671 257147 192699 257175
rect 192485 257085 192513 257113
rect 192547 257085 192575 257113
rect 192609 257085 192637 257113
rect 192671 257085 192699 257113
rect 192485 257023 192513 257051
rect 192547 257023 192575 257051
rect 192609 257023 192637 257051
rect 192671 257023 192699 257051
rect 192485 256961 192513 256989
rect 192547 256961 192575 256989
rect 192609 256961 192637 256989
rect 192671 256961 192699 256989
rect 192485 248147 192513 248175
rect 192547 248147 192575 248175
rect 192609 248147 192637 248175
rect 192671 248147 192699 248175
rect 192485 248085 192513 248113
rect 192547 248085 192575 248113
rect 192609 248085 192637 248113
rect 192671 248085 192699 248113
rect 192485 248023 192513 248051
rect 192547 248023 192575 248051
rect 192609 248023 192637 248051
rect 192671 248023 192699 248051
rect 192485 247961 192513 247989
rect 192547 247961 192575 247989
rect 192609 247961 192637 247989
rect 192671 247961 192699 247989
rect 192485 239147 192513 239175
rect 192547 239147 192575 239175
rect 192609 239147 192637 239175
rect 192671 239147 192699 239175
rect 192485 239085 192513 239113
rect 192547 239085 192575 239113
rect 192609 239085 192637 239113
rect 192671 239085 192699 239113
rect 192485 239023 192513 239051
rect 192547 239023 192575 239051
rect 192609 239023 192637 239051
rect 192671 239023 192699 239051
rect 192485 238961 192513 238989
rect 192547 238961 192575 238989
rect 192609 238961 192637 238989
rect 192671 238961 192699 238989
rect 192485 230147 192513 230175
rect 192547 230147 192575 230175
rect 192609 230147 192637 230175
rect 192671 230147 192699 230175
rect 192485 230085 192513 230113
rect 192547 230085 192575 230113
rect 192609 230085 192637 230113
rect 192671 230085 192699 230113
rect 192485 230023 192513 230051
rect 192547 230023 192575 230051
rect 192609 230023 192637 230051
rect 192671 230023 192699 230051
rect 192485 229961 192513 229989
rect 192547 229961 192575 229989
rect 192609 229961 192637 229989
rect 192671 229961 192699 229989
rect 192485 221147 192513 221175
rect 192547 221147 192575 221175
rect 192609 221147 192637 221175
rect 192671 221147 192699 221175
rect 192485 221085 192513 221113
rect 192547 221085 192575 221113
rect 192609 221085 192637 221113
rect 192671 221085 192699 221113
rect 192485 221023 192513 221051
rect 192547 221023 192575 221051
rect 192609 221023 192637 221051
rect 192671 221023 192699 221051
rect 192485 220961 192513 220989
rect 192547 220961 192575 220989
rect 192609 220961 192637 220989
rect 192671 220961 192699 220989
rect 192485 212147 192513 212175
rect 192547 212147 192575 212175
rect 192609 212147 192637 212175
rect 192671 212147 192699 212175
rect 192485 212085 192513 212113
rect 192547 212085 192575 212113
rect 192609 212085 192637 212113
rect 192671 212085 192699 212113
rect 192485 212023 192513 212051
rect 192547 212023 192575 212051
rect 192609 212023 192637 212051
rect 192671 212023 192699 212051
rect 192485 211961 192513 211989
rect 192547 211961 192575 211989
rect 192609 211961 192637 211989
rect 192671 211961 192699 211989
rect 192485 203147 192513 203175
rect 192547 203147 192575 203175
rect 192609 203147 192637 203175
rect 192671 203147 192699 203175
rect 192485 203085 192513 203113
rect 192547 203085 192575 203113
rect 192609 203085 192637 203113
rect 192671 203085 192699 203113
rect 192485 203023 192513 203051
rect 192547 203023 192575 203051
rect 192609 203023 192637 203051
rect 192671 203023 192699 203051
rect 192485 202961 192513 202989
rect 192547 202961 192575 202989
rect 192609 202961 192637 202989
rect 192671 202961 192699 202989
rect 192485 194147 192513 194175
rect 192547 194147 192575 194175
rect 192609 194147 192637 194175
rect 192671 194147 192699 194175
rect 192485 194085 192513 194113
rect 192547 194085 192575 194113
rect 192609 194085 192637 194113
rect 192671 194085 192699 194113
rect 192485 194023 192513 194051
rect 192547 194023 192575 194051
rect 192609 194023 192637 194051
rect 192671 194023 192699 194051
rect 192485 193961 192513 193989
rect 192547 193961 192575 193989
rect 192609 193961 192637 193989
rect 192671 193961 192699 193989
rect 192485 185147 192513 185175
rect 192547 185147 192575 185175
rect 192609 185147 192637 185175
rect 192671 185147 192699 185175
rect 192485 185085 192513 185113
rect 192547 185085 192575 185113
rect 192609 185085 192637 185113
rect 192671 185085 192699 185113
rect 192485 185023 192513 185051
rect 192547 185023 192575 185051
rect 192609 185023 192637 185051
rect 192671 185023 192699 185051
rect 192485 184961 192513 184989
rect 192547 184961 192575 184989
rect 192609 184961 192637 184989
rect 192671 184961 192699 184989
rect 192485 176147 192513 176175
rect 192547 176147 192575 176175
rect 192609 176147 192637 176175
rect 192671 176147 192699 176175
rect 192485 176085 192513 176113
rect 192547 176085 192575 176113
rect 192609 176085 192637 176113
rect 192671 176085 192699 176113
rect 192485 176023 192513 176051
rect 192547 176023 192575 176051
rect 192609 176023 192637 176051
rect 192671 176023 192699 176051
rect 192485 175961 192513 175989
rect 192547 175961 192575 175989
rect 192609 175961 192637 175989
rect 192671 175961 192699 175989
rect 192485 167147 192513 167175
rect 192547 167147 192575 167175
rect 192609 167147 192637 167175
rect 192671 167147 192699 167175
rect 192485 167085 192513 167113
rect 192547 167085 192575 167113
rect 192609 167085 192637 167113
rect 192671 167085 192699 167113
rect 192485 167023 192513 167051
rect 192547 167023 192575 167051
rect 192609 167023 192637 167051
rect 192671 167023 192699 167051
rect 192485 166961 192513 166989
rect 192547 166961 192575 166989
rect 192609 166961 192637 166989
rect 192671 166961 192699 166989
rect 192485 158147 192513 158175
rect 192547 158147 192575 158175
rect 192609 158147 192637 158175
rect 192671 158147 192699 158175
rect 192485 158085 192513 158113
rect 192547 158085 192575 158113
rect 192609 158085 192637 158113
rect 192671 158085 192699 158113
rect 192485 158023 192513 158051
rect 192547 158023 192575 158051
rect 192609 158023 192637 158051
rect 192671 158023 192699 158051
rect 192485 157961 192513 157989
rect 192547 157961 192575 157989
rect 192609 157961 192637 157989
rect 192671 157961 192699 157989
rect 192485 149147 192513 149175
rect 192547 149147 192575 149175
rect 192609 149147 192637 149175
rect 192671 149147 192699 149175
rect 192485 149085 192513 149113
rect 192547 149085 192575 149113
rect 192609 149085 192637 149113
rect 192671 149085 192699 149113
rect 192485 149023 192513 149051
rect 192547 149023 192575 149051
rect 192609 149023 192637 149051
rect 192671 149023 192699 149051
rect 192485 148961 192513 148989
rect 192547 148961 192575 148989
rect 192609 148961 192637 148989
rect 192671 148961 192699 148989
rect 192485 140147 192513 140175
rect 192547 140147 192575 140175
rect 192609 140147 192637 140175
rect 192671 140147 192699 140175
rect 192485 140085 192513 140113
rect 192547 140085 192575 140113
rect 192609 140085 192637 140113
rect 192671 140085 192699 140113
rect 192485 140023 192513 140051
rect 192547 140023 192575 140051
rect 192609 140023 192637 140051
rect 192671 140023 192699 140051
rect 192485 139961 192513 139989
rect 192547 139961 192575 139989
rect 192609 139961 192637 139989
rect 192671 139961 192699 139989
rect 192485 131147 192513 131175
rect 192547 131147 192575 131175
rect 192609 131147 192637 131175
rect 192671 131147 192699 131175
rect 192485 131085 192513 131113
rect 192547 131085 192575 131113
rect 192609 131085 192637 131113
rect 192671 131085 192699 131113
rect 192485 131023 192513 131051
rect 192547 131023 192575 131051
rect 192609 131023 192637 131051
rect 192671 131023 192699 131051
rect 192485 130961 192513 130989
rect 192547 130961 192575 130989
rect 192609 130961 192637 130989
rect 192671 130961 192699 130989
rect 192485 122147 192513 122175
rect 192547 122147 192575 122175
rect 192609 122147 192637 122175
rect 192671 122147 192699 122175
rect 192485 122085 192513 122113
rect 192547 122085 192575 122113
rect 192609 122085 192637 122113
rect 192671 122085 192699 122113
rect 192485 122023 192513 122051
rect 192547 122023 192575 122051
rect 192609 122023 192637 122051
rect 192671 122023 192699 122051
rect 192485 121961 192513 121989
rect 192547 121961 192575 121989
rect 192609 121961 192637 121989
rect 192671 121961 192699 121989
rect 192485 113147 192513 113175
rect 192547 113147 192575 113175
rect 192609 113147 192637 113175
rect 192671 113147 192699 113175
rect 192485 113085 192513 113113
rect 192547 113085 192575 113113
rect 192609 113085 192637 113113
rect 192671 113085 192699 113113
rect 192485 113023 192513 113051
rect 192547 113023 192575 113051
rect 192609 113023 192637 113051
rect 192671 113023 192699 113051
rect 192485 112961 192513 112989
rect 192547 112961 192575 112989
rect 192609 112961 192637 112989
rect 192671 112961 192699 112989
rect 192485 104147 192513 104175
rect 192547 104147 192575 104175
rect 192609 104147 192637 104175
rect 192671 104147 192699 104175
rect 192485 104085 192513 104113
rect 192547 104085 192575 104113
rect 192609 104085 192637 104113
rect 192671 104085 192699 104113
rect 192485 104023 192513 104051
rect 192547 104023 192575 104051
rect 192609 104023 192637 104051
rect 192671 104023 192699 104051
rect 192485 103961 192513 103989
rect 192547 103961 192575 103989
rect 192609 103961 192637 103989
rect 192671 103961 192699 103989
rect 192485 95147 192513 95175
rect 192547 95147 192575 95175
rect 192609 95147 192637 95175
rect 192671 95147 192699 95175
rect 192485 95085 192513 95113
rect 192547 95085 192575 95113
rect 192609 95085 192637 95113
rect 192671 95085 192699 95113
rect 192485 95023 192513 95051
rect 192547 95023 192575 95051
rect 192609 95023 192637 95051
rect 192671 95023 192699 95051
rect 192485 94961 192513 94989
rect 192547 94961 192575 94989
rect 192609 94961 192637 94989
rect 192671 94961 192699 94989
rect 192485 86147 192513 86175
rect 192547 86147 192575 86175
rect 192609 86147 192637 86175
rect 192671 86147 192699 86175
rect 192485 86085 192513 86113
rect 192547 86085 192575 86113
rect 192609 86085 192637 86113
rect 192671 86085 192699 86113
rect 192485 86023 192513 86051
rect 192547 86023 192575 86051
rect 192609 86023 192637 86051
rect 192671 86023 192699 86051
rect 192485 85961 192513 85989
rect 192547 85961 192575 85989
rect 192609 85961 192637 85989
rect 192671 85961 192699 85989
rect 192485 77147 192513 77175
rect 192547 77147 192575 77175
rect 192609 77147 192637 77175
rect 192671 77147 192699 77175
rect 192485 77085 192513 77113
rect 192547 77085 192575 77113
rect 192609 77085 192637 77113
rect 192671 77085 192699 77113
rect 192485 77023 192513 77051
rect 192547 77023 192575 77051
rect 192609 77023 192637 77051
rect 192671 77023 192699 77051
rect 192485 76961 192513 76989
rect 192547 76961 192575 76989
rect 192609 76961 192637 76989
rect 192671 76961 192699 76989
rect 192485 68147 192513 68175
rect 192547 68147 192575 68175
rect 192609 68147 192637 68175
rect 192671 68147 192699 68175
rect 192485 68085 192513 68113
rect 192547 68085 192575 68113
rect 192609 68085 192637 68113
rect 192671 68085 192699 68113
rect 192485 68023 192513 68051
rect 192547 68023 192575 68051
rect 192609 68023 192637 68051
rect 192671 68023 192699 68051
rect 192485 67961 192513 67989
rect 192547 67961 192575 67989
rect 192609 67961 192637 67989
rect 192671 67961 192699 67989
rect 192485 59147 192513 59175
rect 192547 59147 192575 59175
rect 192609 59147 192637 59175
rect 192671 59147 192699 59175
rect 192485 59085 192513 59113
rect 192547 59085 192575 59113
rect 192609 59085 192637 59113
rect 192671 59085 192699 59113
rect 192485 59023 192513 59051
rect 192547 59023 192575 59051
rect 192609 59023 192637 59051
rect 192671 59023 192699 59051
rect 192485 58961 192513 58989
rect 192547 58961 192575 58989
rect 192609 58961 192637 58989
rect 192671 58961 192699 58989
rect 192485 50147 192513 50175
rect 192547 50147 192575 50175
rect 192609 50147 192637 50175
rect 192671 50147 192699 50175
rect 192485 50085 192513 50113
rect 192547 50085 192575 50113
rect 192609 50085 192637 50113
rect 192671 50085 192699 50113
rect 192485 50023 192513 50051
rect 192547 50023 192575 50051
rect 192609 50023 192637 50051
rect 192671 50023 192699 50051
rect 192485 49961 192513 49989
rect 192547 49961 192575 49989
rect 192609 49961 192637 49989
rect 192671 49961 192699 49989
rect 192485 41147 192513 41175
rect 192547 41147 192575 41175
rect 192609 41147 192637 41175
rect 192671 41147 192699 41175
rect 192485 41085 192513 41113
rect 192547 41085 192575 41113
rect 192609 41085 192637 41113
rect 192671 41085 192699 41113
rect 192485 41023 192513 41051
rect 192547 41023 192575 41051
rect 192609 41023 192637 41051
rect 192671 41023 192699 41051
rect 192485 40961 192513 40989
rect 192547 40961 192575 40989
rect 192609 40961 192637 40989
rect 192671 40961 192699 40989
rect 192485 32147 192513 32175
rect 192547 32147 192575 32175
rect 192609 32147 192637 32175
rect 192671 32147 192699 32175
rect 192485 32085 192513 32113
rect 192547 32085 192575 32113
rect 192609 32085 192637 32113
rect 192671 32085 192699 32113
rect 192485 32023 192513 32051
rect 192547 32023 192575 32051
rect 192609 32023 192637 32051
rect 192671 32023 192699 32051
rect 192485 31961 192513 31989
rect 192547 31961 192575 31989
rect 192609 31961 192637 31989
rect 192671 31961 192699 31989
rect 192485 23147 192513 23175
rect 192547 23147 192575 23175
rect 192609 23147 192637 23175
rect 192671 23147 192699 23175
rect 192485 23085 192513 23113
rect 192547 23085 192575 23113
rect 192609 23085 192637 23113
rect 192671 23085 192699 23113
rect 192485 23023 192513 23051
rect 192547 23023 192575 23051
rect 192609 23023 192637 23051
rect 192671 23023 192699 23051
rect 192485 22961 192513 22989
rect 192547 22961 192575 22989
rect 192609 22961 192637 22989
rect 192671 22961 192699 22989
rect 192485 14147 192513 14175
rect 192547 14147 192575 14175
rect 192609 14147 192637 14175
rect 192671 14147 192699 14175
rect 192485 14085 192513 14113
rect 192547 14085 192575 14113
rect 192609 14085 192637 14113
rect 192671 14085 192699 14113
rect 192485 14023 192513 14051
rect 192547 14023 192575 14051
rect 192609 14023 192637 14051
rect 192671 14023 192699 14051
rect 192485 13961 192513 13989
rect 192547 13961 192575 13989
rect 192609 13961 192637 13989
rect 192671 13961 192699 13989
rect 192485 5147 192513 5175
rect 192547 5147 192575 5175
rect 192609 5147 192637 5175
rect 192671 5147 192699 5175
rect 192485 5085 192513 5113
rect 192547 5085 192575 5113
rect 192609 5085 192637 5113
rect 192671 5085 192699 5113
rect 192485 5023 192513 5051
rect 192547 5023 192575 5051
rect 192609 5023 192637 5051
rect 192671 5023 192699 5051
rect 192485 4961 192513 4989
rect 192547 4961 192575 4989
rect 192609 4961 192637 4989
rect 192671 4961 192699 4989
rect 192485 -588 192513 -560
rect 192547 -588 192575 -560
rect 192609 -588 192637 -560
rect 192671 -588 192699 -560
rect 192485 -650 192513 -622
rect 192547 -650 192575 -622
rect 192609 -650 192637 -622
rect 192671 -650 192699 -622
rect 192485 -712 192513 -684
rect 192547 -712 192575 -684
rect 192609 -712 192637 -684
rect 192671 -712 192699 -684
rect 192485 -774 192513 -746
rect 192547 -774 192575 -746
rect 192609 -774 192637 -746
rect 192671 -774 192699 -746
rect 199625 298578 199653 298606
rect 199687 298578 199715 298606
rect 199749 298578 199777 298606
rect 199811 298578 199839 298606
rect 199625 298516 199653 298544
rect 199687 298516 199715 298544
rect 199749 298516 199777 298544
rect 199811 298516 199839 298544
rect 199625 298454 199653 298482
rect 199687 298454 199715 298482
rect 199749 298454 199777 298482
rect 199811 298454 199839 298482
rect 199625 298392 199653 298420
rect 199687 298392 199715 298420
rect 199749 298392 199777 298420
rect 199811 298392 199839 298420
rect 199625 290147 199653 290175
rect 199687 290147 199715 290175
rect 199749 290147 199777 290175
rect 199811 290147 199839 290175
rect 199625 290085 199653 290113
rect 199687 290085 199715 290113
rect 199749 290085 199777 290113
rect 199811 290085 199839 290113
rect 199625 290023 199653 290051
rect 199687 290023 199715 290051
rect 199749 290023 199777 290051
rect 199811 290023 199839 290051
rect 199625 289961 199653 289989
rect 199687 289961 199715 289989
rect 199749 289961 199777 289989
rect 199811 289961 199839 289989
rect 199625 281147 199653 281175
rect 199687 281147 199715 281175
rect 199749 281147 199777 281175
rect 199811 281147 199839 281175
rect 199625 281085 199653 281113
rect 199687 281085 199715 281113
rect 199749 281085 199777 281113
rect 199811 281085 199839 281113
rect 199625 281023 199653 281051
rect 199687 281023 199715 281051
rect 199749 281023 199777 281051
rect 199811 281023 199839 281051
rect 199625 280961 199653 280989
rect 199687 280961 199715 280989
rect 199749 280961 199777 280989
rect 199811 280961 199839 280989
rect 199625 272147 199653 272175
rect 199687 272147 199715 272175
rect 199749 272147 199777 272175
rect 199811 272147 199839 272175
rect 199625 272085 199653 272113
rect 199687 272085 199715 272113
rect 199749 272085 199777 272113
rect 199811 272085 199839 272113
rect 199625 272023 199653 272051
rect 199687 272023 199715 272051
rect 199749 272023 199777 272051
rect 199811 272023 199839 272051
rect 199625 271961 199653 271989
rect 199687 271961 199715 271989
rect 199749 271961 199777 271989
rect 199811 271961 199839 271989
rect 199625 263147 199653 263175
rect 199687 263147 199715 263175
rect 199749 263147 199777 263175
rect 199811 263147 199839 263175
rect 199625 263085 199653 263113
rect 199687 263085 199715 263113
rect 199749 263085 199777 263113
rect 199811 263085 199839 263113
rect 199625 263023 199653 263051
rect 199687 263023 199715 263051
rect 199749 263023 199777 263051
rect 199811 263023 199839 263051
rect 199625 262961 199653 262989
rect 199687 262961 199715 262989
rect 199749 262961 199777 262989
rect 199811 262961 199839 262989
rect 199625 254147 199653 254175
rect 199687 254147 199715 254175
rect 199749 254147 199777 254175
rect 199811 254147 199839 254175
rect 199625 254085 199653 254113
rect 199687 254085 199715 254113
rect 199749 254085 199777 254113
rect 199811 254085 199839 254113
rect 199625 254023 199653 254051
rect 199687 254023 199715 254051
rect 199749 254023 199777 254051
rect 199811 254023 199839 254051
rect 199625 253961 199653 253989
rect 199687 253961 199715 253989
rect 199749 253961 199777 253989
rect 199811 253961 199839 253989
rect 199625 245147 199653 245175
rect 199687 245147 199715 245175
rect 199749 245147 199777 245175
rect 199811 245147 199839 245175
rect 199625 245085 199653 245113
rect 199687 245085 199715 245113
rect 199749 245085 199777 245113
rect 199811 245085 199839 245113
rect 199625 245023 199653 245051
rect 199687 245023 199715 245051
rect 199749 245023 199777 245051
rect 199811 245023 199839 245051
rect 199625 244961 199653 244989
rect 199687 244961 199715 244989
rect 199749 244961 199777 244989
rect 199811 244961 199839 244989
rect 199625 236147 199653 236175
rect 199687 236147 199715 236175
rect 199749 236147 199777 236175
rect 199811 236147 199839 236175
rect 199625 236085 199653 236113
rect 199687 236085 199715 236113
rect 199749 236085 199777 236113
rect 199811 236085 199839 236113
rect 199625 236023 199653 236051
rect 199687 236023 199715 236051
rect 199749 236023 199777 236051
rect 199811 236023 199839 236051
rect 199625 235961 199653 235989
rect 199687 235961 199715 235989
rect 199749 235961 199777 235989
rect 199811 235961 199839 235989
rect 199625 227147 199653 227175
rect 199687 227147 199715 227175
rect 199749 227147 199777 227175
rect 199811 227147 199839 227175
rect 199625 227085 199653 227113
rect 199687 227085 199715 227113
rect 199749 227085 199777 227113
rect 199811 227085 199839 227113
rect 199625 227023 199653 227051
rect 199687 227023 199715 227051
rect 199749 227023 199777 227051
rect 199811 227023 199839 227051
rect 199625 226961 199653 226989
rect 199687 226961 199715 226989
rect 199749 226961 199777 226989
rect 199811 226961 199839 226989
rect 199625 218147 199653 218175
rect 199687 218147 199715 218175
rect 199749 218147 199777 218175
rect 199811 218147 199839 218175
rect 199625 218085 199653 218113
rect 199687 218085 199715 218113
rect 199749 218085 199777 218113
rect 199811 218085 199839 218113
rect 199625 218023 199653 218051
rect 199687 218023 199715 218051
rect 199749 218023 199777 218051
rect 199811 218023 199839 218051
rect 199625 217961 199653 217989
rect 199687 217961 199715 217989
rect 199749 217961 199777 217989
rect 199811 217961 199839 217989
rect 199625 209147 199653 209175
rect 199687 209147 199715 209175
rect 199749 209147 199777 209175
rect 199811 209147 199839 209175
rect 199625 209085 199653 209113
rect 199687 209085 199715 209113
rect 199749 209085 199777 209113
rect 199811 209085 199839 209113
rect 199625 209023 199653 209051
rect 199687 209023 199715 209051
rect 199749 209023 199777 209051
rect 199811 209023 199839 209051
rect 199625 208961 199653 208989
rect 199687 208961 199715 208989
rect 199749 208961 199777 208989
rect 199811 208961 199839 208989
rect 199625 200147 199653 200175
rect 199687 200147 199715 200175
rect 199749 200147 199777 200175
rect 199811 200147 199839 200175
rect 199625 200085 199653 200113
rect 199687 200085 199715 200113
rect 199749 200085 199777 200113
rect 199811 200085 199839 200113
rect 199625 200023 199653 200051
rect 199687 200023 199715 200051
rect 199749 200023 199777 200051
rect 199811 200023 199839 200051
rect 199625 199961 199653 199989
rect 199687 199961 199715 199989
rect 199749 199961 199777 199989
rect 199811 199961 199839 199989
rect 199625 191147 199653 191175
rect 199687 191147 199715 191175
rect 199749 191147 199777 191175
rect 199811 191147 199839 191175
rect 199625 191085 199653 191113
rect 199687 191085 199715 191113
rect 199749 191085 199777 191113
rect 199811 191085 199839 191113
rect 199625 191023 199653 191051
rect 199687 191023 199715 191051
rect 199749 191023 199777 191051
rect 199811 191023 199839 191051
rect 199625 190961 199653 190989
rect 199687 190961 199715 190989
rect 199749 190961 199777 190989
rect 199811 190961 199839 190989
rect 199625 182147 199653 182175
rect 199687 182147 199715 182175
rect 199749 182147 199777 182175
rect 199811 182147 199839 182175
rect 199625 182085 199653 182113
rect 199687 182085 199715 182113
rect 199749 182085 199777 182113
rect 199811 182085 199839 182113
rect 199625 182023 199653 182051
rect 199687 182023 199715 182051
rect 199749 182023 199777 182051
rect 199811 182023 199839 182051
rect 199625 181961 199653 181989
rect 199687 181961 199715 181989
rect 199749 181961 199777 181989
rect 199811 181961 199839 181989
rect 199625 173147 199653 173175
rect 199687 173147 199715 173175
rect 199749 173147 199777 173175
rect 199811 173147 199839 173175
rect 199625 173085 199653 173113
rect 199687 173085 199715 173113
rect 199749 173085 199777 173113
rect 199811 173085 199839 173113
rect 199625 173023 199653 173051
rect 199687 173023 199715 173051
rect 199749 173023 199777 173051
rect 199811 173023 199839 173051
rect 199625 172961 199653 172989
rect 199687 172961 199715 172989
rect 199749 172961 199777 172989
rect 199811 172961 199839 172989
rect 199625 164147 199653 164175
rect 199687 164147 199715 164175
rect 199749 164147 199777 164175
rect 199811 164147 199839 164175
rect 199625 164085 199653 164113
rect 199687 164085 199715 164113
rect 199749 164085 199777 164113
rect 199811 164085 199839 164113
rect 199625 164023 199653 164051
rect 199687 164023 199715 164051
rect 199749 164023 199777 164051
rect 199811 164023 199839 164051
rect 199625 163961 199653 163989
rect 199687 163961 199715 163989
rect 199749 163961 199777 163989
rect 199811 163961 199839 163989
rect 199625 155147 199653 155175
rect 199687 155147 199715 155175
rect 199749 155147 199777 155175
rect 199811 155147 199839 155175
rect 199625 155085 199653 155113
rect 199687 155085 199715 155113
rect 199749 155085 199777 155113
rect 199811 155085 199839 155113
rect 199625 155023 199653 155051
rect 199687 155023 199715 155051
rect 199749 155023 199777 155051
rect 199811 155023 199839 155051
rect 199625 154961 199653 154989
rect 199687 154961 199715 154989
rect 199749 154961 199777 154989
rect 199811 154961 199839 154989
rect 199625 146147 199653 146175
rect 199687 146147 199715 146175
rect 199749 146147 199777 146175
rect 199811 146147 199839 146175
rect 199625 146085 199653 146113
rect 199687 146085 199715 146113
rect 199749 146085 199777 146113
rect 199811 146085 199839 146113
rect 199625 146023 199653 146051
rect 199687 146023 199715 146051
rect 199749 146023 199777 146051
rect 199811 146023 199839 146051
rect 199625 145961 199653 145989
rect 199687 145961 199715 145989
rect 199749 145961 199777 145989
rect 199811 145961 199839 145989
rect 199625 137147 199653 137175
rect 199687 137147 199715 137175
rect 199749 137147 199777 137175
rect 199811 137147 199839 137175
rect 199625 137085 199653 137113
rect 199687 137085 199715 137113
rect 199749 137085 199777 137113
rect 199811 137085 199839 137113
rect 199625 137023 199653 137051
rect 199687 137023 199715 137051
rect 199749 137023 199777 137051
rect 199811 137023 199839 137051
rect 199625 136961 199653 136989
rect 199687 136961 199715 136989
rect 199749 136961 199777 136989
rect 199811 136961 199839 136989
rect 199625 128147 199653 128175
rect 199687 128147 199715 128175
rect 199749 128147 199777 128175
rect 199811 128147 199839 128175
rect 199625 128085 199653 128113
rect 199687 128085 199715 128113
rect 199749 128085 199777 128113
rect 199811 128085 199839 128113
rect 199625 128023 199653 128051
rect 199687 128023 199715 128051
rect 199749 128023 199777 128051
rect 199811 128023 199839 128051
rect 199625 127961 199653 127989
rect 199687 127961 199715 127989
rect 199749 127961 199777 127989
rect 199811 127961 199839 127989
rect 199625 119147 199653 119175
rect 199687 119147 199715 119175
rect 199749 119147 199777 119175
rect 199811 119147 199839 119175
rect 199625 119085 199653 119113
rect 199687 119085 199715 119113
rect 199749 119085 199777 119113
rect 199811 119085 199839 119113
rect 199625 119023 199653 119051
rect 199687 119023 199715 119051
rect 199749 119023 199777 119051
rect 199811 119023 199839 119051
rect 199625 118961 199653 118989
rect 199687 118961 199715 118989
rect 199749 118961 199777 118989
rect 199811 118961 199839 118989
rect 199625 110147 199653 110175
rect 199687 110147 199715 110175
rect 199749 110147 199777 110175
rect 199811 110147 199839 110175
rect 199625 110085 199653 110113
rect 199687 110085 199715 110113
rect 199749 110085 199777 110113
rect 199811 110085 199839 110113
rect 199625 110023 199653 110051
rect 199687 110023 199715 110051
rect 199749 110023 199777 110051
rect 199811 110023 199839 110051
rect 199625 109961 199653 109989
rect 199687 109961 199715 109989
rect 199749 109961 199777 109989
rect 199811 109961 199839 109989
rect 199625 101147 199653 101175
rect 199687 101147 199715 101175
rect 199749 101147 199777 101175
rect 199811 101147 199839 101175
rect 199625 101085 199653 101113
rect 199687 101085 199715 101113
rect 199749 101085 199777 101113
rect 199811 101085 199839 101113
rect 199625 101023 199653 101051
rect 199687 101023 199715 101051
rect 199749 101023 199777 101051
rect 199811 101023 199839 101051
rect 199625 100961 199653 100989
rect 199687 100961 199715 100989
rect 199749 100961 199777 100989
rect 199811 100961 199839 100989
rect 199625 92147 199653 92175
rect 199687 92147 199715 92175
rect 199749 92147 199777 92175
rect 199811 92147 199839 92175
rect 199625 92085 199653 92113
rect 199687 92085 199715 92113
rect 199749 92085 199777 92113
rect 199811 92085 199839 92113
rect 199625 92023 199653 92051
rect 199687 92023 199715 92051
rect 199749 92023 199777 92051
rect 199811 92023 199839 92051
rect 199625 91961 199653 91989
rect 199687 91961 199715 91989
rect 199749 91961 199777 91989
rect 199811 91961 199839 91989
rect 199625 83147 199653 83175
rect 199687 83147 199715 83175
rect 199749 83147 199777 83175
rect 199811 83147 199839 83175
rect 199625 83085 199653 83113
rect 199687 83085 199715 83113
rect 199749 83085 199777 83113
rect 199811 83085 199839 83113
rect 199625 83023 199653 83051
rect 199687 83023 199715 83051
rect 199749 83023 199777 83051
rect 199811 83023 199839 83051
rect 199625 82961 199653 82989
rect 199687 82961 199715 82989
rect 199749 82961 199777 82989
rect 199811 82961 199839 82989
rect 199625 74147 199653 74175
rect 199687 74147 199715 74175
rect 199749 74147 199777 74175
rect 199811 74147 199839 74175
rect 199625 74085 199653 74113
rect 199687 74085 199715 74113
rect 199749 74085 199777 74113
rect 199811 74085 199839 74113
rect 199625 74023 199653 74051
rect 199687 74023 199715 74051
rect 199749 74023 199777 74051
rect 199811 74023 199839 74051
rect 199625 73961 199653 73989
rect 199687 73961 199715 73989
rect 199749 73961 199777 73989
rect 199811 73961 199839 73989
rect 199625 65147 199653 65175
rect 199687 65147 199715 65175
rect 199749 65147 199777 65175
rect 199811 65147 199839 65175
rect 199625 65085 199653 65113
rect 199687 65085 199715 65113
rect 199749 65085 199777 65113
rect 199811 65085 199839 65113
rect 199625 65023 199653 65051
rect 199687 65023 199715 65051
rect 199749 65023 199777 65051
rect 199811 65023 199839 65051
rect 199625 64961 199653 64989
rect 199687 64961 199715 64989
rect 199749 64961 199777 64989
rect 199811 64961 199839 64989
rect 199625 56147 199653 56175
rect 199687 56147 199715 56175
rect 199749 56147 199777 56175
rect 199811 56147 199839 56175
rect 199625 56085 199653 56113
rect 199687 56085 199715 56113
rect 199749 56085 199777 56113
rect 199811 56085 199839 56113
rect 199625 56023 199653 56051
rect 199687 56023 199715 56051
rect 199749 56023 199777 56051
rect 199811 56023 199839 56051
rect 199625 55961 199653 55989
rect 199687 55961 199715 55989
rect 199749 55961 199777 55989
rect 199811 55961 199839 55989
rect 199625 47147 199653 47175
rect 199687 47147 199715 47175
rect 199749 47147 199777 47175
rect 199811 47147 199839 47175
rect 199625 47085 199653 47113
rect 199687 47085 199715 47113
rect 199749 47085 199777 47113
rect 199811 47085 199839 47113
rect 199625 47023 199653 47051
rect 199687 47023 199715 47051
rect 199749 47023 199777 47051
rect 199811 47023 199839 47051
rect 199625 46961 199653 46989
rect 199687 46961 199715 46989
rect 199749 46961 199777 46989
rect 199811 46961 199839 46989
rect 199625 38147 199653 38175
rect 199687 38147 199715 38175
rect 199749 38147 199777 38175
rect 199811 38147 199839 38175
rect 199625 38085 199653 38113
rect 199687 38085 199715 38113
rect 199749 38085 199777 38113
rect 199811 38085 199839 38113
rect 199625 38023 199653 38051
rect 199687 38023 199715 38051
rect 199749 38023 199777 38051
rect 199811 38023 199839 38051
rect 199625 37961 199653 37989
rect 199687 37961 199715 37989
rect 199749 37961 199777 37989
rect 199811 37961 199839 37989
rect 199625 29147 199653 29175
rect 199687 29147 199715 29175
rect 199749 29147 199777 29175
rect 199811 29147 199839 29175
rect 199625 29085 199653 29113
rect 199687 29085 199715 29113
rect 199749 29085 199777 29113
rect 199811 29085 199839 29113
rect 199625 29023 199653 29051
rect 199687 29023 199715 29051
rect 199749 29023 199777 29051
rect 199811 29023 199839 29051
rect 199625 28961 199653 28989
rect 199687 28961 199715 28989
rect 199749 28961 199777 28989
rect 199811 28961 199839 28989
rect 199625 20147 199653 20175
rect 199687 20147 199715 20175
rect 199749 20147 199777 20175
rect 199811 20147 199839 20175
rect 199625 20085 199653 20113
rect 199687 20085 199715 20113
rect 199749 20085 199777 20113
rect 199811 20085 199839 20113
rect 199625 20023 199653 20051
rect 199687 20023 199715 20051
rect 199749 20023 199777 20051
rect 199811 20023 199839 20051
rect 199625 19961 199653 19989
rect 199687 19961 199715 19989
rect 199749 19961 199777 19989
rect 199811 19961 199839 19989
rect 199625 11147 199653 11175
rect 199687 11147 199715 11175
rect 199749 11147 199777 11175
rect 199811 11147 199839 11175
rect 199625 11085 199653 11113
rect 199687 11085 199715 11113
rect 199749 11085 199777 11113
rect 199811 11085 199839 11113
rect 199625 11023 199653 11051
rect 199687 11023 199715 11051
rect 199749 11023 199777 11051
rect 199811 11023 199839 11051
rect 199625 10961 199653 10989
rect 199687 10961 199715 10989
rect 199749 10961 199777 10989
rect 199811 10961 199839 10989
rect 199625 2147 199653 2175
rect 199687 2147 199715 2175
rect 199749 2147 199777 2175
rect 199811 2147 199839 2175
rect 199625 2085 199653 2113
rect 199687 2085 199715 2113
rect 199749 2085 199777 2113
rect 199811 2085 199839 2113
rect 199625 2023 199653 2051
rect 199687 2023 199715 2051
rect 199749 2023 199777 2051
rect 199811 2023 199839 2051
rect 199625 1961 199653 1989
rect 199687 1961 199715 1989
rect 199749 1961 199777 1989
rect 199811 1961 199839 1989
rect 199625 -108 199653 -80
rect 199687 -108 199715 -80
rect 199749 -108 199777 -80
rect 199811 -108 199839 -80
rect 199625 -170 199653 -142
rect 199687 -170 199715 -142
rect 199749 -170 199777 -142
rect 199811 -170 199839 -142
rect 199625 -232 199653 -204
rect 199687 -232 199715 -204
rect 199749 -232 199777 -204
rect 199811 -232 199839 -204
rect 199625 -294 199653 -266
rect 199687 -294 199715 -266
rect 199749 -294 199777 -266
rect 199811 -294 199839 -266
rect 201485 299058 201513 299086
rect 201547 299058 201575 299086
rect 201609 299058 201637 299086
rect 201671 299058 201699 299086
rect 201485 298996 201513 299024
rect 201547 298996 201575 299024
rect 201609 298996 201637 299024
rect 201671 298996 201699 299024
rect 201485 298934 201513 298962
rect 201547 298934 201575 298962
rect 201609 298934 201637 298962
rect 201671 298934 201699 298962
rect 201485 298872 201513 298900
rect 201547 298872 201575 298900
rect 201609 298872 201637 298900
rect 201671 298872 201699 298900
rect 201485 293147 201513 293175
rect 201547 293147 201575 293175
rect 201609 293147 201637 293175
rect 201671 293147 201699 293175
rect 201485 293085 201513 293113
rect 201547 293085 201575 293113
rect 201609 293085 201637 293113
rect 201671 293085 201699 293113
rect 201485 293023 201513 293051
rect 201547 293023 201575 293051
rect 201609 293023 201637 293051
rect 201671 293023 201699 293051
rect 201485 292961 201513 292989
rect 201547 292961 201575 292989
rect 201609 292961 201637 292989
rect 201671 292961 201699 292989
rect 201485 284147 201513 284175
rect 201547 284147 201575 284175
rect 201609 284147 201637 284175
rect 201671 284147 201699 284175
rect 201485 284085 201513 284113
rect 201547 284085 201575 284113
rect 201609 284085 201637 284113
rect 201671 284085 201699 284113
rect 201485 284023 201513 284051
rect 201547 284023 201575 284051
rect 201609 284023 201637 284051
rect 201671 284023 201699 284051
rect 201485 283961 201513 283989
rect 201547 283961 201575 283989
rect 201609 283961 201637 283989
rect 201671 283961 201699 283989
rect 201485 275147 201513 275175
rect 201547 275147 201575 275175
rect 201609 275147 201637 275175
rect 201671 275147 201699 275175
rect 201485 275085 201513 275113
rect 201547 275085 201575 275113
rect 201609 275085 201637 275113
rect 201671 275085 201699 275113
rect 201485 275023 201513 275051
rect 201547 275023 201575 275051
rect 201609 275023 201637 275051
rect 201671 275023 201699 275051
rect 201485 274961 201513 274989
rect 201547 274961 201575 274989
rect 201609 274961 201637 274989
rect 201671 274961 201699 274989
rect 201485 266147 201513 266175
rect 201547 266147 201575 266175
rect 201609 266147 201637 266175
rect 201671 266147 201699 266175
rect 201485 266085 201513 266113
rect 201547 266085 201575 266113
rect 201609 266085 201637 266113
rect 201671 266085 201699 266113
rect 201485 266023 201513 266051
rect 201547 266023 201575 266051
rect 201609 266023 201637 266051
rect 201671 266023 201699 266051
rect 201485 265961 201513 265989
rect 201547 265961 201575 265989
rect 201609 265961 201637 265989
rect 201671 265961 201699 265989
rect 201485 257147 201513 257175
rect 201547 257147 201575 257175
rect 201609 257147 201637 257175
rect 201671 257147 201699 257175
rect 201485 257085 201513 257113
rect 201547 257085 201575 257113
rect 201609 257085 201637 257113
rect 201671 257085 201699 257113
rect 201485 257023 201513 257051
rect 201547 257023 201575 257051
rect 201609 257023 201637 257051
rect 201671 257023 201699 257051
rect 201485 256961 201513 256989
rect 201547 256961 201575 256989
rect 201609 256961 201637 256989
rect 201671 256961 201699 256989
rect 201485 248147 201513 248175
rect 201547 248147 201575 248175
rect 201609 248147 201637 248175
rect 201671 248147 201699 248175
rect 201485 248085 201513 248113
rect 201547 248085 201575 248113
rect 201609 248085 201637 248113
rect 201671 248085 201699 248113
rect 201485 248023 201513 248051
rect 201547 248023 201575 248051
rect 201609 248023 201637 248051
rect 201671 248023 201699 248051
rect 201485 247961 201513 247989
rect 201547 247961 201575 247989
rect 201609 247961 201637 247989
rect 201671 247961 201699 247989
rect 201485 239147 201513 239175
rect 201547 239147 201575 239175
rect 201609 239147 201637 239175
rect 201671 239147 201699 239175
rect 201485 239085 201513 239113
rect 201547 239085 201575 239113
rect 201609 239085 201637 239113
rect 201671 239085 201699 239113
rect 201485 239023 201513 239051
rect 201547 239023 201575 239051
rect 201609 239023 201637 239051
rect 201671 239023 201699 239051
rect 201485 238961 201513 238989
rect 201547 238961 201575 238989
rect 201609 238961 201637 238989
rect 201671 238961 201699 238989
rect 201485 230147 201513 230175
rect 201547 230147 201575 230175
rect 201609 230147 201637 230175
rect 201671 230147 201699 230175
rect 201485 230085 201513 230113
rect 201547 230085 201575 230113
rect 201609 230085 201637 230113
rect 201671 230085 201699 230113
rect 201485 230023 201513 230051
rect 201547 230023 201575 230051
rect 201609 230023 201637 230051
rect 201671 230023 201699 230051
rect 201485 229961 201513 229989
rect 201547 229961 201575 229989
rect 201609 229961 201637 229989
rect 201671 229961 201699 229989
rect 201485 221147 201513 221175
rect 201547 221147 201575 221175
rect 201609 221147 201637 221175
rect 201671 221147 201699 221175
rect 201485 221085 201513 221113
rect 201547 221085 201575 221113
rect 201609 221085 201637 221113
rect 201671 221085 201699 221113
rect 201485 221023 201513 221051
rect 201547 221023 201575 221051
rect 201609 221023 201637 221051
rect 201671 221023 201699 221051
rect 201485 220961 201513 220989
rect 201547 220961 201575 220989
rect 201609 220961 201637 220989
rect 201671 220961 201699 220989
rect 201485 212147 201513 212175
rect 201547 212147 201575 212175
rect 201609 212147 201637 212175
rect 201671 212147 201699 212175
rect 201485 212085 201513 212113
rect 201547 212085 201575 212113
rect 201609 212085 201637 212113
rect 201671 212085 201699 212113
rect 201485 212023 201513 212051
rect 201547 212023 201575 212051
rect 201609 212023 201637 212051
rect 201671 212023 201699 212051
rect 201485 211961 201513 211989
rect 201547 211961 201575 211989
rect 201609 211961 201637 211989
rect 201671 211961 201699 211989
rect 201485 203147 201513 203175
rect 201547 203147 201575 203175
rect 201609 203147 201637 203175
rect 201671 203147 201699 203175
rect 201485 203085 201513 203113
rect 201547 203085 201575 203113
rect 201609 203085 201637 203113
rect 201671 203085 201699 203113
rect 201485 203023 201513 203051
rect 201547 203023 201575 203051
rect 201609 203023 201637 203051
rect 201671 203023 201699 203051
rect 201485 202961 201513 202989
rect 201547 202961 201575 202989
rect 201609 202961 201637 202989
rect 201671 202961 201699 202989
rect 201485 194147 201513 194175
rect 201547 194147 201575 194175
rect 201609 194147 201637 194175
rect 201671 194147 201699 194175
rect 201485 194085 201513 194113
rect 201547 194085 201575 194113
rect 201609 194085 201637 194113
rect 201671 194085 201699 194113
rect 201485 194023 201513 194051
rect 201547 194023 201575 194051
rect 201609 194023 201637 194051
rect 201671 194023 201699 194051
rect 201485 193961 201513 193989
rect 201547 193961 201575 193989
rect 201609 193961 201637 193989
rect 201671 193961 201699 193989
rect 201485 185147 201513 185175
rect 201547 185147 201575 185175
rect 201609 185147 201637 185175
rect 201671 185147 201699 185175
rect 201485 185085 201513 185113
rect 201547 185085 201575 185113
rect 201609 185085 201637 185113
rect 201671 185085 201699 185113
rect 201485 185023 201513 185051
rect 201547 185023 201575 185051
rect 201609 185023 201637 185051
rect 201671 185023 201699 185051
rect 201485 184961 201513 184989
rect 201547 184961 201575 184989
rect 201609 184961 201637 184989
rect 201671 184961 201699 184989
rect 201485 176147 201513 176175
rect 201547 176147 201575 176175
rect 201609 176147 201637 176175
rect 201671 176147 201699 176175
rect 201485 176085 201513 176113
rect 201547 176085 201575 176113
rect 201609 176085 201637 176113
rect 201671 176085 201699 176113
rect 201485 176023 201513 176051
rect 201547 176023 201575 176051
rect 201609 176023 201637 176051
rect 201671 176023 201699 176051
rect 201485 175961 201513 175989
rect 201547 175961 201575 175989
rect 201609 175961 201637 175989
rect 201671 175961 201699 175989
rect 201485 167147 201513 167175
rect 201547 167147 201575 167175
rect 201609 167147 201637 167175
rect 201671 167147 201699 167175
rect 201485 167085 201513 167113
rect 201547 167085 201575 167113
rect 201609 167085 201637 167113
rect 201671 167085 201699 167113
rect 201485 167023 201513 167051
rect 201547 167023 201575 167051
rect 201609 167023 201637 167051
rect 201671 167023 201699 167051
rect 201485 166961 201513 166989
rect 201547 166961 201575 166989
rect 201609 166961 201637 166989
rect 201671 166961 201699 166989
rect 201485 158147 201513 158175
rect 201547 158147 201575 158175
rect 201609 158147 201637 158175
rect 201671 158147 201699 158175
rect 201485 158085 201513 158113
rect 201547 158085 201575 158113
rect 201609 158085 201637 158113
rect 201671 158085 201699 158113
rect 201485 158023 201513 158051
rect 201547 158023 201575 158051
rect 201609 158023 201637 158051
rect 201671 158023 201699 158051
rect 201485 157961 201513 157989
rect 201547 157961 201575 157989
rect 201609 157961 201637 157989
rect 201671 157961 201699 157989
rect 201485 149147 201513 149175
rect 201547 149147 201575 149175
rect 201609 149147 201637 149175
rect 201671 149147 201699 149175
rect 201485 149085 201513 149113
rect 201547 149085 201575 149113
rect 201609 149085 201637 149113
rect 201671 149085 201699 149113
rect 201485 149023 201513 149051
rect 201547 149023 201575 149051
rect 201609 149023 201637 149051
rect 201671 149023 201699 149051
rect 201485 148961 201513 148989
rect 201547 148961 201575 148989
rect 201609 148961 201637 148989
rect 201671 148961 201699 148989
rect 201485 140147 201513 140175
rect 201547 140147 201575 140175
rect 201609 140147 201637 140175
rect 201671 140147 201699 140175
rect 201485 140085 201513 140113
rect 201547 140085 201575 140113
rect 201609 140085 201637 140113
rect 201671 140085 201699 140113
rect 201485 140023 201513 140051
rect 201547 140023 201575 140051
rect 201609 140023 201637 140051
rect 201671 140023 201699 140051
rect 201485 139961 201513 139989
rect 201547 139961 201575 139989
rect 201609 139961 201637 139989
rect 201671 139961 201699 139989
rect 201485 131147 201513 131175
rect 201547 131147 201575 131175
rect 201609 131147 201637 131175
rect 201671 131147 201699 131175
rect 201485 131085 201513 131113
rect 201547 131085 201575 131113
rect 201609 131085 201637 131113
rect 201671 131085 201699 131113
rect 201485 131023 201513 131051
rect 201547 131023 201575 131051
rect 201609 131023 201637 131051
rect 201671 131023 201699 131051
rect 201485 130961 201513 130989
rect 201547 130961 201575 130989
rect 201609 130961 201637 130989
rect 201671 130961 201699 130989
rect 201485 122147 201513 122175
rect 201547 122147 201575 122175
rect 201609 122147 201637 122175
rect 201671 122147 201699 122175
rect 201485 122085 201513 122113
rect 201547 122085 201575 122113
rect 201609 122085 201637 122113
rect 201671 122085 201699 122113
rect 201485 122023 201513 122051
rect 201547 122023 201575 122051
rect 201609 122023 201637 122051
rect 201671 122023 201699 122051
rect 201485 121961 201513 121989
rect 201547 121961 201575 121989
rect 201609 121961 201637 121989
rect 201671 121961 201699 121989
rect 201485 113147 201513 113175
rect 201547 113147 201575 113175
rect 201609 113147 201637 113175
rect 201671 113147 201699 113175
rect 201485 113085 201513 113113
rect 201547 113085 201575 113113
rect 201609 113085 201637 113113
rect 201671 113085 201699 113113
rect 201485 113023 201513 113051
rect 201547 113023 201575 113051
rect 201609 113023 201637 113051
rect 201671 113023 201699 113051
rect 201485 112961 201513 112989
rect 201547 112961 201575 112989
rect 201609 112961 201637 112989
rect 201671 112961 201699 112989
rect 201485 104147 201513 104175
rect 201547 104147 201575 104175
rect 201609 104147 201637 104175
rect 201671 104147 201699 104175
rect 201485 104085 201513 104113
rect 201547 104085 201575 104113
rect 201609 104085 201637 104113
rect 201671 104085 201699 104113
rect 201485 104023 201513 104051
rect 201547 104023 201575 104051
rect 201609 104023 201637 104051
rect 201671 104023 201699 104051
rect 201485 103961 201513 103989
rect 201547 103961 201575 103989
rect 201609 103961 201637 103989
rect 201671 103961 201699 103989
rect 201485 95147 201513 95175
rect 201547 95147 201575 95175
rect 201609 95147 201637 95175
rect 201671 95147 201699 95175
rect 201485 95085 201513 95113
rect 201547 95085 201575 95113
rect 201609 95085 201637 95113
rect 201671 95085 201699 95113
rect 201485 95023 201513 95051
rect 201547 95023 201575 95051
rect 201609 95023 201637 95051
rect 201671 95023 201699 95051
rect 201485 94961 201513 94989
rect 201547 94961 201575 94989
rect 201609 94961 201637 94989
rect 201671 94961 201699 94989
rect 201485 86147 201513 86175
rect 201547 86147 201575 86175
rect 201609 86147 201637 86175
rect 201671 86147 201699 86175
rect 201485 86085 201513 86113
rect 201547 86085 201575 86113
rect 201609 86085 201637 86113
rect 201671 86085 201699 86113
rect 201485 86023 201513 86051
rect 201547 86023 201575 86051
rect 201609 86023 201637 86051
rect 201671 86023 201699 86051
rect 201485 85961 201513 85989
rect 201547 85961 201575 85989
rect 201609 85961 201637 85989
rect 201671 85961 201699 85989
rect 201485 77147 201513 77175
rect 201547 77147 201575 77175
rect 201609 77147 201637 77175
rect 201671 77147 201699 77175
rect 201485 77085 201513 77113
rect 201547 77085 201575 77113
rect 201609 77085 201637 77113
rect 201671 77085 201699 77113
rect 201485 77023 201513 77051
rect 201547 77023 201575 77051
rect 201609 77023 201637 77051
rect 201671 77023 201699 77051
rect 201485 76961 201513 76989
rect 201547 76961 201575 76989
rect 201609 76961 201637 76989
rect 201671 76961 201699 76989
rect 201485 68147 201513 68175
rect 201547 68147 201575 68175
rect 201609 68147 201637 68175
rect 201671 68147 201699 68175
rect 201485 68085 201513 68113
rect 201547 68085 201575 68113
rect 201609 68085 201637 68113
rect 201671 68085 201699 68113
rect 201485 68023 201513 68051
rect 201547 68023 201575 68051
rect 201609 68023 201637 68051
rect 201671 68023 201699 68051
rect 201485 67961 201513 67989
rect 201547 67961 201575 67989
rect 201609 67961 201637 67989
rect 201671 67961 201699 67989
rect 201485 59147 201513 59175
rect 201547 59147 201575 59175
rect 201609 59147 201637 59175
rect 201671 59147 201699 59175
rect 201485 59085 201513 59113
rect 201547 59085 201575 59113
rect 201609 59085 201637 59113
rect 201671 59085 201699 59113
rect 201485 59023 201513 59051
rect 201547 59023 201575 59051
rect 201609 59023 201637 59051
rect 201671 59023 201699 59051
rect 201485 58961 201513 58989
rect 201547 58961 201575 58989
rect 201609 58961 201637 58989
rect 201671 58961 201699 58989
rect 201485 50147 201513 50175
rect 201547 50147 201575 50175
rect 201609 50147 201637 50175
rect 201671 50147 201699 50175
rect 201485 50085 201513 50113
rect 201547 50085 201575 50113
rect 201609 50085 201637 50113
rect 201671 50085 201699 50113
rect 201485 50023 201513 50051
rect 201547 50023 201575 50051
rect 201609 50023 201637 50051
rect 201671 50023 201699 50051
rect 201485 49961 201513 49989
rect 201547 49961 201575 49989
rect 201609 49961 201637 49989
rect 201671 49961 201699 49989
rect 201485 41147 201513 41175
rect 201547 41147 201575 41175
rect 201609 41147 201637 41175
rect 201671 41147 201699 41175
rect 201485 41085 201513 41113
rect 201547 41085 201575 41113
rect 201609 41085 201637 41113
rect 201671 41085 201699 41113
rect 201485 41023 201513 41051
rect 201547 41023 201575 41051
rect 201609 41023 201637 41051
rect 201671 41023 201699 41051
rect 201485 40961 201513 40989
rect 201547 40961 201575 40989
rect 201609 40961 201637 40989
rect 201671 40961 201699 40989
rect 201485 32147 201513 32175
rect 201547 32147 201575 32175
rect 201609 32147 201637 32175
rect 201671 32147 201699 32175
rect 201485 32085 201513 32113
rect 201547 32085 201575 32113
rect 201609 32085 201637 32113
rect 201671 32085 201699 32113
rect 201485 32023 201513 32051
rect 201547 32023 201575 32051
rect 201609 32023 201637 32051
rect 201671 32023 201699 32051
rect 201485 31961 201513 31989
rect 201547 31961 201575 31989
rect 201609 31961 201637 31989
rect 201671 31961 201699 31989
rect 201485 23147 201513 23175
rect 201547 23147 201575 23175
rect 201609 23147 201637 23175
rect 201671 23147 201699 23175
rect 201485 23085 201513 23113
rect 201547 23085 201575 23113
rect 201609 23085 201637 23113
rect 201671 23085 201699 23113
rect 201485 23023 201513 23051
rect 201547 23023 201575 23051
rect 201609 23023 201637 23051
rect 201671 23023 201699 23051
rect 201485 22961 201513 22989
rect 201547 22961 201575 22989
rect 201609 22961 201637 22989
rect 201671 22961 201699 22989
rect 201485 14147 201513 14175
rect 201547 14147 201575 14175
rect 201609 14147 201637 14175
rect 201671 14147 201699 14175
rect 201485 14085 201513 14113
rect 201547 14085 201575 14113
rect 201609 14085 201637 14113
rect 201671 14085 201699 14113
rect 201485 14023 201513 14051
rect 201547 14023 201575 14051
rect 201609 14023 201637 14051
rect 201671 14023 201699 14051
rect 201485 13961 201513 13989
rect 201547 13961 201575 13989
rect 201609 13961 201637 13989
rect 201671 13961 201699 13989
rect 201485 5147 201513 5175
rect 201547 5147 201575 5175
rect 201609 5147 201637 5175
rect 201671 5147 201699 5175
rect 201485 5085 201513 5113
rect 201547 5085 201575 5113
rect 201609 5085 201637 5113
rect 201671 5085 201699 5113
rect 201485 5023 201513 5051
rect 201547 5023 201575 5051
rect 201609 5023 201637 5051
rect 201671 5023 201699 5051
rect 201485 4961 201513 4989
rect 201547 4961 201575 4989
rect 201609 4961 201637 4989
rect 201671 4961 201699 4989
rect 201485 -588 201513 -560
rect 201547 -588 201575 -560
rect 201609 -588 201637 -560
rect 201671 -588 201699 -560
rect 201485 -650 201513 -622
rect 201547 -650 201575 -622
rect 201609 -650 201637 -622
rect 201671 -650 201699 -622
rect 201485 -712 201513 -684
rect 201547 -712 201575 -684
rect 201609 -712 201637 -684
rect 201671 -712 201699 -684
rect 201485 -774 201513 -746
rect 201547 -774 201575 -746
rect 201609 -774 201637 -746
rect 201671 -774 201699 -746
rect 208625 298578 208653 298606
rect 208687 298578 208715 298606
rect 208749 298578 208777 298606
rect 208811 298578 208839 298606
rect 208625 298516 208653 298544
rect 208687 298516 208715 298544
rect 208749 298516 208777 298544
rect 208811 298516 208839 298544
rect 208625 298454 208653 298482
rect 208687 298454 208715 298482
rect 208749 298454 208777 298482
rect 208811 298454 208839 298482
rect 208625 298392 208653 298420
rect 208687 298392 208715 298420
rect 208749 298392 208777 298420
rect 208811 298392 208839 298420
rect 208625 290147 208653 290175
rect 208687 290147 208715 290175
rect 208749 290147 208777 290175
rect 208811 290147 208839 290175
rect 208625 290085 208653 290113
rect 208687 290085 208715 290113
rect 208749 290085 208777 290113
rect 208811 290085 208839 290113
rect 208625 290023 208653 290051
rect 208687 290023 208715 290051
rect 208749 290023 208777 290051
rect 208811 290023 208839 290051
rect 208625 289961 208653 289989
rect 208687 289961 208715 289989
rect 208749 289961 208777 289989
rect 208811 289961 208839 289989
rect 208625 281147 208653 281175
rect 208687 281147 208715 281175
rect 208749 281147 208777 281175
rect 208811 281147 208839 281175
rect 208625 281085 208653 281113
rect 208687 281085 208715 281113
rect 208749 281085 208777 281113
rect 208811 281085 208839 281113
rect 208625 281023 208653 281051
rect 208687 281023 208715 281051
rect 208749 281023 208777 281051
rect 208811 281023 208839 281051
rect 208625 280961 208653 280989
rect 208687 280961 208715 280989
rect 208749 280961 208777 280989
rect 208811 280961 208839 280989
rect 208625 272147 208653 272175
rect 208687 272147 208715 272175
rect 208749 272147 208777 272175
rect 208811 272147 208839 272175
rect 208625 272085 208653 272113
rect 208687 272085 208715 272113
rect 208749 272085 208777 272113
rect 208811 272085 208839 272113
rect 208625 272023 208653 272051
rect 208687 272023 208715 272051
rect 208749 272023 208777 272051
rect 208811 272023 208839 272051
rect 208625 271961 208653 271989
rect 208687 271961 208715 271989
rect 208749 271961 208777 271989
rect 208811 271961 208839 271989
rect 208625 263147 208653 263175
rect 208687 263147 208715 263175
rect 208749 263147 208777 263175
rect 208811 263147 208839 263175
rect 208625 263085 208653 263113
rect 208687 263085 208715 263113
rect 208749 263085 208777 263113
rect 208811 263085 208839 263113
rect 208625 263023 208653 263051
rect 208687 263023 208715 263051
rect 208749 263023 208777 263051
rect 208811 263023 208839 263051
rect 208625 262961 208653 262989
rect 208687 262961 208715 262989
rect 208749 262961 208777 262989
rect 208811 262961 208839 262989
rect 208625 254147 208653 254175
rect 208687 254147 208715 254175
rect 208749 254147 208777 254175
rect 208811 254147 208839 254175
rect 208625 254085 208653 254113
rect 208687 254085 208715 254113
rect 208749 254085 208777 254113
rect 208811 254085 208839 254113
rect 208625 254023 208653 254051
rect 208687 254023 208715 254051
rect 208749 254023 208777 254051
rect 208811 254023 208839 254051
rect 208625 253961 208653 253989
rect 208687 253961 208715 253989
rect 208749 253961 208777 253989
rect 208811 253961 208839 253989
rect 208625 245147 208653 245175
rect 208687 245147 208715 245175
rect 208749 245147 208777 245175
rect 208811 245147 208839 245175
rect 208625 245085 208653 245113
rect 208687 245085 208715 245113
rect 208749 245085 208777 245113
rect 208811 245085 208839 245113
rect 208625 245023 208653 245051
rect 208687 245023 208715 245051
rect 208749 245023 208777 245051
rect 208811 245023 208839 245051
rect 208625 244961 208653 244989
rect 208687 244961 208715 244989
rect 208749 244961 208777 244989
rect 208811 244961 208839 244989
rect 208625 236147 208653 236175
rect 208687 236147 208715 236175
rect 208749 236147 208777 236175
rect 208811 236147 208839 236175
rect 208625 236085 208653 236113
rect 208687 236085 208715 236113
rect 208749 236085 208777 236113
rect 208811 236085 208839 236113
rect 208625 236023 208653 236051
rect 208687 236023 208715 236051
rect 208749 236023 208777 236051
rect 208811 236023 208839 236051
rect 208625 235961 208653 235989
rect 208687 235961 208715 235989
rect 208749 235961 208777 235989
rect 208811 235961 208839 235989
rect 208625 227147 208653 227175
rect 208687 227147 208715 227175
rect 208749 227147 208777 227175
rect 208811 227147 208839 227175
rect 208625 227085 208653 227113
rect 208687 227085 208715 227113
rect 208749 227085 208777 227113
rect 208811 227085 208839 227113
rect 208625 227023 208653 227051
rect 208687 227023 208715 227051
rect 208749 227023 208777 227051
rect 208811 227023 208839 227051
rect 208625 226961 208653 226989
rect 208687 226961 208715 226989
rect 208749 226961 208777 226989
rect 208811 226961 208839 226989
rect 208625 218147 208653 218175
rect 208687 218147 208715 218175
rect 208749 218147 208777 218175
rect 208811 218147 208839 218175
rect 208625 218085 208653 218113
rect 208687 218085 208715 218113
rect 208749 218085 208777 218113
rect 208811 218085 208839 218113
rect 208625 218023 208653 218051
rect 208687 218023 208715 218051
rect 208749 218023 208777 218051
rect 208811 218023 208839 218051
rect 208625 217961 208653 217989
rect 208687 217961 208715 217989
rect 208749 217961 208777 217989
rect 208811 217961 208839 217989
rect 208625 209147 208653 209175
rect 208687 209147 208715 209175
rect 208749 209147 208777 209175
rect 208811 209147 208839 209175
rect 208625 209085 208653 209113
rect 208687 209085 208715 209113
rect 208749 209085 208777 209113
rect 208811 209085 208839 209113
rect 208625 209023 208653 209051
rect 208687 209023 208715 209051
rect 208749 209023 208777 209051
rect 208811 209023 208839 209051
rect 208625 208961 208653 208989
rect 208687 208961 208715 208989
rect 208749 208961 208777 208989
rect 208811 208961 208839 208989
rect 208625 200147 208653 200175
rect 208687 200147 208715 200175
rect 208749 200147 208777 200175
rect 208811 200147 208839 200175
rect 208625 200085 208653 200113
rect 208687 200085 208715 200113
rect 208749 200085 208777 200113
rect 208811 200085 208839 200113
rect 208625 200023 208653 200051
rect 208687 200023 208715 200051
rect 208749 200023 208777 200051
rect 208811 200023 208839 200051
rect 208625 199961 208653 199989
rect 208687 199961 208715 199989
rect 208749 199961 208777 199989
rect 208811 199961 208839 199989
rect 208625 191147 208653 191175
rect 208687 191147 208715 191175
rect 208749 191147 208777 191175
rect 208811 191147 208839 191175
rect 208625 191085 208653 191113
rect 208687 191085 208715 191113
rect 208749 191085 208777 191113
rect 208811 191085 208839 191113
rect 208625 191023 208653 191051
rect 208687 191023 208715 191051
rect 208749 191023 208777 191051
rect 208811 191023 208839 191051
rect 208625 190961 208653 190989
rect 208687 190961 208715 190989
rect 208749 190961 208777 190989
rect 208811 190961 208839 190989
rect 208625 182147 208653 182175
rect 208687 182147 208715 182175
rect 208749 182147 208777 182175
rect 208811 182147 208839 182175
rect 208625 182085 208653 182113
rect 208687 182085 208715 182113
rect 208749 182085 208777 182113
rect 208811 182085 208839 182113
rect 208625 182023 208653 182051
rect 208687 182023 208715 182051
rect 208749 182023 208777 182051
rect 208811 182023 208839 182051
rect 208625 181961 208653 181989
rect 208687 181961 208715 181989
rect 208749 181961 208777 181989
rect 208811 181961 208839 181989
rect 208625 173147 208653 173175
rect 208687 173147 208715 173175
rect 208749 173147 208777 173175
rect 208811 173147 208839 173175
rect 208625 173085 208653 173113
rect 208687 173085 208715 173113
rect 208749 173085 208777 173113
rect 208811 173085 208839 173113
rect 208625 173023 208653 173051
rect 208687 173023 208715 173051
rect 208749 173023 208777 173051
rect 208811 173023 208839 173051
rect 208625 172961 208653 172989
rect 208687 172961 208715 172989
rect 208749 172961 208777 172989
rect 208811 172961 208839 172989
rect 208625 164147 208653 164175
rect 208687 164147 208715 164175
rect 208749 164147 208777 164175
rect 208811 164147 208839 164175
rect 208625 164085 208653 164113
rect 208687 164085 208715 164113
rect 208749 164085 208777 164113
rect 208811 164085 208839 164113
rect 208625 164023 208653 164051
rect 208687 164023 208715 164051
rect 208749 164023 208777 164051
rect 208811 164023 208839 164051
rect 208625 163961 208653 163989
rect 208687 163961 208715 163989
rect 208749 163961 208777 163989
rect 208811 163961 208839 163989
rect 208625 155147 208653 155175
rect 208687 155147 208715 155175
rect 208749 155147 208777 155175
rect 208811 155147 208839 155175
rect 208625 155085 208653 155113
rect 208687 155085 208715 155113
rect 208749 155085 208777 155113
rect 208811 155085 208839 155113
rect 208625 155023 208653 155051
rect 208687 155023 208715 155051
rect 208749 155023 208777 155051
rect 208811 155023 208839 155051
rect 208625 154961 208653 154989
rect 208687 154961 208715 154989
rect 208749 154961 208777 154989
rect 208811 154961 208839 154989
rect 208625 146147 208653 146175
rect 208687 146147 208715 146175
rect 208749 146147 208777 146175
rect 208811 146147 208839 146175
rect 208625 146085 208653 146113
rect 208687 146085 208715 146113
rect 208749 146085 208777 146113
rect 208811 146085 208839 146113
rect 208625 146023 208653 146051
rect 208687 146023 208715 146051
rect 208749 146023 208777 146051
rect 208811 146023 208839 146051
rect 208625 145961 208653 145989
rect 208687 145961 208715 145989
rect 208749 145961 208777 145989
rect 208811 145961 208839 145989
rect 208625 137147 208653 137175
rect 208687 137147 208715 137175
rect 208749 137147 208777 137175
rect 208811 137147 208839 137175
rect 208625 137085 208653 137113
rect 208687 137085 208715 137113
rect 208749 137085 208777 137113
rect 208811 137085 208839 137113
rect 208625 137023 208653 137051
rect 208687 137023 208715 137051
rect 208749 137023 208777 137051
rect 208811 137023 208839 137051
rect 208625 136961 208653 136989
rect 208687 136961 208715 136989
rect 208749 136961 208777 136989
rect 208811 136961 208839 136989
rect 208625 128147 208653 128175
rect 208687 128147 208715 128175
rect 208749 128147 208777 128175
rect 208811 128147 208839 128175
rect 208625 128085 208653 128113
rect 208687 128085 208715 128113
rect 208749 128085 208777 128113
rect 208811 128085 208839 128113
rect 208625 128023 208653 128051
rect 208687 128023 208715 128051
rect 208749 128023 208777 128051
rect 208811 128023 208839 128051
rect 208625 127961 208653 127989
rect 208687 127961 208715 127989
rect 208749 127961 208777 127989
rect 208811 127961 208839 127989
rect 208625 119147 208653 119175
rect 208687 119147 208715 119175
rect 208749 119147 208777 119175
rect 208811 119147 208839 119175
rect 208625 119085 208653 119113
rect 208687 119085 208715 119113
rect 208749 119085 208777 119113
rect 208811 119085 208839 119113
rect 208625 119023 208653 119051
rect 208687 119023 208715 119051
rect 208749 119023 208777 119051
rect 208811 119023 208839 119051
rect 208625 118961 208653 118989
rect 208687 118961 208715 118989
rect 208749 118961 208777 118989
rect 208811 118961 208839 118989
rect 208625 110147 208653 110175
rect 208687 110147 208715 110175
rect 208749 110147 208777 110175
rect 208811 110147 208839 110175
rect 208625 110085 208653 110113
rect 208687 110085 208715 110113
rect 208749 110085 208777 110113
rect 208811 110085 208839 110113
rect 208625 110023 208653 110051
rect 208687 110023 208715 110051
rect 208749 110023 208777 110051
rect 208811 110023 208839 110051
rect 208625 109961 208653 109989
rect 208687 109961 208715 109989
rect 208749 109961 208777 109989
rect 208811 109961 208839 109989
rect 208625 101147 208653 101175
rect 208687 101147 208715 101175
rect 208749 101147 208777 101175
rect 208811 101147 208839 101175
rect 208625 101085 208653 101113
rect 208687 101085 208715 101113
rect 208749 101085 208777 101113
rect 208811 101085 208839 101113
rect 208625 101023 208653 101051
rect 208687 101023 208715 101051
rect 208749 101023 208777 101051
rect 208811 101023 208839 101051
rect 208625 100961 208653 100989
rect 208687 100961 208715 100989
rect 208749 100961 208777 100989
rect 208811 100961 208839 100989
rect 208625 92147 208653 92175
rect 208687 92147 208715 92175
rect 208749 92147 208777 92175
rect 208811 92147 208839 92175
rect 208625 92085 208653 92113
rect 208687 92085 208715 92113
rect 208749 92085 208777 92113
rect 208811 92085 208839 92113
rect 208625 92023 208653 92051
rect 208687 92023 208715 92051
rect 208749 92023 208777 92051
rect 208811 92023 208839 92051
rect 208625 91961 208653 91989
rect 208687 91961 208715 91989
rect 208749 91961 208777 91989
rect 208811 91961 208839 91989
rect 208625 83147 208653 83175
rect 208687 83147 208715 83175
rect 208749 83147 208777 83175
rect 208811 83147 208839 83175
rect 208625 83085 208653 83113
rect 208687 83085 208715 83113
rect 208749 83085 208777 83113
rect 208811 83085 208839 83113
rect 208625 83023 208653 83051
rect 208687 83023 208715 83051
rect 208749 83023 208777 83051
rect 208811 83023 208839 83051
rect 208625 82961 208653 82989
rect 208687 82961 208715 82989
rect 208749 82961 208777 82989
rect 208811 82961 208839 82989
rect 208625 74147 208653 74175
rect 208687 74147 208715 74175
rect 208749 74147 208777 74175
rect 208811 74147 208839 74175
rect 208625 74085 208653 74113
rect 208687 74085 208715 74113
rect 208749 74085 208777 74113
rect 208811 74085 208839 74113
rect 208625 74023 208653 74051
rect 208687 74023 208715 74051
rect 208749 74023 208777 74051
rect 208811 74023 208839 74051
rect 208625 73961 208653 73989
rect 208687 73961 208715 73989
rect 208749 73961 208777 73989
rect 208811 73961 208839 73989
rect 208625 65147 208653 65175
rect 208687 65147 208715 65175
rect 208749 65147 208777 65175
rect 208811 65147 208839 65175
rect 208625 65085 208653 65113
rect 208687 65085 208715 65113
rect 208749 65085 208777 65113
rect 208811 65085 208839 65113
rect 208625 65023 208653 65051
rect 208687 65023 208715 65051
rect 208749 65023 208777 65051
rect 208811 65023 208839 65051
rect 208625 64961 208653 64989
rect 208687 64961 208715 64989
rect 208749 64961 208777 64989
rect 208811 64961 208839 64989
rect 208625 56147 208653 56175
rect 208687 56147 208715 56175
rect 208749 56147 208777 56175
rect 208811 56147 208839 56175
rect 208625 56085 208653 56113
rect 208687 56085 208715 56113
rect 208749 56085 208777 56113
rect 208811 56085 208839 56113
rect 208625 56023 208653 56051
rect 208687 56023 208715 56051
rect 208749 56023 208777 56051
rect 208811 56023 208839 56051
rect 208625 55961 208653 55989
rect 208687 55961 208715 55989
rect 208749 55961 208777 55989
rect 208811 55961 208839 55989
rect 208625 47147 208653 47175
rect 208687 47147 208715 47175
rect 208749 47147 208777 47175
rect 208811 47147 208839 47175
rect 208625 47085 208653 47113
rect 208687 47085 208715 47113
rect 208749 47085 208777 47113
rect 208811 47085 208839 47113
rect 208625 47023 208653 47051
rect 208687 47023 208715 47051
rect 208749 47023 208777 47051
rect 208811 47023 208839 47051
rect 208625 46961 208653 46989
rect 208687 46961 208715 46989
rect 208749 46961 208777 46989
rect 208811 46961 208839 46989
rect 208625 38147 208653 38175
rect 208687 38147 208715 38175
rect 208749 38147 208777 38175
rect 208811 38147 208839 38175
rect 208625 38085 208653 38113
rect 208687 38085 208715 38113
rect 208749 38085 208777 38113
rect 208811 38085 208839 38113
rect 208625 38023 208653 38051
rect 208687 38023 208715 38051
rect 208749 38023 208777 38051
rect 208811 38023 208839 38051
rect 208625 37961 208653 37989
rect 208687 37961 208715 37989
rect 208749 37961 208777 37989
rect 208811 37961 208839 37989
rect 208625 29147 208653 29175
rect 208687 29147 208715 29175
rect 208749 29147 208777 29175
rect 208811 29147 208839 29175
rect 208625 29085 208653 29113
rect 208687 29085 208715 29113
rect 208749 29085 208777 29113
rect 208811 29085 208839 29113
rect 208625 29023 208653 29051
rect 208687 29023 208715 29051
rect 208749 29023 208777 29051
rect 208811 29023 208839 29051
rect 208625 28961 208653 28989
rect 208687 28961 208715 28989
rect 208749 28961 208777 28989
rect 208811 28961 208839 28989
rect 208625 20147 208653 20175
rect 208687 20147 208715 20175
rect 208749 20147 208777 20175
rect 208811 20147 208839 20175
rect 208625 20085 208653 20113
rect 208687 20085 208715 20113
rect 208749 20085 208777 20113
rect 208811 20085 208839 20113
rect 208625 20023 208653 20051
rect 208687 20023 208715 20051
rect 208749 20023 208777 20051
rect 208811 20023 208839 20051
rect 208625 19961 208653 19989
rect 208687 19961 208715 19989
rect 208749 19961 208777 19989
rect 208811 19961 208839 19989
rect 208625 11147 208653 11175
rect 208687 11147 208715 11175
rect 208749 11147 208777 11175
rect 208811 11147 208839 11175
rect 208625 11085 208653 11113
rect 208687 11085 208715 11113
rect 208749 11085 208777 11113
rect 208811 11085 208839 11113
rect 208625 11023 208653 11051
rect 208687 11023 208715 11051
rect 208749 11023 208777 11051
rect 208811 11023 208839 11051
rect 208625 10961 208653 10989
rect 208687 10961 208715 10989
rect 208749 10961 208777 10989
rect 208811 10961 208839 10989
rect 208625 2147 208653 2175
rect 208687 2147 208715 2175
rect 208749 2147 208777 2175
rect 208811 2147 208839 2175
rect 208625 2085 208653 2113
rect 208687 2085 208715 2113
rect 208749 2085 208777 2113
rect 208811 2085 208839 2113
rect 208625 2023 208653 2051
rect 208687 2023 208715 2051
rect 208749 2023 208777 2051
rect 208811 2023 208839 2051
rect 208625 1961 208653 1989
rect 208687 1961 208715 1989
rect 208749 1961 208777 1989
rect 208811 1961 208839 1989
rect 208625 -108 208653 -80
rect 208687 -108 208715 -80
rect 208749 -108 208777 -80
rect 208811 -108 208839 -80
rect 208625 -170 208653 -142
rect 208687 -170 208715 -142
rect 208749 -170 208777 -142
rect 208811 -170 208839 -142
rect 208625 -232 208653 -204
rect 208687 -232 208715 -204
rect 208749 -232 208777 -204
rect 208811 -232 208839 -204
rect 208625 -294 208653 -266
rect 208687 -294 208715 -266
rect 208749 -294 208777 -266
rect 208811 -294 208839 -266
rect 210485 299058 210513 299086
rect 210547 299058 210575 299086
rect 210609 299058 210637 299086
rect 210671 299058 210699 299086
rect 210485 298996 210513 299024
rect 210547 298996 210575 299024
rect 210609 298996 210637 299024
rect 210671 298996 210699 299024
rect 210485 298934 210513 298962
rect 210547 298934 210575 298962
rect 210609 298934 210637 298962
rect 210671 298934 210699 298962
rect 210485 298872 210513 298900
rect 210547 298872 210575 298900
rect 210609 298872 210637 298900
rect 210671 298872 210699 298900
rect 210485 293147 210513 293175
rect 210547 293147 210575 293175
rect 210609 293147 210637 293175
rect 210671 293147 210699 293175
rect 210485 293085 210513 293113
rect 210547 293085 210575 293113
rect 210609 293085 210637 293113
rect 210671 293085 210699 293113
rect 210485 293023 210513 293051
rect 210547 293023 210575 293051
rect 210609 293023 210637 293051
rect 210671 293023 210699 293051
rect 210485 292961 210513 292989
rect 210547 292961 210575 292989
rect 210609 292961 210637 292989
rect 210671 292961 210699 292989
rect 210485 284147 210513 284175
rect 210547 284147 210575 284175
rect 210609 284147 210637 284175
rect 210671 284147 210699 284175
rect 210485 284085 210513 284113
rect 210547 284085 210575 284113
rect 210609 284085 210637 284113
rect 210671 284085 210699 284113
rect 210485 284023 210513 284051
rect 210547 284023 210575 284051
rect 210609 284023 210637 284051
rect 210671 284023 210699 284051
rect 210485 283961 210513 283989
rect 210547 283961 210575 283989
rect 210609 283961 210637 283989
rect 210671 283961 210699 283989
rect 210485 275147 210513 275175
rect 210547 275147 210575 275175
rect 210609 275147 210637 275175
rect 210671 275147 210699 275175
rect 210485 275085 210513 275113
rect 210547 275085 210575 275113
rect 210609 275085 210637 275113
rect 210671 275085 210699 275113
rect 210485 275023 210513 275051
rect 210547 275023 210575 275051
rect 210609 275023 210637 275051
rect 210671 275023 210699 275051
rect 210485 274961 210513 274989
rect 210547 274961 210575 274989
rect 210609 274961 210637 274989
rect 210671 274961 210699 274989
rect 210485 266147 210513 266175
rect 210547 266147 210575 266175
rect 210609 266147 210637 266175
rect 210671 266147 210699 266175
rect 210485 266085 210513 266113
rect 210547 266085 210575 266113
rect 210609 266085 210637 266113
rect 210671 266085 210699 266113
rect 210485 266023 210513 266051
rect 210547 266023 210575 266051
rect 210609 266023 210637 266051
rect 210671 266023 210699 266051
rect 210485 265961 210513 265989
rect 210547 265961 210575 265989
rect 210609 265961 210637 265989
rect 210671 265961 210699 265989
rect 210485 257147 210513 257175
rect 210547 257147 210575 257175
rect 210609 257147 210637 257175
rect 210671 257147 210699 257175
rect 210485 257085 210513 257113
rect 210547 257085 210575 257113
rect 210609 257085 210637 257113
rect 210671 257085 210699 257113
rect 210485 257023 210513 257051
rect 210547 257023 210575 257051
rect 210609 257023 210637 257051
rect 210671 257023 210699 257051
rect 210485 256961 210513 256989
rect 210547 256961 210575 256989
rect 210609 256961 210637 256989
rect 210671 256961 210699 256989
rect 210485 248147 210513 248175
rect 210547 248147 210575 248175
rect 210609 248147 210637 248175
rect 210671 248147 210699 248175
rect 210485 248085 210513 248113
rect 210547 248085 210575 248113
rect 210609 248085 210637 248113
rect 210671 248085 210699 248113
rect 210485 248023 210513 248051
rect 210547 248023 210575 248051
rect 210609 248023 210637 248051
rect 210671 248023 210699 248051
rect 210485 247961 210513 247989
rect 210547 247961 210575 247989
rect 210609 247961 210637 247989
rect 210671 247961 210699 247989
rect 210485 239147 210513 239175
rect 210547 239147 210575 239175
rect 210609 239147 210637 239175
rect 210671 239147 210699 239175
rect 210485 239085 210513 239113
rect 210547 239085 210575 239113
rect 210609 239085 210637 239113
rect 210671 239085 210699 239113
rect 210485 239023 210513 239051
rect 210547 239023 210575 239051
rect 210609 239023 210637 239051
rect 210671 239023 210699 239051
rect 210485 238961 210513 238989
rect 210547 238961 210575 238989
rect 210609 238961 210637 238989
rect 210671 238961 210699 238989
rect 210485 230147 210513 230175
rect 210547 230147 210575 230175
rect 210609 230147 210637 230175
rect 210671 230147 210699 230175
rect 210485 230085 210513 230113
rect 210547 230085 210575 230113
rect 210609 230085 210637 230113
rect 210671 230085 210699 230113
rect 210485 230023 210513 230051
rect 210547 230023 210575 230051
rect 210609 230023 210637 230051
rect 210671 230023 210699 230051
rect 210485 229961 210513 229989
rect 210547 229961 210575 229989
rect 210609 229961 210637 229989
rect 210671 229961 210699 229989
rect 210485 221147 210513 221175
rect 210547 221147 210575 221175
rect 210609 221147 210637 221175
rect 210671 221147 210699 221175
rect 210485 221085 210513 221113
rect 210547 221085 210575 221113
rect 210609 221085 210637 221113
rect 210671 221085 210699 221113
rect 210485 221023 210513 221051
rect 210547 221023 210575 221051
rect 210609 221023 210637 221051
rect 210671 221023 210699 221051
rect 210485 220961 210513 220989
rect 210547 220961 210575 220989
rect 210609 220961 210637 220989
rect 210671 220961 210699 220989
rect 210485 212147 210513 212175
rect 210547 212147 210575 212175
rect 210609 212147 210637 212175
rect 210671 212147 210699 212175
rect 210485 212085 210513 212113
rect 210547 212085 210575 212113
rect 210609 212085 210637 212113
rect 210671 212085 210699 212113
rect 210485 212023 210513 212051
rect 210547 212023 210575 212051
rect 210609 212023 210637 212051
rect 210671 212023 210699 212051
rect 210485 211961 210513 211989
rect 210547 211961 210575 211989
rect 210609 211961 210637 211989
rect 210671 211961 210699 211989
rect 210485 203147 210513 203175
rect 210547 203147 210575 203175
rect 210609 203147 210637 203175
rect 210671 203147 210699 203175
rect 210485 203085 210513 203113
rect 210547 203085 210575 203113
rect 210609 203085 210637 203113
rect 210671 203085 210699 203113
rect 210485 203023 210513 203051
rect 210547 203023 210575 203051
rect 210609 203023 210637 203051
rect 210671 203023 210699 203051
rect 210485 202961 210513 202989
rect 210547 202961 210575 202989
rect 210609 202961 210637 202989
rect 210671 202961 210699 202989
rect 210485 194147 210513 194175
rect 210547 194147 210575 194175
rect 210609 194147 210637 194175
rect 210671 194147 210699 194175
rect 210485 194085 210513 194113
rect 210547 194085 210575 194113
rect 210609 194085 210637 194113
rect 210671 194085 210699 194113
rect 210485 194023 210513 194051
rect 210547 194023 210575 194051
rect 210609 194023 210637 194051
rect 210671 194023 210699 194051
rect 210485 193961 210513 193989
rect 210547 193961 210575 193989
rect 210609 193961 210637 193989
rect 210671 193961 210699 193989
rect 210485 185147 210513 185175
rect 210547 185147 210575 185175
rect 210609 185147 210637 185175
rect 210671 185147 210699 185175
rect 210485 185085 210513 185113
rect 210547 185085 210575 185113
rect 210609 185085 210637 185113
rect 210671 185085 210699 185113
rect 210485 185023 210513 185051
rect 210547 185023 210575 185051
rect 210609 185023 210637 185051
rect 210671 185023 210699 185051
rect 210485 184961 210513 184989
rect 210547 184961 210575 184989
rect 210609 184961 210637 184989
rect 210671 184961 210699 184989
rect 210485 176147 210513 176175
rect 210547 176147 210575 176175
rect 210609 176147 210637 176175
rect 210671 176147 210699 176175
rect 210485 176085 210513 176113
rect 210547 176085 210575 176113
rect 210609 176085 210637 176113
rect 210671 176085 210699 176113
rect 210485 176023 210513 176051
rect 210547 176023 210575 176051
rect 210609 176023 210637 176051
rect 210671 176023 210699 176051
rect 210485 175961 210513 175989
rect 210547 175961 210575 175989
rect 210609 175961 210637 175989
rect 210671 175961 210699 175989
rect 210485 167147 210513 167175
rect 210547 167147 210575 167175
rect 210609 167147 210637 167175
rect 210671 167147 210699 167175
rect 210485 167085 210513 167113
rect 210547 167085 210575 167113
rect 210609 167085 210637 167113
rect 210671 167085 210699 167113
rect 210485 167023 210513 167051
rect 210547 167023 210575 167051
rect 210609 167023 210637 167051
rect 210671 167023 210699 167051
rect 210485 166961 210513 166989
rect 210547 166961 210575 166989
rect 210609 166961 210637 166989
rect 210671 166961 210699 166989
rect 210485 158147 210513 158175
rect 210547 158147 210575 158175
rect 210609 158147 210637 158175
rect 210671 158147 210699 158175
rect 210485 158085 210513 158113
rect 210547 158085 210575 158113
rect 210609 158085 210637 158113
rect 210671 158085 210699 158113
rect 210485 158023 210513 158051
rect 210547 158023 210575 158051
rect 210609 158023 210637 158051
rect 210671 158023 210699 158051
rect 210485 157961 210513 157989
rect 210547 157961 210575 157989
rect 210609 157961 210637 157989
rect 210671 157961 210699 157989
rect 210485 149147 210513 149175
rect 210547 149147 210575 149175
rect 210609 149147 210637 149175
rect 210671 149147 210699 149175
rect 210485 149085 210513 149113
rect 210547 149085 210575 149113
rect 210609 149085 210637 149113
rect 210671 149085 210699 149113
rect 210485 149023 210513 149051
rect 210547 149023 210575 149051
rect 210609 149023 210637 149051
rect 210671 149023 210699 149051
rect 210485 148961 210513 148989
rect 210547 148961 210575 148989
rect 210609 148961 210637 148989
rect 210671 148961 210699 148989
rect 210485 140147 210513 140175
rect 210547 140147 210575 140175
rect 210609 140147 210637 140175
rect 210671 140147 210699 140175
rect 210485 140085 210513 140113
rect 210547 140085 210575 140113
rect 210609 140085 210637 140113
rect 210671 140085 210699 140113
rect 210485 140023 210513 140051
rect 210547 140023 210575 140051
rect 210609 140023 210637 140051
rect 210671 140023 210699 140051
rect 210485 139961 210513 139989
rect 210547 139961 210575 139989
rect 210609 139961 210637 139989
rect 210671 139961 210699 139989
rect 210485 131147 210513 131175
rect 210547 131147 210575 131175
rect 210609 131147 210637 131175
rect 210671 131147 210699 131175
rect 210485 131085 210513 131113
rect 210547 131085 210575 131113
rect 210609 131085 210637 131113
rect 210671 131085 210699 131113
rect 210485 131023 210513 131051
rect 210547 131023 210575 131051
rect 210609 131023 210637 131051
rect 210671 131023 210699 131051
rect 210485 130961 210513 130989
rect 210547 130961 210575 130989
rect 210609 130961 210637 130989
rect 210671 130961 210699 130989
rect 210485 122147 210513 122175
rect 210547 122147 210575 122175
rect 210609 122147 210637 122175
rect 210671 122147 210699 122175
rect 210485 122085 210513 122113
rect 210547 122085 210575 122113
rect 210609 122085 210637 122113
rect 210671 122085 210699 122113
rect 210485 122023 210513 122051
rect 210547 122023 210575 122051
rect 210609 122023 210637 122051
rect 210671 122023 210699 122051
rect 210485 121961 210513 121989
rect 210547 121961 210575 121989
rect 210609 121961 210637 121989
rect 210671 121961 210699 121989
rect 210485 113147 210513 113175
rect 210547 113147 210575 113175
rect 210609 113147 210637 113175
rect 210671 113147 210699 113175
rect 210485 113085 210513 113113
rect 210547 113085 210575 113113
rect 210609 113085 210637 113113
rect 210671 113085 210699 113113
rect 210485 113023 210513 113051
rect 210547 113023 210575 113051
rect 210609 113023 210637 113051
rect 210671 113023 210699 113051
rect 210485 112961 210513 112989
rect 210547 112961 210575 112989
rect 210609 112961 210637 112989
rect 210671 112961 210699 112989
rect 210485 104147 210513 104175
rect 210547 104147 210575 104175
rect 210609 104147 210637 104175
rect 210671 104147 210699 104175
rect 210485 104085 210513 104113
rect 210547 104085 210575 104113
rect 210609 104085 210637 104113
rect 210671 104085 210699 104113
rect 210485 104023 210513 104051
rect 210547 104023 210575 104051
rect 210609 104023 210637 104051
rect 210671 104023 210699 104051
rect 210485 103961 210513 103989
rect 210547 103961 210575 103989
rect 210609 103961 210637 103989
rect 210671 103961 210699 103989
rect 210485 95147 210513 95175
rect 210547 95147 210575 95175
rect 210609 95147 210637 95175
rect 210671 95147 210699 95175
rect 210485 95085 210513 95113
rect 210547 95085 210575 95113
rect 210609 95085 210637 95113
rect 210671 95085 210699 95113
rect 210485 95023 210513 95051
rect 210547 95023 210575 95051
rect 210609 95023 210637 95051
rect 210671 95023 210699 95051
rect 210485 94961 210513 94989
rect 210547 94961 210575 94989
rect 210609 94961 210637 94989
rect 210671 94961 210699 94989
rect 210485 86147 210513 86175
rect 210547 86147 210575 86175
rect 210609 86147 210637 86175
rect 210671 86147 210699 86175
rect 210485 86085 210513 86113
rect 210547 86085 210575 86113
rect 210609 86085 210637 86113
rect 210671 86085 210699 86113
rect 210485 86023 210513 86051
rect 210547 86023 210575 86051
rect 210609 86023 210637 86051
rect 210671 86023 210699 86051
rect 210485 85961 210513 85989
rect 210547 85961 210575 85989
rect 210609 85961 210637 85989
rect 210671 85961 210699 85989
rect 210485 77147 210513 77175
rect 210547 77147 210575 77175
rect 210609 77147 210637 77175
rect 210671 77147 210699 77175
rect 210485 77085 210513 77113
rect 210547 77085 210575 77113
rect 210609 77085 210637 77113
rect 210671 77085 210699 77113
rect 210485 77023 210513 77051
rect 210547 77023 210575 77051
rect 210609 77023 210637 77051
rect 210671 77023 210699 77051
rect 210485 76961 210513 76989
rect 210547 76961 210575 76989
rect 210609 76961 210637 76989
rect 210671 76961 210699 76989
rect 210485 68147 210513 68175
rect 210547 68147 210575 68175
rect 210609 68147 210637 68175
rect 210671 68147 210699 68175
rect 210485 68085 210513 68113
rect 210547 68085 210575 68113
rect 210609 68085 210637 68113
rect 210671 68085 210699 68113
rect 210485 68023 210513 68051
rect 210547 68023 210575 68051
rect 210609 68023 210637 68051
rect 210671 68023 210699 68051
rect 210485 67961 210513 67989
rect 210547 67961 210575 67989
rect 210609 67961 210637 67989
rect 210671 67961 210699 67989
rect 210485 59147 210513 59175
rect 210547 59147 210575 59175
rect 210609 59147 210637 59175
rect 210671 59147 210699 59175
rect 210485 59085 210513 59113
rect 210547 59085 210575 59113
rect 210609 59085 210637 59113
rect 210671 59085 210699 59113
rect 210485 59023 210513 59051
rect 210547 59023 210575 59051
rect 210609 59023 210637 59051
rect 210671 59023 210699 59051
rect 210485 58961 210513 58989
rect 210547 58961 210575 58989
rect 210609 58961 210637 58989
rect 210671 58961 210699 58989
rect 210485 50147 210513 50175
rect 210547 50147 210575 50175
rect 210609 50147 210637 50175
rect 210671 50147 210699 50175
rect 210485 50085 210513 50113
rect 210547 50085 210575 50113
rect 210609 50085 210637 50113
rect 210671 50085 210699 50113
rect 210485 50023 210513 50051
rect 210547 50023 210575 50051
rect 210609 50023 210637 50051
rect 210671 50023 210699 50051
rect 210485 49961 210513 49989
rect 210547 49961 210575 49989
rect 210609 49961 210637 49989
rect 210671 49961 210699 49989
rect 210485 41147 210513 41175
rect 210547 41147 210575 41175
rect 210609 41147 210637 41175
rect 210671 41147 210699 41175
rect 210485 41085 210513 41113
rect 210547 41085 210575 41113
rect 210609 41085 210637 41113
rect 210671 41085 210699 41113
rect 210485 41023 210513 41051
rect 210547 41023 210575 41051
rect 210609 41023 210637 41051
rect 210671 41023 210699 41051
rect 210485 40961 210513 40989
rect 210547 40961 210575 40989
rect 210609 40961 210637 40989
rect 210671 40961 210699 40989
rect 210485 32147 210513 32175
rect 210547 32147 210575 32175
rect 210609 32147 210637 32175
rect 210671 32147 210699 32175
rect 210485 32085 210513 32113
rect 210547 32085 210575 32113
rect 210609 32085 210637 32113
rect 210671 32085 210699 32113
rect 210485 32023 210513 32051
rect 210547 32023 210575 32051
rect 210609 32023 210637 32051
rect 210671 32023 210699 32051
rect 210485 31961 210513 31989
rect 210547 31961 210575 31989
rect 210609 31961 210637 31989
rect 210671 31961 210699 31989
rect 210485 23147 210513 23175
rect 210547 23147 210575 23175
rect 210609 23147 210637 23175
rect 210671 23147 210699 23175
rect 210485 23085 210513 23113
rect 210547 23085 210575 23113
rect 210609 23085 210637 23113
rect 210671 23085 210699 23113
rect 210485 23023 210513 23051
rect 210547 23023 210575 23051
rect 210609 23023 210637 23051
rect 210671 23023 210699 23051
rect 210485 22961 210513 22989
rect 210547 22961 210575 22989
rect 210609 22961 210637 22989
rect 210671 22961 210699 22989
rect 210485 14147 210513 14175
rect 210547 14147 210575 14175
rect 210609 14147 210637 14175
rect 210671 14147 210699 14175
rect 210485 14085 210513 14113
rect 210547 14085 210575 14113
rect 210609 14085 210637 14113
rect 210671 14085 210699 14113
rect 210485 14023 210513 14051
rect 210547 14023 210575 14051
rect 210609 14023 210637 14051
rect 210671 14023 210699 14051
rect 210485 13961 210513 13989
rect 210547 13961 210575 13989
rect 210609 13961 210637 13989
rect 210671 13961 210699 13989
rect 210485 5147 210513 5175
rect 210547 5147 210575 5175
rect 210609 5147 210637 5175
rect 210671 5147 210699 5175
rect 210485 5085 210513 5113
rect 210547 5085 210575 5113
rect 210609 5085 210637 5113
rect 210671 5085 210699 5113
rect 210485 5023 210513 5051
rect 210547 5023 210575 5051
rect 210609 5023 210637 5051
rect 210671 5023 210699 5051
rect 210485 4961 210513 4989
rect 210547 4961 210575 4989
rect 210609 4961 210637 4989
rect 210671 4961 210699 4989
rect 210485 -588 210513 -560
rect 210547 -588 210575 -560
rect 210609 -588 210637 -560
rect 210671 -588 210699 -560
rect 210485 -650 210513 -622
rect 210547 -650 210575 -622
rect 210609 -650 210637 -622
rect 210671 -650 210699 -622
rect 210485 -712 210513 -684
rect 210547 -712 210575 -684
rect 210609 -712 210637 -684
rect 210671 -712 210699 -684
rect 210485 -774 210513 -746
rect 210547 -774 210575 -746
rect 210609 -774 210637 -746
rect 210671 -774 210699 -746
rect 217625 298578 217653 298606
rect 217687 298578 217715 298606
rect 217749 298578 217777 298606
rect 217811 298578 217839 298606
rect 217625 298516 217653 298544
rect 217687 298516 217715 298544
rect 217749 298516 217777 298544
rect 217811 298516 217839 298544
rect 217625 298454 217653 298482
rect 217687 298454 217715 298482
rect 217749 298454 217777 298482
rect 217811 298454 217839 298482
rect 217625 298392 217653 298420
rect 217687 298392 217715 298420
rect 217749 298392 217777 298420
rect 217811 298392 217839 298420
rect 217625 290147 217653 290175
rect 217687 290147 217715 290175
rect 217749 290147 217777 290175
rect 217811 290147 217839 290175
rect 217625 290085 217653 290113
rect 217687 290085 217715 290113
rect 217749 290085 217777 290113
rect 217811 290085 217839 290113
rect 217625 290023 217653 290051
rect 217687 290023 217715 290051
rect 217749 290023 217777 290051
rect 217811 290023 217839 290051
rect 217625 289961 217653 289989
rect 217687 289961 217715 289989
rect 217749 289961 217777 289989
rect 217811 289961 217839 289989
rect 217625 281147 217653 281175
rect 217687 281147 217715 281175
rect 217749 281147 217777 281175
rect 217811 281147 217839 281175
rect 217625 281085 217653 281113
rect 217687 281085 217715 281113
rect 217749 281085 217777 281113
rect 217811 281085 217839 281113
rect 217625 281023 217653 281051
rect 217687 281023 217715 281051
rect 217749 281023 217777 281051
rect 217811 281023 217839 281051
rect 217625 280961 217653 280989
rect 217687 280961 217715 280989
rect 217749 280961 217777 280989
rect 217811 280961 217839 280989
rect 217625 272147 217653 272175
rect 217687 272147 217715 272175
rect 217749 272147 217777 272175
rect 217811 272147 217839 272175
rect 217625 272085 217653 272113
rect 217687 272085 217715 272113
rect 217749 272085 217777 272113
rect 217811 272085 217839 272113
rect 217625 272023 217653 272051
rect 217687 272023 217715 272051
rect 217749 272023 217777 272051
rect 217811 272023 217839 272051
rect 217625 271961 217653 271989
rect 217687 271961 217715 271989
rect 217749 271961 217777 271989
rect 217811 271961 217839 271989
rect 217625 263147 217653 263175
rect 217687 263147 217715 263175
rect 217749 263147 217777 263175
rect 217811 263147 217839 263175
rect 217625 263085 217653 263113
rect 217687 263085 217715 263113
rect 217749 263085 217777 263113
rect 217811 263085 217839 263113
rect 217625 263023 217653 263051
rect 217687 263023 217715 263051
rect 217749 263023 217777 263051
rect 217811 263023 217839 263051
rect 217625 262961 217653 262989
rect 217687 262961 217715 262989
rect 217749 262961 217777 262989
rect 217811 262961 217839 262989
rect 217625 254147 217653 254175
rect 217687 254147 217715 254175
rect 217749 254147 217777 254175
rect 217811 254147 217839 254175
rect 217625 254085 217653 254113
rect 217687 254085 217715 254113
rect 217749 254085 217777 254113
rect 217811 254085 217839 254113
rect 217625 254023 217653 254051
rect 217687 254023 217715 254051
rect 217749 254023 217777 254051
rect 217811 254023 217839 254051
rect 217625 253961 217653 253989
rect 217687 253961 217715 253989
rect 217749 253961 217777 253989
rect 217811 253961 217839 253989
rect 217625 245147 217653 245175
rect 217687 245147 217715 245175
rect 217749 245147 217777 245175
rect 217811 245147 217839 245175
rect 217625 245085 217653 245113
rect 217687 245085 217715 245113
rect 217749 245085 217777 245113
rect 217811 245085 217839 245113
rect 217625 245023 217653 245051
rect 217687 245023 217715 245051
rect 217749 245023 217777 245051
rect 217811 245023 217839 245051
rect 217625 244961 217653 244989
rect 217687 244961 217715 244989
rect 217749 244961 217777 244989
rect 217811 244961 217839 244989
rect 217625 236147 217653 236175
rect 217687 236147 217715 236175
rect 217749 236147 217777 236175
rect 217811 236147 217839 236175
rect 217625 236085 217653 236113
rect 217687 236085 217715 236113
rect 217749 236085 217777 236113
rect 217811 236085 217839 236113
rect 217625 236023 217653 236051
rect 217687 236023 217715 236051
rect 217749 236023 217777 236051
rect 217811 236023 217839 236051
rect 217625 235961 217653 235989
rect 217687 235961 217715 235989
rect 217749 235961 217777 235989
rect 217811 235961 217839 235989
rect 217625 227147 217653 227175
rect 217687 227147 217715 227175
rect 217749 227147 217777 227175
rect 217811 227147 217839 227175
rect 217625 227085 217653 227113
rect 217687 227085 217715 227113
rect 217749 227085 217777 227113
rect 217811 227085 217839 227113
rect 217625 227023 217653 227051
rect 217687 227023 217715 227051
rect 217749 227023 217777 227051
rect 217811 227023 217839 227051
rect 217625 226961 217653 226989
rect 217687 226961 217715 226989
rect 217749 226961 217777 226989
rect 217811 226961 217839 226989
rect 217625 218147 217653 218175
rect 217687 218147 217715 218175
rect 217749 218147 217777 218175
rect 217811 218147 217839 218175
rect 217625 218085 217653 218113
rect 217687 218085 217715 218113
rect 217749 218085 217777 218113
rect 217811 218085 217839 218113
rect 217625 218023 217653 218051
rect 217687 218023 217715 218051
rect 217749 218023 217777 218051
rect 217811 218023 217839 218051
rect 217625 217961 217653 217989
rect 217687 217961 217715 217989
rect 217749 217961 217777 217989
rect 217811 217961 217839 217989
rect 217625 209147 217653 209175
rect 217687 209147 217715 209175
rect 217749 209147 217777 209175
rect 217811 209147 217839 209175
rect 217625 209085 217653 209113
rect 217687 209085 217715 209113
rect 217749 209085 217777 209113
rect 217811 209085 217839 209113
rect 217625 209023 217653 209051
rect 217687 209023 217715 209051
rect 217749 209023 217777 209051
rect 217811 209023 217839 209051
rect 217625 208961 217653 208989
rect 217687 208961 217715 208989
rect 217749 208961 217777 208989
rect 217811 208961 217839 208989
rect 217625 200147 217653 200175
rect 217687 200147 217715 200175
rect 217749 200147 217777 200175
rect 217811 200147 217839 200175
rect 217625 200085 217653 200113
rect 217687 200085 217715 200113
rect 217749 200085 217777 200113
rect 217811 200085 217839 200113
rect 217625 200023 217653 200051
rect 217687 200023 217715 200051
rect 217749 200023 217777 200051
rect 217811 200023 217839 200051
rect 217625 199961 217653 199989
rect 217687 199961 217715 199989
rect 217749 199961 217777 199989
rect 217811 199961 217839 199989
rect 217625 191147 217653 191175
rect 217687 191147 217715 191175
rect 217749 191147 217777 191175
rect 217811 191147 217839 191175
rect 217625 191085 217653 191113
rect 217687 191085 217715 191113
rect 217749 191085 217777 191113
rect 217811 191085 217839 191113
rect 217625 191023 217653 191051
rect 217687 191023 217715 191051
rect 217749 191023 217777 191051
rect 217811 191023 217839 191051
rect 217625 190961 217653 190989
rect 217687 190961 217715 190989
rect 217749 190961 217777 190989
rect 217811 190961 217839 190989
rect 217625 182147 217653 182175
rect 217687 182147 217715 182175
rect 217749 182147 217777 182175
rect 217811 182147 217839 182175
rect 217625 182085 217653 182113
rect 217687 182085 217715 182113
rect 217749 182085 217777 182113
rect 217811 182085 217839 182113
rect 217625 182023 217653 182051
rect 217687 182023 217715 182051
rect 217749 182023 217777 182051
rect 217811 182023 217839 182051
rect 217625 181961 217653 181989
rect 217687 181961 217715 181989
rect 217749 181961 217777 181989
rect 217811 181961 217839 181989
rect 217625 173147 217653 173175
rect 217687 173147 217715 173175
rect 217749 173147 217777 173175
rect 217811 173147 217839 173175
rect 217625 173085 217653 173113
rect 217687 173085 217715 173113
rect 217749 173085 217777 173113
rect 217811 173085 217839 173113
rect 217625 173023 217653 173051
rect 217687 173023 217715 173051
rect 217749 173023 217777 173051
rect 217811 173023 217839 173051
rect 217625 172961 217653 172989
rect 217687 172961 217715 172989
rect 217749 172961 217777 172989
rect 217811 172961 217839 172989
rect 217625 164147 217653 164175
rect 217687 164147 217715 164175
rect 217749 164147 217777 164175
rect 217811 164147 217839 164175
rect 217625 164085 217653 164113
rect 217687 164085 217715 164113
rect 217749 164085 217777 164113
rect 217811 164085 217839 164113
rect 217625 164023 217653 164051
rect 217687 164023 217715 164051
rect 217749 164023 217777 164051
rect 217811 164023 217839 164051
rect 217625 163961 217653 163989
rect 217687 163961 217715 163989
rect 217749 163961 217777 163989
rect 217811 163961 217839 163989
rect 217625 155147 217653 155175
rect 217687 155147 217715 155175
rect 217749 155147 217777 155175
rect 217811 155147 217839 155175
rect 217625 155085 217653 155113
rect 217687 155085 217715 155113
rect 217749 155085 217777 155113
rect 217811 155085 217839 155113
rect 217625 155023 217653 155051
rect 217687 155023 217715 155051
rect 217749 155023 217777 155051
rect 217811 155023 217839 155051
rect 217625 154961 217653 154989
rect 217687 154961 217715 154989
rect 217749 154961 217777 154989
rect 217811 154961 217839 154989
rect 217625 146147 217653 146175
rect 217687 146147 217715 146175
rect 217749 146147 217777 146175
rect 217811 146147 217839 146175
rect 217625 146085 217653 146113
rect 217687 146085 217715 146113
rect 217749 146085 217777 146113
rect 217811 146085 217839 146113
rect 217625 146023 217653 146051
rect 217687 146023 217715 146051
rect 217749 146023 217777 146051
rect 217811 146023 217839 146051
rect 217625 145961 217653 145989
rect 217687 145961 217715 145989
rect 217749 145961 217777 145989
rect 217811 145961 217839 145989
rect 217625 137147 217653 137175
rect 217687 137147 217715 137175
rect 217749 137147 217777 137175
rect 217811 137147 217839 137175
rect 217625 137085 217653 137113
rect 217687 137085 217715 137113
rect 217749 137085 217777 137113
rect 217811 137085 217839 137113
rect 217625 137023 217653 137051
rect 217687 137023 217715 137051
rect 217749 137023 217777 137051
rect 217811 137023 217839 137051
rect 217625 136961 217653 136989
rect 217687 136961 217715 136989
rect 217749 136961 217777 136989
rect 217811 136961 217839 136989
rect 217625 128147 217653 128175
rect 217687 128147 217715 128175
rect 217749 128147 217777 128175
rect 217811 128147 217839 128175
rect 217625 128085 217653 128113
rect 217687 128085 217715 128113
rect 217749 128085 217777 128113
rect 217811 128085 217839 128113
rect 217625 128023 217653 128051
rect 217687 128023 217715 128051
rect 217749 128023 217777 128051
rect 217811 128023 217839 128051
rect 217625 127961 217653 127989
rect 217687 127961 217715 127989
rect 217749 127961 217777 127989
rect 217811 127961 217839 127989
rect 217625 119147 217653 119175
rect 217687 119147 217715 119175
rect 217749 119147 217777 119175
rect 217811 119147 217839 119175
rect 217625 119085 217653 119113
rect 217687 119085 217715 119113
rect 217749 119085 217777 119113
rect 217811 119085 217839 119113
rect 217625 119023 217653 119051
rect 217687 119023 217715 119051
rect 217749 119023 217777 119051
rect 217811 119023 217839 119051
rect 217625 118961 217653 118989
rect 217687 118961 217715 118989
rect 217749 118961 217777 118989
rect 217811 118961 217839 118989
rect 217625 110147 217653 110175
rect 217687 110147 217715 110175
rect 217749 110147 217777 110175
rect 217811 110147 217839 110175
rect 217625 110085 217653 110113
rect 217687 110085 217715 110113
rect 217749 110085 217777 110113
rect 217811 110085 217839 110113
rect 217625 110023 217653 110051
rect 217687 110023 217715 110051
rect 217749 110023 217777 110051
rect 217811 110023 217839 110051
rect 217625 109961 217653 109989
rect 217687 109961 217715 109989
rect 217749 109961 217777 109989
rect 217811 109961 217839 109989
rect 217625 101147 217653 101175
rect 217687 101147 217715 101175
rect 217749 101147 217777 101175
rect 217811 101147 217839 101175
rect 217625 101085 217653 101113
rect 217687 101085 217715 101113
rect 217749 101085 217777 101113
rect 217811 101085 217839 101113
rect 217625 101023 217653 101051
rect 217687 101023 217715 101051
rect 217749 101023 217777 101051
rect 217811 101023 217839 101051
rect 217625 100961 217653 100989
rect 217687 100961 217715 100989
rect 217749 100961 217777 100989
rect 217811 100961 217839 100989
rect 217625 92147 217653 92175
rect 217687 92147 217715 92175
rect 217749 92147 217777 92175
rect 217811 92147 217839 92175
rect 217625 92085 217653 92113
rect 217687 92085 217715 92113
rect 217749 92085 217777 92113
rect 217811 92085 217839 92113
rect 217625 92023 217653 92051
rect 217687 92023 217715 92051
rect 217749 92023 217777 92051
rect 217811 92023 217839 92051
rect 217625 91961 217653 91989
rect 217687 91961 217715 91989
rect 217749 91961 217777 91989
rect 217811 91961 217839 91989
rect 217625 83147 217653 83175
rect 217687 83147 217715 83175
rect 217749 83147 217777 83175
rect 217811 83147 217839 83175
rect 217625 83085 217653 83113
rect 217687 83085 217715 83113
rect 217749 83085 217777 83113
rect 217811 83085 217839 83113
rect 217625 83023 217653 83051
rect 217687 83023 217715 83051
rect 217749 83023 217777 83051
rect 217811 83023 217839 83051
rect 217625 82961 217653 82989
rect 217687 82961 217715 82989
rect 217749 82961 217777 82989
rect 217811 82961 217839 82989
rect 217625 74147 217653 74175
rect 217687 74147 217715 74175
rect 217749 74147 217777 74175
rect 217811 74147 217839 74175
rect 217625 74085 217653 74113
rect 217687 74085 217715 74113
rect 217749 74085 217777 74113
rect 217811 74085 217839 74113
rect 217625 74023 217653 74051
rect 217687 74023 217715 74051
rect 217749 74023 217777 74051
rect 217811 74023 217839 74051
rect 217625 73961 217653 73989
rect 217687 73961 217715 73989
rect 217749 73961 217777 73989
rect 217811 73961 217839 73989
rect 217625 65147 217653 65175
rect 217687 65147 217715 65175
rect 217749 65147 217777 65175
rect 217811 65147 217839 65175
rect 217625 65085 217653 65113
rect 217687 65085 217715 65113
rect 217749 65085 217777 65113
rect 217811 65085 217839 65113
rect 217625 65023 217653 65051
rect 217687 65023 217715 65051
rect 217749 65023 217777 65051
rect 217811 65023 217839 65051
rect 217625 64961 217653 64989
rect 217687 64961 217715 64989
rect 217749 64961 217777 64989
rect 217811 64961 217839 64989
rect 217625 56147 217653 56175
rect 217687 56147 217715 56175
rect 217749 56147 217777 56175
rect 217811 56147 217839 56175
rect 217625 56085 217653 56113
rect 217687 56085 217715 56113
rect 217749 56085 217777 56113
rect 217811 56085 217839 56113
rect 217625 56023 217653 56051
rect 217687 56023 217715 56051
rect 217749 56023 217777 56051
rect 217811 56023 217839 56051
rect 217625 55961 217653 55989
rect 217687 55961 217715 55989
rect 217749 55961 217777 55989
rect 217811 55961 217839 55989
rect 217625 47147 217653 47175
rect 217687 47147 217715 47175
rect 217749 47147 217777 47175
rect 217811 47147 217839 47175
rect 217625 47085 217653 47113
rect 217687 47085 217715 47113
rect 217749 47085 217777 47113
rect 217811 47085 217839 47113
rect 217625 47023 217653 47051
rect 217687 47023 217715 47051
rect 217749 47023 217777 47051
rect 217811 47023 217839 47051
rect 217625 46961 217653 46989
rect 217687 46961 217715 46989
rect 217749 46961 217777 46989
rect 217811 46961 217839 46989
rect 217625 38147 217653 38175
rect 217687 38147 217715 38175
rect 217749 38147 217777 38175
rect 217811 38147 217839 38175
rect 217625 38085 217653 38113
rect 217687 38085 217715 38113
rect 217749 38085 217777 38113
rect 217811 38085 217839 38113
rect 217625 38023 217653 38051
rect 217687 38023 217715 38051
rect 217749 38023 217777 38051
rect 217811 38023 217839 38051
rect 217625 37961 217653 37989
rect 217687 37961 217715 37989
rect 217749 37961 217777 37989
rect 217811 37961 217839 37989
rect 217625 29147 217653 29175
rect 217687 29147 217715 29175
rect 217749 29147 217777 29175
rect 217811 29147 217839 29175
rect 217625 29085 217653 29113
rect 217687 29085 217715 29113
rect 217749 29085 217777 29113
rect 217811 29085 217839 29113
rect 217625 29023 217653 29051
rect 217687 29023 217715 29051
rect 217749 29023 217777 29051
rect 217811 29023 217839 29051
rect 217625 28961 217653 28989
rect 217687 28961 217715 28989
rect 217749 28961 217777 28989
rect 217811 28961 217839 28989
rect 217625 20147 217653 20175
rect 217687 20147 217715 20175
rect 217749 20147 217777 20175
rect 217811 20147 217839 20175
rect 217625 20085 217653 20113
rect 217687 20085 217715 20113
rect 217749 20085 217777 20113
rect 217811 20085 217839 20113
rect 217625 20023 217653 20051
rect 217687 20023 217715 20051
rect 217749 20023 217777 20051
rect 217811 20023 217839 20051
rect 217625 19961 217653 19989
rect 217687 19961 217715 19989
rect 217749 19961 217777 19989
rect 217811 19961 217839 19989
rect 217625 11147 217653 11175
rect 217687 11147 217715 11175
rect 217749 11147 217777 11175
rect 217811 11147 217839 11175
rect 217625 11085 217653 11113
rect 217687 11085 217715 11113
rect 217749 11085 217777 11113
rect 217811 11085 217839 11113
rect 217625 11023 217653 11051
rect 217687 11023 217715 11051
rect 217749 11023 217777 11051
rect 217811 11023 217839 11051
rect 217625 10961 217653 10989
rect 217687 10961 217715 10989
rect 217749 10961 217777 10989
rect 217811 10961 217839 10989
rect 217625 2147 217653 2175
rect 217687 2147 217715 2175
rect 217749 2147 217777 2175
rect 217811 2147 217839 2175
rect 217625 2085 217653 2113
rect 217687 2085 217715 2113
rect 217749 2085 217777 2113
rect 217811 2085 217839 2113
rect 217625 2023 217653 2051
rect 217687 2023 217715 2051
rect 217749 2023 217777 2051
rect 217811 2023 217839 2051
rect 217625 1961 217653 1989
rect 217687 1961 217715 1989
rect 217749 1961 217777 1989
rect 217811 1961 217839 1989
rect 217625 -108 217653 -80
rect 217687 -108 217715 -80
rect 217749 -108 217777 -80
rect 217811 -108 217839 -80
rect 217625 -170 217653 -142
rect 217687 -170 217715 -142
rect 217749 -170 217777 -142
rect 217811 -170 217839 -142
rect 217625 -232 217653 -204
rect 217687 -232 217715 -204
rect 217749 -232 217777 -204
rect 217811 -232 217839 -204
rect 217625 -294 217653 -266
rect 217687 -294 217715 -266
rect 217749 -294 217777 -266
rect 217811 -294 217839 -266
rect 219485 299058 219513 299086
rect 219547 299058 219575 299086
rect 219609 299058 219637 299086
rect 219671 299058 219699 299086
rect 219485 298996 219513 299024
rect 219547 298996 219575 299024
rect 219609 298996 219637 299024
rect 219671 298996 219699 299024
rect 219485 298934 219513 298962
rect 219547 298934 219575 298962
rect 219609 298934 219637 298962
rect 219671 298934 219699 298962
rect 219485 298872 219513 298900
rect 219547 298872 219575 298900
rect 219609 298872 219637 298900
rect 219671 298872 219699 298900
rect 219485 293147 219513 293175
rect 219547 293147 219575 293175
rect 219609 293147 219637 293175
rect 219671 293147 219699 293175
rect 219485 293085 219513 293113
rect 219547 293085 219575 293113
rect 219609 293085 219637 293113
rect 219671 293085 219699 293113
rect 219485 293023 219513 293051
rect 219547 293023 219575 293051
rect 219609 293023 219637 293051
rect 219671 293023 219699 293051
rect 219485 292961 219513 292989
rect 219547 292961 219575 292989
rect 219609 292961 219637 292989
rect 219671 292961 219699 292989
rect 219485 284147 219513 284175
rect 219547 284147 219575 284175
rect 219609 284147 219637 284175
rect 219671 284147 219699 284175
rect 219485 284085 219513 284113
rect 219547 284085 219575 284113
rect 219609 284085 219637 284113
rect 219671 284085 219699 284113
rect 219485 284023 219513 284051
rect 219547 284023 219575 284051
rect 219609 284023 219637 284051
rect 219671 284023 219699 284051
rect 219485 283961 219513 283989
rect 219547 283961 219575 283989
rect 219609 283961 219637 283989
rect 219671 283961 219699 283989
rect 219485 275147 219513 275175
rect 219547 275147 219575 275175
rect 219609 275147 219637 275175
rect 219671 275147 219699 275175
rect 219485 275085 219513 275113
rect 219547 275085 219575 275113
rect 219609 275085 219637 275113
rect 219671 275085 219699 275113
rect 219485 275023 219513 275051
rect 219547 275023 219575 275051
rect 219609 275023 219637 275051
rect 219671 275023 219699 275051
rect 219485 274961 219513 274989
rect 219547 274961 219575 274989
rect 219609 274961 219637 274989
rect 219671 274961 219699 274989
rect 219485 266147 219513 266175
rect 219547 266147 219575 266175
rect 219609 266147 219637 266175
rect 219671 266147 219699 266175
rect 219485 266085 219513 266113
rect 219547 266085 219575 266113
rect 219609 266085 219637 266113
rect 219671 266085 219699 266113
rect 219485 266023 219513 266051
rect 219547 266023 219575 266051
rect 219609 266023 219637 266051
rect 219671 266023 219699 266051
rect 219485 265961 219513 265989
rect 219547 265961 219575 265989
rect 219609 265961 219637 265989
rect 219671 265961 219699 265989
rect 219485 257147 219513 257175
rect 219547 257147 219575 257175
rect 219609 257147 219637 257175
rect 219671 257147 219699 257175
rect 219485 257085 219513 257113
rect 219547 257085 219575 257113
rect 219609 257085 219637 257113
rect 219671 257085 219699 257113
rect 219485 257023 219513 257051
rect 219547 257023 219575 257051
rect 219609 257023 219637 257051
rect 219671 257023 219699 257051
rect 219485 256961 219513 256989
rect 219547 256961 219575 256989
rect 219609 256961 219637 256989
rect 219671 256961 219699 256989
rect 219485 248147 219513 248175
rect 219547 248147 219575 248175
rect 219609 248147 219637 248175
rect 219671 248147 219699 248175
rect 219485 248085 219513 248113
rect 219547 248085 219575 248113
rect 219609 248085 219637 248113
rect 219671 248085 219699 248113
rect 219485 248023 219513 248051
rect 219547 248023 219575 248051
rect 219609 248023 219637 248051
rect 219671 248023 219699 248051
rect 219485 247961 219513 247989
rect 219547 247961 219575 247989
rect 219609 247961 219637 247989
rect 219671 247961 219699 247989
rect 219485 239147 219513 239175
rect 219547 239147 219575 239175
rect 219609 239147 219637 239175
rect 219671 239147 219699 239175
rect 219485 239085 219513 239113
rect 219547 239085 219575 239113
rect 219609 239085 219637 239113
rect 219671 239085 219699 239113
rect 219485 239023 219513 239051
rect 219547 239023 219575 239051
rect 219609 239023 219637 239051
rect 219671 239023 219699 239051
rect 219485 238961 219513 238989
rect 219547 238961 219575 238989
rect 219609 238961 219637 238989
rect 219671 238961 219699 238989
rect 219485 230147 219513 230175
rect 219547 230147 219575 230175
rect 219609 230147 219637 230175
rect 219671 230147 219699 230175
rect 219485 230085 219513 230113
rect 219547 230085 219575 230113
rect 219609 230085 219637 230113
rect 219671 230085 219699 230113
rect 219485 230023 219513 230051
rect 219547 230023 219575 230051
rect 219609 230023 219637 230051
rect 219671 230023 219699 230051
rect 219485 229961 219513 229989
rect 219547 229961 219575 229989
rect 219609 229961 219637 229989
rect 219671 229961 219699 229989
rect 219485 221147 219513 221175
rect 219547 221147 219575 221175
rect 219609 221147 219637 221175
rect 219671 221147 219699 221175
rect 219485 221085 219513 221113
rect 219547 221085 219575 221113
rect 219609 221085 219637 221113
rect 219671 221085 219699 221113
rect 219485 221023 219513 221051
rect 219547 221023 219575 221051
rect 219609 221023 219637 221051
rect 219671 221023 219699 221051
rect 219485 220961 219513 220989
rect 219547 220961 219575 220989
rect 219609 220961 219637 220989
rect 219671 220961 219699 220989
rect 219485 212147 219513 212175
rect 219547 212147 219575 212175
rect 219609 212147 219637 212175
rect 219671 212147 219699 212175
rect 219485 212085 219513 212113
rect 219547 212085 219575 212113
rect 219609 212085 219637 212113
rect 219671 212085 219699 212113
rect 219485 212023 219513 212051
rect 219547 212023 219575 212051
rect 219609 212023 219637 212051
rect 219671 212023 219699 212051
rect 219485 211961 219513 211989
rect 219547 211961 219575 211989
rect 219609 211961 219637 211989
rect 219671 211961 219699 211989
rect 219485 203147 219513 203175
rect 219547 203147 219575 203175
rect 219609 203147 219637 203175
rect 219671 203147 219699 203175
rect 219485 203085 219513 203113
rect 219547 203085 219575 203113
rect 219609 203085 219637 203113
rect 219671 203085 219699 203113
rect 219485 203023 219513 203051
rect 219547 203023 219575 203051
rect 219609 203023 219637 203051
rect 219671 203023 219699 203051
rect 219485 202961 219513 202989
rect 219547 202961 219575 202989
rect 219609 202961 219637 202989
rect 219671 202961 219699 202989
rect 219485 194147 219513 194175
rect 219547 194147 219575 194175
rect 219609 194147 219637 194175
rect 219671 194147 219699 194175
rect 219485 194085 219513 194113
rect 219547 194085 219575 194113
rect 219609 194085 219637 194113
rect 219671 194085 219699 194113
rect 219485 194023 219513 194051
rect 219547 194023 219575 194051
rect 219609 194023 219637 194051
rect 219671 194023 219699 194051
rect 219485 193961 219513 193989
rect 219547 193961 219575 193989
rect 219609 193961 219637 193989
rect 219671 193961 219699 193989
rect 219485 185147 219513 185175
rect 219547 185147 219575 185175
rect 219609 185147 219637 185175
rect 219671 185147 219699 185175
rect 219485 185085 219513 185113
rect 219547 185085 219575 185113
rect 219609 185085 219637 185113
rect 219671 185085 219699 185113
rect 219485 185023 219513 185051
rect 219547 185023 219575 185051
rect 219609 185023 219637 185051
rect 219671 185023 219699 185051
rect 219485 184961 219513 184989
rect 219547 184961 219575 184989
rect 219609 184961 219637 184989
rect 219671 184961 219699 184989
rect 219485 176147 219513 176175
rect 219547 176147 219575 176175
rect 219609 176147 219637 176175
rect 219671 176147 219699 176175
rect 219485 176085 219513 176113
rect 219547 176085 219575 176113
rect 219609 176085 219637 176113
rect 219671 176085 219699 176113
rect 219485 176023 219513 176051
rect 219547 176023 219575 176051
rect 219609 176023 219637 176051
rect 219671 176023 219699 176051
rect 219485 175961 219513 175989
rect 219547 175961 219575 175989
rect 219609 175961 219637 175989
rect 219671 175961 219699 175989
rect 219485 167147 219513 167175
rect 219547 167147 219575 167175
rect 219609 167147 219637 167175
rect 219671 167147 219699 167175
rect 219485 167085 219513 167113
rect 219547 167085 219575 167113
rect 219609 167085 219637 167113
rect 219671 167085 219699 167113
rect 219485 167023 219513 167051
rect 219547 167023 219575 167051
rect 219609 167023 219637 167051
rect 219671 167023 219699 167051
rect 219485 166961 219513 166989
rect 219547 166961 219575 166989
rect 219609 166961 219637 166989
rect 219671 166961 219699 166989
rect 219485 158147 219513 158175
rect 219547 158147 219575 158175
rect 219609 158147 219637 158175
rect 219671 158147 219699 158175
rect 219485 158085 219513 158113
rect 219547 158085 219575 158113
rect 219609 158085 219637 158113
rect 219671 158085 219699 158113
rect 219485 158023 219513 158051
rect 219547 158023 219575 158051
rect 219609 158023 219637 158051
rect 219671 158023 219699 158051
rect 219485 157961 219513 157989
rect 219547 157961 219575 157989
rect 219609 157961 219637 157989
rect 219671 157961 219699 157989
rect 219485 149147 219513 149175
rect 219547 149147 219575 149175
rect 219609 149147 219637 149175
rect 219671 149147 219699 149175
rect 219485 149085 219513 149113
rect 219547 149085 219575 149113
rect 219609 149085 219637 149113
rect 219671 149085 219699 149113
rect 219485 149023 219513 149051
rect 219547 149023 219575 149051
rect 219609 149023 219637 149051
rect 219671 149023 219699 149051
rect 219485 148961 219513 148989
rect 219547 148961 219575 148989
rect 219609 148961 219637 148989
rect 219671 148961 219699 148989
rect 219485 140147 219513 140175
rect 219547 140147 219575 140175
rect 219609 140147 219637 140175
rect 219671 140147 219699 140175
rect 219485 140085 219513 140113
rect 219547 140085 219575 140113
rect 219609 140085 219637 140113
rect 219671 140085 219699 140113
rect 219485 140023 219513 140051
rect 219547 140023 219575 140051
rect 219609 140023 219637 140051
rect 219671 140023 219699 140051
rect 219485 139961 219513 139989
rect 219547 139961 219575 139989
rect 219609 139961 219637 139989
rect 219671 139961 219699 139989
rect 219485 131147 219513 131175
rect 219547 131147 219575 131175
rect 219609 131147 219637 131175
rect 219671 131147 219699 131175
rect 219485 131085 219513 131113
rect 219547 131085 219575 131113
rect 219609 131085 219637 131113
rect 219671 131085 219699 131113
rect 219485 131023 219513 131051
rect 219547 131023 219575 131051
rect 219609 131023 219637 131051
rect 219671 131023 219699 131051
rect 219485 130961 219513 130989
rect 219547 130961 219575 130989
rect 219609 130961 219637 130989
rect 219671 130961 219699 130989
rect 219485 122147 219513 122175
rect 219547 122147 219575 122175
rect 219609 122147 219637 122175
rect 219671 122147 219699 122175
rect 219485 122085 219513 122113
rect 219547 122085 219575 122113
rect 219609 122085 219637 122113
rect 219671 122085 219699 122113
rect 219485 122023 219513 122051
rect 219547 122023 219575 122051
rect 219609 122023 219637 122051
rect 219671 122023 219699 122051
rect 219485 121961 219513 121989
rect 219547 121961 219575 121989
rect 219609 121961 219637 121989
rect 219671 121961 219699 121989
rect 219485 113147 219513 113175
rect 219547 113147 219575 113175
rect 219609 113147 219637 113175
rect 219671 113147 219699 113175
rect 219485 113085 219513 113113
rect 219547 113085 219575 113113
rect 219609 113085 219637 113113
rect 219671 113085 219699 113113
rect 219485 113023 219513 113051
rect 219547 113023 219575 113051
rect 219609 113023 219637 113051
rect 219671 113023 219699 113051
rect 219485 112961 219513 112989
rect 219547 112961 219575 112989
rect 219609 112961 219637 112989
rect 219671 112961 219699 112989
rect 219485 104147 219513 104175
rect 219547 104147 219575 104175
rect 219609 104147 219637 104175
rect 219671 104147 219699 104175
rect 219485 104085 219513 104113
rect 219547 104085 219575 104113
rect 219609 104085 219637 104113
rect 219671 104085 219699 104113
rect 219485 104023 219513 104051
rect 219547 104023 219575 104051
rect 219609 104023 219637 104051
rect 219671 104023 219699 104051
rect 219485 103961 219513 103989
rect 219547 103961 219575 103989
rect 219609 103961 219637 103989
rect 219671 103961 219699 103989
rect 219485 95147 219513 95175
rect 219547 95147 219575 95175
rect 219609 95147 219637 95175
rect 219671 95147 219699 95175
rect 219485 95085 219513 95113
rect 219547 95085 219575 95113
rect 219609 95085 219637 95113
rect 219671 95085 219699 95113
rect 219485 95023 219513 95051
rect 219547 95023 219575 95051
rect 219609 95023 219637 95051
rect 219671 95023 219699 95051
rect 219485 94961 219513 94989
rect 219547 94961 219575 94989
rect 219609 94961 219637 94989
rect 219671 94961 219699 94989
rect 219485 86147 219513 86175
rect 219547 86147 219575 86175
rect 219609 86147 219637 86175
rect 219671 86147 219699 86175
rect 219485 86085 219513 86113
rect 219547 86085 219575 86113
rect 219609 86085 219637 86113
rect 219671 86085 219699 86113
rect 219485 86023 219513 86051
rect 219547 86023 219575 86051
rect 219609 86023 219637 86051
rect 219671 86023 219699 86051
rect 219485 85961 219513 85989
rect 219547 85961 219575 85989
rect 219609 85961 219637 85989
rect 219671 85961 219699 85989
rect 219485 77147 219513 77175
rect 219547 77147 219575 77175
rect 219609 77147 219637 77175
rect 219671 77147 219699 77175
rect 219485 77085 219513 77113
rect 219547 77085 219575 77113
rect 219609 77085 219637 77113
rect 219671 77085 219699 77113
rect 219485 77023 219513 77051
rect 219547 77023 219575 77051
rect 219609 77023 219637 77051
rect 219671 77023 219699 77051
rect 219485 76961 219513 76989
rect 219547 76961 219575 76989
rect 219609 76961 219637 76989
rect 219671 76961 219699 76989
rect 219485 68147 219513 68175
rect 219547 68147 219575 68175
rect 219609 68147 219637 68175
rect 219671 68147 219699 68175
rect 219485 68085 219513 68113
rect 219547 68085 219575 68113
rect 219609 68085 219637 68113
rect 219671 68085 219699 68113
rect 219485 68023 219513 68051
rect 219547 68023 219575 68051
rect 219609 68023 219637 68051
rect 219671 68023 219699 68051
rect 219485 67961 219513 67989
rect 219547 67961 219575 67989
rect 219609 67961 219637 67989
rect 219671 67961 219699 67989
rect 219485 59147 219513 59175
rect 219547 59147 219575 59175
rect 219609 59147 219637 59175
rect 219671 59147 219699 59175
rect 219485 59085 219513 59113
rect 219547 59085 219575 59113
rect 219609 59085 219637 59113
rect 219671 59085 219699 59113
rect 219485 59023 219513 59051
rect 219547 59023 219575 59051
rect 219609 59023 219637 59051
rect 219671 59023 219699 59051
rect 219485 58961 219513 58989
rect 219547 58961 219575 58989
rect 219609 58961 219637 58989
rect 219671 58961 219699 58989
rect 219485 50147 219513 50175
rect 219547 50147 219575 50175
rect 219609 50147 219637 50175
rect 219671 50147 219699 50175
rect 219485 50085 219513 50113
rect 219547 50085 219575 50113
rect 219609 50085 219637 50113
rect 219671 50085 219699 50113
rect 219485 50023 219513 50051
rect 219547 50023 219575 50051
rect 219609 50023 219637 50051
rect 219671 50023 219699 50051
rect 219485 49961 219513 49989
rect 219547 49961 219575 49989
rect 219609 49961 219637 49989
rect 219671 49961 219699 49989
rect 219485 41147 219513 41175
rect 219547 41147 219575 41175
rect 219609 41147 219637 41175
rect 219671 41147 219699 41175
rect 219485 41085 219513 41113
rect 219547 41085 219575 41113
rect 219609 41085 219637 41113
rect 219671 41085 219699 41113
rect 219485 41023 219513 41051
rect 219547 41023 219575 41051
rect 219609 41023 219637 41051
rect 219671 41023 219699 41051
rect 219485 40961 219513 40989
rect 219547 40961 219575 40989
rect 219609 40961 219637 40989
rect 219671 40961 219699 40989
rect 219485 32147 219513 32175
rect 219547 32147 219575 32175
rect 219609 32147 219637 32175
rect 219671 32147 219699 32175
rect 219485 32085 219513 32113
rect 219547 32085 219575 32113
rect 219609 32085 219637 32113
rect 219671 32085 219699 32113
rect 219485 32023 219513 32051
rect 219547 32023 219575 32051
rect 219609 32023 219637 32051
rect 219671 32023 219699 32051
rect 219485 31961 219513 31989
rect 219547 31961 219575 31989
rect 219609 31961 219637 31989
rect 219671 31961 219699 31989
rect 219485 23147 219513 23175
rect 219547 23147 219575 23175
rect 219609 23147 219637 23175
rect 219671 23147 219699 23175
rect 219485 23085 219513 23113
rect 219547 23085 219575 23113
rect 219609 23085 219637 23113
rect 219671 23085 219699 23113
rect 219485 23023 219513 23051
rect 219547 23023 219575 23051
rect 219609 23023 219637 23051
rect 219671 23023 219699 23051
rect 219485 22961 219513 22989
rect 219547 22961 219575 22989
rect 219609 22961 219637 22989
rect 219671 22961 219699 22989
rect 219485 14147 219513 14175
rect 219547 14147 219575 14175
rect 219609 14147 219637 14175
rect 219671 14147 219699 14175
rect 219485 14085 219513 14113
rect 219547 14085 219575 14113
rect 219609 14085 219637 14113
rect 219671 14085 219699 14113
rect 219485 14023 219513 14051
rect 219547 14023 219575 14051
rect 219609 14023 219637 14051
rect 219671 14023 219699 14051
rect 219485 13961 219513 13989
rect 219547 13961 219575 13989
rect 219609 13961 219637 13989
rect 219671 13961 219699 13989
rect 219485 5147 219513 5175
rect 219547 5147 219575 5175
rect 219609 5147 219637 5175
rect 219671 5147 219699 5175
rect 219485 5085 219513 5113
rect 219547 5085 219575 5113
rect 219609 5085 219637 5113
rect 219671 5085 219699 5113
rect 219485 5023 219513 5051
rect 219547 5023 219575 5051
rect 219609 5023 219637 5051
rect 219671 5023 219699 5051
rect 219485 4961 219513 4989
rect 219547 4961 219575 4989
rect 219609 4961 219637 4989
rect 219671 4961 219699 4989
rect 219485 -588 219513 -560
rect 219547 -588 219575 -560
rect 219609 -588 219637 -560
rect 219671 -588 219699 -560
rect 219485 -650 219513 -622
rect 219547 -650 219575 -622
rect 219609 -650 219637 -622
rect 219671 -650 219699 -622
rect 219485 -712 219513 -684
rect 219547 -712 219575 -684
rect 219609 -712 219637 -684
rect 219671 -712 219699 -684
rect 219485 -774 219513 -746
rect 219547 -774 219575 -746
rect 219609 -774 219637 -746
rect 219671 -774 219699 -746
rect 226625 298578 226653 298606
rect 226687 298578 226715 298606
rect 226749 298578 226777 298606
rect 226811 298578 226839 298606
rect 226625 298516 226653 298544
rect 226687 298516 226715 298544
rect 226749 298516 226777 298544
rect 226811 298516 226839 298544
rect 226625 298454 226653 298482
rect 226687 298454 226715 298482
rect 226749 298454 226777 298482
rect 226811 298454 226839 298482
rect 226625 298392 226653 298420
rect 226687 298392 226715 298420
rect 226749 298392 226777 298420
rect 226811 298392 226839 298420
rect 226625 290147 226653 290175
rect 226687 290147 226715 290175
rect 226749 290147 226777 290175
rect 226811 290147 226839 290175
rect 226625 290085 226653 290113
rect 226687 290085 226715 290113
rect 226749 290085 226777 290113
rect 226811 290085 226839 290113
rect 226625 290023 226653 290051
rect 226687 290023 226715 290051
rect 226749 290023 226777 290051
rect 226811 290023 226839 290051
rect 226625 289961 226653 289989
rect 226687 289961 226715 289989
rect 226749 289961 226777 289989
rect 226811 289961 226839 289989
rect 226625 281147 226653 281175
rect 226687 281147 226715 281175
rect 226749 281147 226777 281175
rect 226811 281147 226839 281175
rect 226625 281085 226653 281113
rect 226687 281085 226715 281113
rect 226749 281085 226777 281113
rect 226811 281085 226839 281113
rect 226625 281023 226653 281051
rect 226687 281023 226715 281051
rect 226749 281023 226777 281051
rect 226811 281023 226839 281051
rect 226625 280961 226653 280989
rect 226687 280961 226715 280989
rect 226749 280961 226777 280989
rect 226811 280961 226839 280989
rect 226625 272147 226653 272175
rect 226687 272147 226715 272175
rect 226749 272147 226777 272175
rect 226811 272147 226839 272175
rect 226625 272085 226653 272113
rect 226687 272085 226715 272113
rect 226749 272085 226777 272113
rect 226811 272085 226839 272113
rect 226625 272023 226653 272051
rect 226687 272023 226715 272051
rect 226749 272023 226777 272051
rect 226811 272023 226839 272051
rect 226625 271961 226653 271989
rect 226687 271961 226715 271989
rect 226749 271961 226777 271989
rect 226811 271961 226839 271989
rect 226625 263147 226653 263175
rect 226687 263147 226715 263175
rect 226749 263147 226777 263175
rect 226811 263147 226839 263175
rect 226625 263085 226653 263113
rect 226687 263085 226715 263113
rect 226749 263085 226777 263113
rect 226811 263085 226839 263113
rect 226625 263023 226653 263051
rect 226687 263023 226715 263051
rect 226749 263023 226777 263051
rect 226811 263023 226839 263051
rect 226625 262961 226653 262989
rect 226687 262961 226715 262989
rect 226749 262961 226777 262989
rect 226811 262961 226839 262989
rect 226625 254147 226653 254175
rect 226687 254147 226715 254175
rect 226749 254147 226777 254175
rect 226811 254147 226839 254175
rect 226625 254085 226653 254113
rect 226687 254085 226715 254113
rect 226749 254085 226777 254113
rect 226811 254085 226839 254113
rect 226625 254023 226653 254051
rect 226687 254023 226715 254051
rect 226749 254023 226777 254051
rect 226811 254023 226839 254051
rect 226625 253961 226653 253989
rect 226687 253961 226715 253989
rect 226749 253961 226777 253989
rect 226811 253961 226839 253989
rect 226625 245147 226653 245175
rect 226687 245147 226715 245175
rect 226749 245147 226777 245175
rect 226811 245147 226839 245175
rect 226625 245085 226653 245113
rect 226687 245085 226715 245113
rect 226749 245085 226777 245113
rect 226811 245085 226839 245113
rect 226625 245023 226653 245051
rect 226687 245023 226715 245051
rect 226749 245023 226777 245051
rect 226811 245023 226839 245051
rect 226625 244961 226653 244989
rect 226687 244961 226715 244989
rect 226749 244961 226777 244989
rect 226811 244961 226839 244989
rect 226625 236147 226653 236175
rect 226687 236147 226715 236175
rect 226749 236147 226777 236175
rect 226811 236147 226839 236175
rect 226625 236085 226653 236113
rect 226687 236085 226715 236113
rect 226749 236085 226777 236113
rect 226811 236085 226839 236113
rect 226625 236023 226653 236051
rect 226687 236023 226715 236051
rect 226749 236023 226777 236051
rect 226811 236023 226839 236051
rect 226625 235961 226653 235989
rect 226687 235961 226715 235989
rect 226749 235961 226777 235989
rect 226811 235961 226839 235989
rect 226625 227147 226653 227175
rect 226687 227147 226715 227175
rect 226749 227147 226777 227175
rect 226811 227147 226839 227175
rect 226625 227085 226653 227113
rect 226687 227085 226715 227113
rect 226749 227085 226777 227113
rect 226811 227085 226839 227113
rect 226625 227023 226653 227051
rect 226687 227023 226715 227051
rect 226749 227023 226777 227051
rect 226811 227023 226839 227051
rect 226625 226961 226653 226989
rect 226687 226961 226715 226989
rect 226749 226961 226777 226989
rect 226811 226961 226839 226989
rect 226625 218147 226653 218175
rect 226687 218147 226715 218175
rect 226749 218147 226777 218175
rect 226811 218147 226839 218175
rect 226625 218085 226653 218113
rect 226687 218085 226715 218113
rect 226749 218085 226777 218113
rect 226811 218085 226839 218113
rect 226625 218023 226653 218051
rect 226687 218023 226715 218051
rect 226749 218023 226777 218051
rect 226811 218023 226839 218051
rect 226625 217961 226653 217989
rect 226687 217961 226715 217989
rect 226749 217961 226777 217989
rect 226811 217961 226839 217989
rect 226625 209147 226653 209175
rect 226687 209147 226715 209175
rect 226749 209147 226777 209175
rect 226811 209147 226839 209175
rect 226625 209085 226653 209113
rect 226687 209085 226715 209113
rect 226749 209085 226777 209113
rect 226811 209085 226839 209113
rect 226625 209023 226653 209051
rect 226687 209023 226715 209051
rect 226749 209023 226777 209051
rect 226811 209023 226839 209051
rect 226625 208961 226653 208989
rect 226687 208961 226715 208989
rect 226749 208961 226777 208989
rect 226811 208961 226839 208989
rect 226625 200147 226653 200175
rect 226687 200147 226715 200175
rect 226749 200147 226777 200175
rect 226811 200147 226839 200175
rect 226625 200085 226653 200113
rect 226687 200085 226715 200113
rect 226749 200085 226777 200113
rect 226811 200085 226839 200113
rect 226625 200023 226653 200051
rect 226687 200023 226715 200051
rect 226749 200023 226777 200051
rect 226811 200023 226839 200051
rect 226625 199961 226653 199989
rect 226687 199961 226715 199989
rect 226749 199961 226777 199989
rect 226811 199961 226839 199989
rect 226625 191147 226653 191175
rect 226687 191147 226715 191175
rect 226749 191147 226777 191175
rect 226811 191147 226839 191175
rect 226625 191085 226653 191113
rect 226687 191085 226715 191113
rect 226749 191085 226777 191113
rect 226811 191085 226839 191113
rect 226625 191023 226653 191051
rect 226687 191023 226715 191051
rect 226749 191023 226777 191051
rect 226811 191023 226839 191051
rect 226625 190961 226653 190989
rect 226687 190961 226715 190989
rect 226749 190961 226777 190989
rect 226811 190961 226839 190989
rect 226625 182147 226653 182175
rect 226687 182147 226715 182175
rect 226749 182147 226777 182175
rect 226811 182147 226839 182175
rect 226625 182085 226653 182113
rect 226687 182085 226715 182113
rect 226749 182085 226777 182113
rect 226811 182085 226839 182113
rect 226625 182023 226653 182051
rect 226687 182023 226715 182051
rect 226749 182023 226777 182051
rect 226811 182023 226839 182051
rect 226625 181961 226653 181989
rect 226687 181961 226715 181989
rect 226749 181961 226777 181989
rect 226811 181961 226839 181989
rect 226625 173147 226653 173175
rect 226687 173147 226715 173175
rect 226749 173147 226777 173175
rect 226811 173147 226839 173175
rect 226625 173085 226653 173113
rect 226687 173085 226715 173113
rect 226749 173085 226777 173113
rect 226811 173085 226839 173113
rect 226625 173023 226653 173051
rect 226687 173023 226715 173051
rect 226749 173023 226777 173051
rect 226811 173023 226839 173051
rect 226625 172961 226653 172989
rect 226687 172961 226715 172989
rect 226749 172961 226777 172989
rect 226811 172961 226839 172989
rect 226625 164147 226653 164175
rect 226687 164147 226715 164175
rect 226749 164147 226777 164175
rect 226811 164147 226839 164175
rect 226625 164085 226653 164113
rect 226687 164085 226715 164113
rect 226749 164085 226777 164113
rect 226811 164085 226839 164113
rect 226625 164023 226653 164051
rect 226687 164023 226715 164051
rect 226749 164023 226777 164051
rect 226811 164023 226839 164051
rect 226625 163961 226653 163989
rect 226687 163961 226715 163989
rect 226749 163961 226777 163989
rect 226811 163961 226839 163989
rect 226625 155147 226653 155175
rect 226687 155147 226715 155175
rect 226749 155147 226777 155175
rect 226811 155147 226839 155175
rect 226625 155085 226653 155113
rect 226687 155085 226715 155113
rect 226749 155085 226777 155113
rect 226811 155085 226839 155113
rect 226625 155023 226653 155051
rect 226687 155023 226715 155051
rect 226749 155023 226777 155051
rect 226811 155023 226839 155051
rect 226625 154961 226653 154989
rect 226687 154961 226715 154989
rect 226749 154961 226777 154989
rect 226811 154961 226839 154989
rect 226625 146147 226653 146175
rect 226687 146147 226715 146175
rect 226749 146147 226777 146175
rect 226811 146147 226839 146175
rect 226625 146085 226653 146113
rect 226687 146085 226715 146113
rect 226749 146085 226777 146113
rect 226811 146085 226839 146113
rect 226625 146023 226653 146051
rect 226687 146023 226715 146051
rect 226749 146023 226777 146051
rect 226811 146023 226839 146051
rect 226625 145961 226653 145989
rect 226687 145961 226715 145989
rect 226749 145961 226777 145989
rect 226811 145961 226839 145989
rect 226625 137147 226653 137175
rect 226687 137147 226715 137175
rect 226749 137147 226777 137175
rect 226811 137147 226839 137175
rect 226625 137085 226653 137113
rect 226687 137085 226715 137113
rect 226749 137085 226777 137113
rect 226811 137085 226839 137113
rect 226625 137023 226653 137051
rect 226687 137023 226715 137051
rect 226749 137023 226777 137051
rect 226811 137023 226839 137051
rect 226625 136961 226653 136989
rect 226687 136961 226715 136989
rect 226749 136961 226777 136989
rect 226811 136961 226839 136989
rect 226625 128147 226653 128175
rect 226687 128147 226715 128175
rect 226749 128147 226777 128175
rect 226811 128147 226839 128175
rect 226625 128085 226653 128113
rect 226687 128085 226715 128113
rect 226749 128085 226777 128113
rect 226811 128085 226839 128113
rect 226625 128023 226653 128051
rect 226687 128023 226715 128051
rect 226749 128023 226777 128051
rect 226811 128023 226839 128051
rect 226625 127961 226653 127989
rect 226687 127961 226715 127989
rect 226749 127961 226777 127989
rect 226811 127961 226839 127989
rect 226625 119147 226653 119175
rect 226687 119147 226715 119175
rect 226749 119147 226777 119175
rect 226811 119147 226839 119175
rect 226625 119085 226653 119113
rect 226687 119085 226715 119113
rect 226749 119085 226777 119113
rect 226811 119085 226839 119113
rect 226625 119023 226653 119051
rect 226687 119023 226715 119051
rect 226749 119023 226777 119051
rect 226811 119023 226839 119051
rect 226625 118961 226653 118989
rect 226687 118961 226715 118989
rect 226749 118961 226777 118989
rect 226811 118961 226839 118989
rect 226625 110147 226653 110175
rect 226687 110147 226715 110175
rect 226749 110147 226777 110175
rect 226811 110147 226839 110175
rect 226625 110085 226653 110113
rect 226687 110085 226715 110113
rect 226749 110085 226777 110113
rect 226811 110085 226839 110113
rect 226625 110023 226653 110051
rect 226687 110023 226715 110051
rect 226749 110023 226777 110051
rect 226811 110023 226839 110051
rect 226625 109961 226653 109989
rect 226687 109961 226715 109989
rect 226749 109961 226777 109989
rect 226811 109961 226839 109989
rect 226625 101147 226653 101175
rect 226687 101147 226715 101175
rect 226749 101147 226777 101175
rect 226811 101147 226839 101175
rect 226625 101085 226653 101113
rect 226687 101085 226715 101113
rect 226749 101085 226777 101113
rect 226811 101085 226839 101113
rect 226625 101023 226653 101051
rect 226687 101023 226715 101051
rect 226749 101023 226777 101051
rect 226811 101023 226839 101051
rect 226625 100961 226653 100989
rect 226687 100961 226715 100989
rect 226749 100961 226777 100989
rect 226811 100961 226839 100989
rect 226625 92147 226653 92175
rect 226687 92147 226715 92175
rect 226749 92147 226777 92175
rect 226811 92147 226839 92175
rect 226625 92085 226653 92113
rect 226687 92085 226715 92113
rect 226749 92085 226777 92113
rect 226811 92085 226839 92113
rect 226625 92023 226653 92051
rect 226687 92023 226715 92051
rect 226749 92023 226777 92051
rect 226811 92023 226839 92051
rect 226625 91961 226653 91989
rect 226687 91961 226715 91989
rect 226749 91961 226777 91989
rect 226811 91961 226839 91989
rect 226625 83147 226653 83175
rect 226687 83147 226715 83175
rect 226749 83147 226777 83175
rect 226811 83147 226839 83175
rect 226625 83085 226653 83113
rect 226687 83085 226715 83113
rect 226749 83085 226777 83113
rect 226811 83085 226839 83113
rect 226625 83023 226653 83051
rect 226687 83023 226715 83051
rect 226749 83023 226777 83051
rect 226811 83023 226839 83051
rect 226625 82961 226653 82989
rect 226687 82961 226715 82989
rect 226749 82961 226777 82989
rect 226811 82961 226839 82989
rect 226625 74147 226653 74175
rect 226687 74147 226715 74175
rect 226749 74147 226777 74175
rect 226811 74147 226839 74175
rect 226625 74085 226653 74113
rect 226687 74085 226715 74113
rect 226749 74085 226777 74113
rect 226811 74085 226839 74113
rect 226625 74023 226653 74051
rect 226687 74023 226715 74051
rect 226749 74023 226777 74051
rect 226811 74023 226839 74051
rect 226625 73961 226653 73989
rect 226687 73961 226715 73989
rect 226749 73961 226777 73989
rect 226811 73961 226839 73989
rect 226625 65147 226653 65175
rect 226687 65147 226715 65175
rect 226749 65147 226777 65175
rect 226811 65147 226839 65175
rect 226625 65085 226653 65113
rect 226687 65085 226715 65113
rect 226749 65085 226777 65113
rect 226811 65085 226839 65113
rect 226625 65023 226653 65051
rect 226687 65023 226715 65051
rect 226749 65023 226777 65051
rect 226811 65023 226839 65051
rect 226625 64961 226653 64989
rect 226687 64961 226715 64989
rect 226749 64961 226777 64989
rect 226811 64961 226839 64989
rect 226625 56147 226653 56175
rect 226687 56147 226715 56175
rect 226749 56147 226777 56175
rect 226811 56147 226839 56175
rect 226625 56085 226653 56113
rect 226687 56085 226715 56113
rect 226749 56085 226777 56113
rect 226811 56085 226839 56113
rect 226625 56023 226653 56051
rect 226687 56023 226715 56051
rect 226749 56023 226777 56051
rect 226811 56023 226839 56051
rect 226625 55961 226653 55989
rect 226687 55961 226715 55989
rect 226749 55961 226777 55989
rect 226811 55961 226839 55989
rect 226625 47147 226653 47175
rect 226687 47147 226715 47175
rect 226749 47147 226777 47175
rect 226811 47147 226839 47175
rect 226625 47085 226653 47113
rect 226687 47085 226715 47113
rect 226749 47085 226777 47113
rect 226811 47085 226839 47113
rect 226625 47023 226653 47051
rect 226687 47023 226715 47051
rect 226749 47023 226777 47051
rect 226811 47023 226839 47051
rect 226625 46961 226653 46989
rect 226687 46961 226715 46989
rect 226749 46961 226777 46989
rect 226811 46961 226839 46989
rect 226625 38147 226653 38175
rect 226687 38147 226715 38175
rect 226749 38147 226777 38175
rect 226811 38147 226839 38175
rect 226625 38085 226653 38113
rect 226687 38085 226715 38113
rect 226749 38085 226777 38113
rect 226811 38085 226839 38113
rect 226625 38023 226653 38051
rect 226687 38023 226715 38051
rect 226749 38023 226777 38051
rect 226811 38023 226839 38051
rect 226625 37961 226653 37989
rect 226687 37961 226715 37989
rect 226749 37961 226777 37989
rect 226811 37961 226839 37989
rect 226625 29147 226653 29175
rect 226687 29147 226715 29175
rect 226749 29147 226777 29175
rect 226811 29147 226839 29175
rect 226625 29085 226653 29113
rect 226687 29085 226715 29113
rect 226749 29085 226777 29113
rect 226811 29085 226839 29113
rect 226625 29023 226653 29051
rect 226687 29023 226715 29051
rect 226749 29023 226777 29051
rect 226811 29023 226839 29051
rect 226625 28961 226653 28989
rect 226687 28961 226715 28989
rect 226749 28961 226777 28989
rect 226811 28961 226839 28989
rect 226625 20147 226653 20175
rect 226687 20147 226715 20175
rect 226749 20147 226777 20175
rect 226811 20147 226839 20175
rect 226625 20085 226653 20113
rect 226687 20085 226715 20113
rect 226749 20085 226777 20113
rect 226811 20085 226839 20113
rect 226625 20023 226653 20051
rect 226687 20023 226715 20051
rect 226749 20023 226777 20051
rect 226811 20023 226839 20051
rect 226625 19961 226653 19989
rect 226687 19961 226715 19989
rect 226749 19961 226777 19989
rect 226811 19961 226839 19989
rect 226625 11147 226653 11175
rect 226687 11147 226715 11175
rect 226749 11147 226777 11175
rect 226811 11147 226839 11175
rect 226625 11085 226653 11113
rect 226687 11085 226715 11113
rect 226749 11085 226777 11113
rect 226811 11085 226839 11113
rect 226625 11023 226653 11051
rect 226687 11023 226715 11051
rect 226749 11023 226777 11051
rect 226811 11023 226839 11051
rect 226625 10961 226653 10989
rect 226687 10961 226715 10989
rect 226749 10961 226777 10989
rect 226811 10961 226839 10989
rect 226625 2147 226653 2175
rect 226687 2147 226715 2175
rect 226749 2147 226777 2175
rect 226811 2147 226839 2175
rect 226625 2085 226653 2113
rect 226687 2085 226715 2113
rect 226749 2085 226777 2113
rect 226811 2085 226839 2113
rect 226625 2023 226653 2051
rect 226687 2023 226715 2051
rect 226749 2023 226777 2051
rect 226811 2023 226839 2051
rect 226625 1961 226653 1989
rect 226687 1961 226715 1989
rect 226749 1961 226777 1989
rect 226811 1961 226839 1989
rect 226625 -108 226653 -80
rect 226687 -108 226715 -80
rect 226749 -108 226777 -80
rect 226811 -108 226839 -80
rect 226625 -170 226653 -142
rect 226687 -170 226715 -142
rect 226749 -170 226777 -142
rect 226811 -170 226839 -142
rect 226625 -232 226653 -204
rect 226687 -232 226715 -204
rect 226749 -232 226777 -204
rect 226811 -232 226839 -204
rect 226625 -294 226653 -266
rect 226687 -294 226715 -266
rect 226749 -294 226777 -266
rect 226811 -294 226839 -266
rect 228485 299058 228513 299086
rect 228547 299058 228575 299086
rect 228609 299058 228637 299086
rect 228671 299058 228699 299086
rect 228485 298996 228513 299024
rect 228547 298996 228575 299024
rect 228609 298996 228637 299024
rect 228671 298996 228699 299024
rect 228485 298934 228513 298962
rect 228547 298934 228575 298962
rect 228609 298934 228637 298962
rect 228671 298934 228699 298962
rect 228485 298872 228513 298900
rect 228547 298872 228575 298900
rect 228609 298872 228637 298900
rect 228671 298872 228699 298900
rect 228485 293147 228513 293175
rect 228547 293147 228575 293175
rect 228609 293147 228637 293175
rect 228671 293147 228699 293175
rect 228485 293085 228513 293113
rect 228547 293085 228575 293113
rect 228609 293085 228637 293113
rect 228671 293085 228699 293113
rect 228485 293023 228513 293051
rect 228547 293023 228575 293051
rect 228609 293023 228637 293051
rect 228671 293023 228699 293051
rect 228485 292961 228513 292989
rect 228547 292961 228575 292989
rect 228609 292961 228637 292989
rect 228671 292961 228699 292989
rect 228485 284147 228513 284175
rect 228547 284147 228575 284175
rect 228609 284147 228637 284175
rect 228671 284147 228699 284175
rect 228485 284085 228513 284113
rect 228547 284085 228575 284113
rect 228609 284085 228637 284113
rect 228671 284085 228699 284113
rect 228485 284023 228513 284051
rect 228547 284023 228575 284051
rect 228609 284023 228637 284051
rect 228671 284023 228699 284051
rect 228485 283961 228513 283989
rect 228547 283961 228575 283989
rect 228609 283961 228637 283989
rect 228671 283961 228699 283989
rect 228485 275147 228513 275175
rect 228547 275147 228575 275175
rect 228609 275147 228637 275175
rect 228671 275147 228699 275175
rect 228485 275085 228513 275113
rect 228547 275085 228575 275113
rect 228609 275085 228637 275113
rect 228671 275085 228699 275113
rect 228485 275023 228513 275051
rect 228547 275023 228575 275051
rect 228609 275023 228637 275051
rect 228671 275023 228699 275051
rect 228485 274961 228513 274989
rect 228547 274961 228575 274989
rect 228609 274961 228637 274989
rect 228671 274961 228699 274989
rect 228485 266147 228513 266175
rect 228547 266147 228575 266175
rect 228609 266147 228637 266175
rect 228671 266147 228699 266175
rect 228485 266085 228513 266113
rect 228547 266085 228575 266113
rect 228609 266085 228637 266113
rect 228671 266085 228699 266113
rect 228485 266023 228513 266051
rect 228547 266023 228575 266051
rect 228609 266023 228637 266051
rect 228671 266023 228699 266051
rect 228485 265961 228513 265989
rect 228547 265961 228575 265989
rect 228609 265961 228637 265989
rect 228671 265961 228699 265989
rect 228485 257147 228513 257175
rect 228547 257147 228575 257175
rect 228609 257147 228637 257175
rect 228671 257147 228699 257175
rect 228485 257085 228513 257113
rect 228547 257085 228575 257113
rect 228609 257085 228637 257113
rect 228671 257085 228699 257113
rect 228485 257023 228513 257051
rect 228547 257023 228575 257051
rect 228609 257023 228637 257051
rect 228671 257023 228699 257051
rect 228485 256961 228513 256989
rect 228547 256961 228575 256989
rect 228609 256961 228637 256989
rect 228671 256961 228699 256989
rect 228485 248147 228513 248175
rect 228547 248147 228575 248175
rect 228609 248147 228637 248175
rect 228671 248147 228699 248175
rect 228485 248085 228513 248113
rect 228547 248085 228575 248113
rect 228609 248085 228637 248113
rect 228671 248085 228699 248113
rect 228485 248023 228513 248051
rect 228547 248023 228575 248051
rect 228609 248023 228637 248051
rect 228671 248023 228699 248051
rect 228485 247961 228513 247989
rect 228547 247961 228575 247989
rect 228609 247961 228637 247989
rect 228671 247961 228699 247989
rect 228485 239147 228513 239175
rect 228547 239147 228575 239175
rect 228609 239147 228637 239175
rect 228671 239147 228699 239175
rect 228485 239085 228513 239113
rect 228547 239085 228575 239113
rect 228609 239085 228637 239113
rect 228671 239085 228699 239113
rect 228485 239023 228513 239051
rect 228547 239023 228575 239051
rect 228609 239023 228637 239051
rect 228671 239023 228699 239051
rect 228485 238961 228513 238989
rect 228547 238961 228575 238989
rect 228609 238961 228637 238989
rect 228671 238961 228699 238989
rect 228485 230147 228513 230175
rect 228547 230147 228575 230175
rect 228609 230147 228637 230175
rect 228671 230147 228699 230175
rect 228485 230085 228513 230113
rect 228547 230085 228575 230113
rect 228609 230085 228637 230113
rect 228671 230085 228699 230113
rect 228485 230023 228513 230051
rect 228547 230023 228575 230051
rect 228609 230023 228637 230051
rect 228671 230023 228699 230051
rect 228485 229961 228513 229989
rect 228547 229961 228575 229989
rect 228609 229961 228637 229989
rect 228671 229961 228699 229989
rect 228485 221147 228513 221175
rect 228547 221147 228575 221175
rect 228609 221147 228637 221175
rect 228671 221147 228699 221175
rect 228485 221085 228513 221113
rect 228547 221085 228575 221113
rect 228609 221085 228637 221113
rect 228671 221085 228699 221113
rect 228485 221023 228513 221051
rect 228547 221023 228575 221051
rect 228609 221023 228637 221051
rect 228671 221023 228699 221051
rect 228485 220961 228513 220989
rect 228547 220961 228575 220989
rect 228609 220961 228637 220989
rect 228671 220961 228699 220989
rect 228485 212147 228513 212175
rect 228547 212147 228575 212175
rect 228609 212147 228637 212175
rect 228671 212147 228699 212175
rect 228485 212085 228513 212113
rect 228547 212085 228575 212113
rect 228609 212085 228637 212113
rect 228671 212085 228699 212113
rect 228485 212023 228513 212051
rect 228547 212023 228575 212051
rect 228609 212023 228637 212051
rect 228671 212023 228699 212051
rect 228485 211961 228513 211989
rect 228547 211961 228575 211989
rect 228609 211961 228637 211989
rect 228671 211961 228699 211989
rect 228485 203147 228513 203175
rect 228547 203147 228575 203175
rect 228609 203147 228637 203175
rect 228671 203147 228699 203175
rect 228485 203085 228513 203113
rect 228547 203085 228575 203113
rect 228609 203085 228637 203113
rect 228671 203085 228699 203113
rect 228485 203023 228513 203051
rect 228547 203023 228575 203051
rect 228609 203023 228637 203051
rect 228671 203023 228699 203051
rect 228485 202961 228513 202989
rect 228547 202961 228575 202989
rect 228609 202961 228637 202989
rect 228671 202961 228699 202989
rect 228485 194147 228513 194175
rect 228547 194147 228575 194175
rect 228609 194147 228637 194175
rect 228671 194147 228699 194175
rect 228485 194085 228513 194113
rect 228547 194085 228575 194113
rect 228609 194085 228637 194113
rect 228671 194085 228699 194113
rect 228485 194023 228513 194051
rect 228547 194023 228575 194051
rect 228609 194023 228637 194051
rect 228671 194023 228699 194051
rect 228485 193961 228513 193989
rect 228547 193961 228575 193989
rect 228609 193961 228637 193989
rect 228671 193961 228699 193989
rect 228485 185147 228513 185175
rect 228547 185147 228575 185175
rect 228609 185147 228637 185175
rect 228671 185147 228699 185175
rect 228485 185085 228513 185113
rect 228547 185085 228575 185113
rect 228609 185085 228637 185113
rect 228671 185085 228699 185113
rect 228485 185023 228513 185051
rect 228547 185023 228575 185051
rect 228609 185023 228637 185051
rect 228671 185023 228699 185051
rect 228485 184961 228513 184989
rect 228547 184961 228575 184989
rect 228609 184961 228637 184989
rect 228671 184961 228699 184989
rect 228485 176147 228513 176175
rect 228547 176147 228575 176175
rect 228609 176147 228637 176175
rect 228671 176147 228699 176175
rect 228485 176085 228513 176113
rect 228547 176085 228575 176113
rect 228609 176085 228637 176113
rect 228671 176085 228699 176113
rect 228485 176023 228513 176051
rect 228547 176023 228575 176051
rect 228609 176023 228637 176051
rect 228671 176023 228699 176051
rect 228485 175961 228513 175989
rect 228547 175961 228575 175989
rect 228609 175961 228637 175989
rect 228671 175961 228699 175989
rect 228485 167147 228513 167175
rect 228547 167147 228575 167175
rect 228609 167147 228637 167175
rect 228671 167147 228699 167175
rect 228485 167085 228513 167113
rect 228547 167085 228575 167113
rect 228609 167085 228637 167113
rect 228671 167085 228699 167113
rect 228485 167023 228513 167051
rect 228547 167023 228575 167051
rect 228609 167023 228637 167051
rect 228671 167023 228699 167051
rect 228485 166961 228513 166989
rect 228547 166961 228575 166989
rect 228609 166961 228637 166989
rect 228671 166961 228699 166989
rect 228485 158147 228513 158175
rect 228547 158147 228575 158175
rect 228609 158147 228637 158175
rect 228671 158147 228699 158175
rect 228485 158085 228513 158113
rect 228547 158085 228575 158113
rect 228609 158085 228637 158113
rect 228671 158085 228699 158113
rect 228485 158023 228513 158051
rect 228547 158023 228575 158051
rect 228609 158023 228637 158051
rect 228671 158023 228699 158051
rect 228485 157961 228513 157989
rect 228547 157961 228575 157989
rect 228609 157961 228637 157989
rect 228671 157961 228699 157989
rect 228485 149147 228513 149175
rect 228547 149147 228575 149175
rect 228609 149147 228637 149175
rect 228671 149147 228699 149175
rect 228485 149085 228513 149113
rect 228547 149085 228575 149113
rect 228609 149085 228637 149113
rect 228671 149085 228699 149113
rect 228485 149023 228513 149051
rect 228547 149023 228575 149051
rect 228609 149023 228637 149051
rect 228671 149023 228699 149051
rect 228485 148961 228513 148989
rect 228547 148961 228575 148989
rect 228609 148961 228637 148989
rect 228671 148961 228699 148989
rect 228485 140147 228513 140175
rect 228547 140147 228575 140175
rect 228609 140147 228637 140175
rect 228671 140147 228699 140175
rect 228485 140085 228513 140113
rect 228547 140085 228575 140113
rect 228609 140085 228637 140113
rect 228671 140085 228699 140113
rect 228485 140023 228513 140051
rect 228547 140023 228575 140051
rect 228609 140023 228637 140051
rect 228671 140023 228699 140051
rect 228485 139961 228513 139989
rect 228547 139961 228575 139989
rect 228609 139961 228637 139989
rect 228671 139961 228699 139989
rect 228485 131147 228513 131175
rect 228547 131147 228575 131175
rect 228609 131147 228637 131175
rect 228671 131147 228699 131175
rect 228485 131085 228513 131113
rect 228547 131085 228575 131113
rect 228609 131085 228637 131113
rect 228671 131085 228699 131113
rect 228485 131023 228513 131051
rect 228547 131023 228575 131051
rect 228609 131023 228637 131051
rect 228671 131023 228699 131051
rect 228485 130961 228513 130989
rect 228547 130961 228575 130989
rect 228609 130961 228637 130989
rect 228671 130961 228699 130989
rect 228485 122147 228513 122175
rect 228547 122147 228575 122175
rect 228609 122147 228637 122175
rect 228671 122147 228699 122175
rect 228485 122085 228513 122113
rect 228547 122085 228575 122113
rect 228609 122085 228637 122113
rect 228671 122085 228699 122113
rect 228485 122023 228513 122051
rect 228547 122023 228575 122051
rect 228609 122023 228637 122051
rect 228671 122023 228699 122051
rect 228485 121961 228513 121989
rect 228547 121961 228575 121989
rect 228609 121961 228637 121989
rect 228671 121961 228699 121989
rect 228485 113147 228513 113175
rect 228547 113147 228575 113175
rect 228609 113147 228637 113175
rect 228671 113147 228699 113175
rect 228485 113085 228513 113113
rect 228547 113085 228575 113113
rect 228609 113085 228637 113113
rect 228671 113085 228699 113113
rect 228485 113023 228513 113051
rect 228547 113023 228575 113051
rect 228609 113023 228637 113051
rect 228671 113023 228699 113051
rect 228485 112961 228513 112989
rect 228547 112961 228575 112989
rect 228609 112961 228637 112989
rect 228671 112961 228699 112989
rect 228485 104147 228513 104175
rect 228547 104147 228575 104175
rect 228609 104147 228637 104175
rect 228671 104147 228699 104175
rect 228485 104085 228513 104113
rect 228547 104085 228575 104113
rect 228609 104085 228637 104113
rect 228671 104085 228699 104113
rect 228485 104023 228513 104051
rect 228547 104023 228575 104051
rect 228609 104023 228637 104051
rect 228671 104023 228699 104051
rect 228485 103961 228513 103989
rect 228547 103961 228575 103989
rect 228609 103961 228637 103989
rect 228671 103961 228699 103989
rect 228485 95147 228513 95175
rect 228547 95147 228575 95175
rect 228609 95147 228637 95175
rect 228671 95147 228699 95175
rect 228485 95085 228513 95113
rect 228547 95085 228575 95113
rect 228609 95085 228637 95113
rect 228671 95085 228699 95113
rect 228485 95023 228513 95051
rect 228547 95023 228575 95051
rect 228609 95023 228637 95051
rect 228671 95023 228699 95051
rect 228485 94961 228513 94989
rect 228547 94961 228575 94989
rect 228609 94961 228637 94989
rect 228671 94961 228699 94989
rect 228485 86147 228513 86175
rect 228547 86147 228575 86175
rect 228609 86147 228637 86175
rect 228671 86147 228699 86175
rect 228485 86085 228513 86113
rect 228547 86085 228575 86113
rect 228609 86085 228637 86113
rect 228671 86085 228699 86113
rect 228485 86023 228513 86051
rect 228547 86023 228575 86051
rect 228609 86023 228637 86051
rect 228671 86023 228699 86051
rect 228485 85961 228513 85989
rect 228547 85961 228575 85989
rect 228609 85961 228637 85989
rect 228671 85961 228699 85989
rect 228485 77147 228513 77175
rect 228547 77147 228575 77175
rect 228609 77147 228637 77175
rect 228671 77147 228699 77175
rect 228485 77085 228513 77113
rect 228547 77085 228575 77113
rect 228609 77085 228637 77113
rect 228671 77085 228699 77113
rect 228485 77023 228513 77051
rect 228547 77023 228575 77051
rect 228609 77023 228637 77051
rect 228671 77023 228699 77051
rect 228485 76961 228513 76989
rect 228547 76961 228575 76989
rect 228609 76961 228637 76989
rect 228671 76961 228699 76989
rect 228485 68147 228513 68175
rect 228547 68147 228575 68175
rect 228609 68147 228637 68175
rect 228671 68147 228699 68175
rect 228485 68085 228513 68113
rect 228547 68085 228575 68113
rect 228609 68085 228637 68113
rect 228671 68085 228699 68113
rect 228485 68023 228513 68051
rect 228547 68023 228575 68051
rect 228609 68023 228637 68051
rect 228671 68023 228699 68051
rect 228485 67961 228513 67989
rect 228547 67961 228575 67989
rect 228609 67961 228637 67989
rect 228671 67961 228699 67989
rect 228485 59147 228513 59175
rect 228547 59147 228575 59175
rect 228609 59147 228637 59175
rect 228671 59147 228699 59175
rect 228485 59085 228513 59113
rect 228547 59085 228575 59113
rect 228609 59085 228637 59113
rect 228671 59085 228699 59113
rect 228485 59023 228513 59051
rect 228547 59023 228575 59051
rect 228609 59023 228637 59051
rect 228671 59023 228699 59051
rect 228485 58961 228513 58989
rect 228547 58961 228575 58989
rect 228609 58961 228637 58989
rect 228671 58961 228699 58989
rect 228485 50147 228513 50175
rect 228547 50147 228575 50175
rect 228609 50147 228637 50175
rect 228671 50147 228699 50175
rect 228485 50085 228513 50113
rect 228547 50085 228575 50113
rect 228609 50085 228637 50113
rect 228671 50085 228699 50113
rect 228485 50023 228513 50051
rect 228547 50023 228575 50051
rect 228609 50023 228637 50051
rect 228671 50023 228699 50051
rect 228485 49961 228513 49989
rect 228547 49961 228575 49989
rect 228609 49961 228637 49989
rect 228671 49961 228699 49989
rect 228485 41147 228513 41175
rect 228547 41147 228575 41175
rect 228609 41147 228637 41175
rect 228671 41147 228699 41175
rect 228485 41085 228513 41113
rect 228547 41085 228575 41113
rect 228609 41085 228637 41113
rect 228671 41085 228699 41113
rect 228485 41023 228513 41051
rect 228547 41023 228575 41051
rect 228609 41023 228637 41051
rect 228671 41023 228699 41051
rect 228485 40961 228513 40989
rect 228547 40961 228575 40989
rect 228609 40961 228637 40989
rect 228671 40961 228699 40989
rect 228485 32147 228513 32175
rect 228547 32147 228575 32175
rect 228609 32147 228637 32175
rect 228671 32147 228699 32175
rect 228485 32085 228513 32113
rect 228547 32085 228575 32113
rect 228609 32085 228637 32113
rect 228671 32085 228699 32113
rect 228485 32023 228513 32051
rect 228547 32023 228575 32051
rect 228609 32023 228637 32051
rect 228671 32023 228699 32051
rect 228485 31961 228513 31989
rect 228547 31961 228575 31989
rect 228609 31961 228637 31989
rect 228671 31961 228699 31989
rect 228485 23147 228513 23175
rect 228547 23147 228575 23175
rect 228609 23147 228637 23175
rect 228671 23147 228699 23175
rect 228485 23085 228513 23113
rect 228547 23085 228575 23113
rect 228609 23085 228637 23113
rect 228671 23085 228699 23113
rect 228485 23023 228513 23051
rect 228547 23023 228575 23051
rect 228609 23023 228637 23051
rect 228671 23023 228699 23051
rect 228485 22961 228513 22989
rect 228547 22961 228575 22989
rect 228609 22961 228637 22989
rect 228671 22961 228699 22989
rect 228485 14147 228513 14175
rect 228547 14147 228575 14175
rect 228609 14147 228637 14175
rect 228671 14147 228699 14175
rect 228485 14085 228513 14113
rect 228547 14085 228575 14113
rect 228609 14085 228637 14113
rect 228671 14085 228699 14113
rect 228485 14023 228513 14051
rect 228547 14023 228575 14051
rect 228609 14023 228637 14051
rect 228671 14023 228699 14051
rect 228485 13961 228513 13989
rect 228547 13961 228575 13989
rect 228609 13961 228637 13989
rect 228671 13961 228699 13989
rect 228485 5147 228513 5175
rect 228547 5147 228575 5175
rect 228609 5147 228637 5175
rect 228671 5147 228699 5175
rect 228485 5085 228513 5113
rect 228547 5085 228575 5113
rect 228609 5085 228637 5113
rect 228671 5085 228699 5113
rect 228485 5023 228513 5051
rect 228547 5023 228575 5051
rect 228609 5023 228637 5051
rect 228671 5023 228699 5051
rect 228485 4961 228513 4989
rect 228547 4961 228575 4989
rect 228609 4961 228637 4989
rect 228671 4961 228699 4989
rect 228485 -588 228513 -560
rect 228547 -588 228575 -560
rect 228609 -588 228637 -560
rect 228671 -588 228699 -560
rect 228485 -650 228513 -622
rect 228547 -650 228575 -622
rect 228609 -650 228637 -622
rect 228671 -650 228699 -622
rect 228485 -712 228513 -684
rect 228547 -712 228575 -684
rect 228609 -712 228637 -684
rect 228671 -712 228699 -684
rect 228485 -774 228513 -746
rect 228547 -774 228575 -746
rect 228609 -774 228637 -746
rect 228671 -774 228699 -746
rect 235625 298578 235653 298606
rect 235687 298578 235715 298606
rect 235749 298578 235777 298606
rect 235811 298578 235839 298606
rect 235625 298516 235653 298544
rect 235687 298516 235715 298544
rect 235749 298516 235777 298544
rect 235811 298516 235839 298544
rect 235625 298454 235653 298482
rect 235687 298454 235715 298482
rect 235749 298454 235777 298482
rect 235811 298454 235839 298482
rect 235625 298392 235653 298420
rect 235687 298392 235715 298420
rect 235749 298392 235777 298420
rect 235811 298392 235839 298420
rect 235625 290147 235653 290175
rect 235687 290147 235715 290175
rect 235749 290147 235777 290175
rect 235811 290147 235839 290175
rect 235625 290085 235653 290113
rect 235687 290085 235715 290113
rect 235749 290085 235777 290113
rect 235811 290085 235839 290113
rect 235625 290023 235653 290051
rect 235687 290023 235715 290051
rect 235749 290023 235777 290051
rect 235811 290023 235839 290051
rect 235625 289961 235653 289989
rect 235687 289961 235715 289989
rect 235749 289961 235777 289989
rect 235811 289961 235839 289989
rect 235625 281147 235653 281175
rect 235687 281147 235715 281175
rect 235749 281147 235777 281175
rect 235811 281147 235839 281175
rect 235625 281085 235653 281113
rect 235687 281085 235715 281113
rect 235749 281085 235777 281113
rect 235811 281085 235839 281113
rect 235625 281023 235653 281051
rect 235687 281023 235715 281051
rect 235749 281023 235777 281051
rect 235811 281023 235839 281051
rect 235625 280961 235653 280989
rect 235687 280961 235715 280989
rect 235749 280961 235777 280989
rect 235811 280961 235839 280989
rect 235625 272147 235653 272175
rect 235687 272147 235715 272175
rect 235749 272147 235777 272175
rect 235811 272147 235839 272175
rect 235625 272085 235653 272113
rect 235687 272085 235715 272113
rect 235749 272085 235777 272113
rect 235811 272085 235839 272113
rect 235625 272023 235653 272051
rect 235687 272023 235715 272051
rect 235749 272023 235777 272051
rect 235811 272023 235839 272051
rect 235625 271961 235653 271989
rect 235687 271961 235715 271989
rect 235749 271961 235777 271989
rect 235811 271961 235839 271989
rect 235625 263147 235653 263175
rect 235687 263147 235715 263175
rect 235749 263147 235777 263175
rect 235811 263147 235839 263175
rect 235625 263085 235653 263113
rect 235687 263085 235715 263113
rect 235749 263085 235777 263113
rect 235811 263085 235839 263113
rect 235625 263023 235653 263051
rect 235687 263023 235715 263051
rect 235749 263023 235777 263051
rect 235811 263023 235839 263051
rect 235625 262961 235653 262989
rect 235687 262961 235715 262989
rect 235749 262961 235777 262989
rect 235811 262961 235839 262989
rect 235625 254147 235653 254175
rect 235687 254147 235715 254175
rect 235749 254147 235777 254175
rect 235811 254147 235839 254175
rect 235625 254085 235653 254113
rect 235687 254085 235715 254113
rect 235749 254085 235777 254113
rect 235811 254085 235839 254113
rect 235625 254023 235653 254051
rect 235687 254023 235715 254051
rect 235749 254023 235777 254051
rect 235811 254023 235839 254051
rect 235625 253961 235653 253989
rect 235687 253961 235715 253989
rect 235749 253961 235777 253989
rect 235811 253961 235839 253989
rect 235625 245147 235653 245175
rect 235687 245147 235715 245175
rect 235749 245147 235777 245175
rect 235811 245147 235839 245175
rect 235625 245085 235653 245113
rect 235687 245085 235715 245113
rect 235749 245085 235777 245113
rect 235811 245085 235839 245113
rect 235625 245023 235653 245051
rect 235687 245023 235715 245051
rect 235749 245023 235777 245051
rect 235811 245023 235839 245051
rect 235625 244961 235653 244989
rect 235687 244961 235715 244989
rect 235749 244961 235777 244989
rect 235811 244961 235839 244989
rect 235625 236147 235653 236175
rect 235687 236147 235715 236175
rect 235749 236147 235777 236175
rect 235811 236147 235839 236175
rect 235625 236085 235653 236113
rect 235687 236085 235715 236113
rect 235749 236085 235777 236113
rect 235811 236085 235839 236113
rect 235625 236023 235653 236051
rect 235687 236023 235715 236051
rect 235749 236023 235777 236051
rect 235811 236023 235839 236051
rect 235625 235961 235653 235989
rect 235687 235961 235715 235989
rect 235749 235961 235777 235989
rect 235811 235961 235839 235989
rect 235625 227147 235653 227175
rect 235687 227147 235715 227175
rect 235749 227147 235777 227175
rect 235811 227147 235839 227175
rect 235625 227085 235653 227113
rect 235687 227085 235715 227113
rect 235749 227085 235777 227113
rect 235811 227085 235839 227113
rect 235625 227023 235653 227051
rect 235687 227023 235715 227051
rect 235749 227023 235777 227051
rect 235811 227023 235839 227051
rect 235625 226961 235653 226989
rect 235687 226961 235715 226989
rect 235749 226961 235777 226989
rect 235811 226961 235839 226989
rect 235625 218147 235653 218175
rect 235687 218147 235715 218175
rect 235749 218147 235777 218175
rect 235811 218147 235839 218175
rect 235625 218085 235653 218113
rect 235687 218085 235715 218113
rect 235749 218085 235777 218113
rect 235811 218085 235839 218113
rect 235625 218023 235653 218051
rect 235687 218023 235715 218051
rect 235749 218023 235777 218051
rect 235811 218023 235839 218051
rect 235625 217961 235653 217989
rect 235687 217961 235715 217989
rect 235749 217961 235777 217989
rect 235811 217961 235839 217989
rect 235625 209147 235653 209175
rect 235687 209147 235715 209175
rect 235749 209147 235777 209175
rect 235811 209147 235839 209175
rect 235625 209085 235653 209113
rect 235687 209085 235715 209113
rect 235749 209085 235777 209113
rect 235811 209085 235839 209113
rect 235625 209023 235653 209051
rect 235687 209023 235715 209051
rect 235749 209023 235777 209051
rect 235811 209023 235839 209051
rect 235625 208961 235653 208989
rect 235687 208961 235715 208989
rect 235749 208961 235777 208989
rect 235811 208961 235839 208989
rect 235625 200147 235653 200175
rect 235687 200147 235715 200175
rect 235749 200147 235777 200175
rect 235811 200147 235839 200175
rect 235625 200085 235653 200113
rect 235687 200085 235715 200113
rect 235749 200085 235777 200113
rect 235811 200085 235839 200113
rect 235625 200023 235653 200051
rect 235687 200023 235715 200051
rect 235749 200023 235777 200051
rect 235811 200023 235839 200051
rect 235625 199961 235653 199989
rect 235687 199961 235715 199989
rect 235749 199961 235777 199989
rect 235811 199961 235839 199989
rect 235625 191147 235653 191175
rect 235687 191147 235715 191175
rect 235749 191147 235777 191175
rect 235811 191147 235839 191175
rect 235625 191085 235653 191113
rect 235687 191085 235715 191113
rect 235749 191085 235777 191113
rect 235811 191085 235839 191113
rect 235625 191023 235653 191051
rect 235687 191023 235715 191051
rect 235749 191023 235777 191051
rect 235811 191023 235839 191051
rect 235625 190961 235653 190989
rect 235687 190961 235715 190989
rect 235749 190961 235777 190989
rect 235811 190961 235839 190989
rect 235625 182147 235653 182175
rect 235687 182147 235715 182175
rect 235749 182147 235777 182175
rect 235811 182147 235839 182175
rect 235625 182085 235653 182113
rect 235687 182085 235715 182113
rect 235749 182085 235777 182113
rect 235811 182085 235839 182113
rect 235625 182023 235653 182051
rect 235687 182023 235715 182051
rect 235749 182023 235777 182051
rect 235811 182023 235839 182051
rect 235625 181961 235653 181989
rect 235687 181961 235715 181989
rect 235749 181961 235777 181989
rect 235811 181961 235839 181989
rect 235625 173147 235653 173175
rect 235687 173147 235715 173175
rect 235749 173147 235777 173175
rect 235811 173147 235839 173175
rect 235625 173085 235653 173113
rect 235687 173085 235715 173113
rect 235749 173085 235777 173113
rect 235811 173085 235839 173113
rect 235625 173023 235653 173051
rect 235687 173023 235715 173051
rect 235749 173023 235777 173051
rect 235811 173023 235839 173051
rect 235625 172961 235653 172989
rect 235687 172961 235715 172989
rect 235749 172961 235777 172989
rect 235811 172961 235839 172989
rect 235625 164147 235653 164175
rect 235687 164147 235715 164175
rect 235749 164147 235777 164175
rect 235811 164147 235839 164175
rect 235625 164085 235653 164113
rect 235687 164085 235715 164113
rect 235749 164085 235777 164113
rect 235811 164085 235839 164113
rect 235625 164023 235653 164051
rect 235687 164023 235715 164051
rect 235749 164023 235777 164051
rect 235811 164023 235839 164051
rect 235625 163961 235653 163989
rect 235687 163961 235715 163989
rect 235749 163961 235777 163989
rect 235811 163961 235839 163989
rect 235625 155147 235653 155175
rect 235687 155147 235715 155175
rect 235749 155147 235777 155175
rect 235811 155147 235839 155175
rect 235625 155085 235653 155113
rect 235687 155085 235715 155113
rect 235749 155085 235777 155113
rect 235811 155085 235839 155113
rect 235625 155023 235653 155051
rect 235687 155023 235715 155051
rect 235749 155023 235777 155051
rect 235811 155023 235839 155051
rect 235625 154961 235653 154989
rect 235687 154961 235715 154989
rect 235749 154961 235777 154989
rect 235811 154961 235839 154989
rect 235625 146147 235653 146175
rect 235687 146147 235715 146175
rect 235749 146147 235777 146175
rect 235811 146147 235839 146175
rect 235625 146085 235653 146113
rect 235687 146085 235715 146113
rect 235749 146085 235777 146113
rect 235811 146085 235839 146113
rect 235625 146023 235653 146051
rect 235687 146023 235715 146051
rect 235749 146023 235777 146051
rect 235811 146023 235839 146051
rect 235625 145961 235653 145989
rect 235687 145961 235715 145989
rect 235749 145961 235777 145989
rect 235811 145961 235839 145989
rect 235625 137147 235653 137175
rect 235687 137147 235715 137175
rect 235749 137147 235777 137175
rect 235811 137147 235839 137175
rect 235625 137085 235653 137113
rect 235687 137085 235715 137113
rect 235749 137085 235777 137113
rect 235811 137085 235839 137113
rect 235625 137023 235653 137051
rect 235687 137023 235715 137051
rect 235749 137023 235777 137051
rect 235811 137023 235839 137051
rect 235625 136961 235653 136989
rect 235687 136961 235715 136989
rect 235749 136961 235777 136989
rect 235811 136961 235839 136989
rect 235625 128147 235653 128175
rect 235687 128147 235715 128175
rect 235749 128147 235777 128175
rect 235811 128147 235839 128175
rect 235625 128085 235653 128113
rect 235687 128085 235715 128113
rect 235749 128085 235777 128113
rect 235811 128085 235839 128113
rect 235625 128023 235653 128051
rect 235687 128023 235715 128051
rect 235749 128023 235777 128051
rect 235811 128023 235839 128051
rect 235625 127961 235653 127989
rect 235687 127961 235715 127989
rect 235749 127961 235777 127989
rect 235811 127961 235839 127989
rect 235625 119147 235653 119175
rect 235687 119147 235715 119175
rect 235749 119147 235777 119175
rect 235811 119147 235839 119175
rect 235625 119085 235653 119113
rect 235687 119085 235715 119113
rect 235749 119085 235777 119113
rect 235811 119085 235839 119113
rect 235625 119023 235653 119051
rect 235687 119023 235715 119051
rect 235749 119023 235777 119051
rect 235811 119023 235839 119051
rect 235625 118961 235653 118989
rect 235687 118961 235715 118989
rect 235749 118961 235777 118989
rect 235811 118961 235839 118989
rect 235625 110147 235653 110175
rect 235687 110147 235715 110175
rect 235749 110147 235777 110175
rect 235811 110147 235839 110175
rect 235625 110085 235653 110113
rect 235687 110085 235715 110113
rect 235749 110085 235777 110113
rect 235811 110085 235839 110113
rect 235625 110023 235653 110051
rect 235687 110023 235715 110051
rect 235749 110023 235777 110051
rect 235811 110023 235839 110051
rect 235625 109961 235653 109989
rect 235687 109961 235715 109989
rect 235749 109961 235777 109989
rect 235811 109961 235839 109989
rect 235625 101147 235653 101175
rect 235687 101147 235715 101175
rect 235749 101147 235777 101175
rect 235811 101147 235839 101175
rect 235625 101085 235653 101113
rect 235687 101085 235715 101113
rect 235749 101085 235777 101113
rect 235811 101085 235839 101113
rect 235625 101023 235653 101051
rect 235687 101023 235715 101051
rect 235749 101023 235777 101051
rect 235811 101023 235839 101051
rect 235625 100961 235653 100989
rect 235687 100961 235715 100989
rect 235749 100961 235777 100989
rect 235811 100961 235839 100989
rect 235625 92147 235653 92175
rect 235687 92147 235715 92175
rect 235749 92147 235777 92175
rect 235811 92147 235839 92175
rect 235625 92085 235653 92113
rect 235687 92085 235715 92113
rect 235749 92085 235777 92113
rect 235811 92085 235839 92113
rect 235625 92023 235653 92051
rect 235687 92023 235715 92051
rect 235749 92023 235777 92051
rect 235811 92023 235839 92051
rect 235625 91961 235653 91989
rect 235687 91961 235715 91989
rect 235749 91961 235777 91989
rect 235811 91961 235839 91989
rect 235625 83147 235653 83175
rect 235687 83147 235715 83175
rect 235749 83147 235777 83175
rect 235811 83147 235839 83175
rect 235625 83085 235653 83113
rect 235687 83085 235715 83113
rect 235749 83085 235777 83113
rect 235811 83085 235839 83113
rect 235625 83023 235653 83051
rect 235687 83023 235715 83051
rect 235749 83023 235777 83051
rect 235811 83023 235839 83051
rect 235625 82961 235653 82989
rect 235687 82961 235715 82989
rect 235749 82961 235777 82989
rect 235811 82961 235839 82989
rect 235625 74147 235653 74175
rect 235687 74147 235715 74175
rect 235749 74147 235777 74175
rect 235811 74147 235839 74175
rect 235625 74085 235653 74113
rect 235687 74085 235715 74113
rect 235749 74085 235777 74113
rect 235811 74085 235839 74113
rect 235625 74023 235653 74051
rect 235687 74023 235715 74051
rect 235749 74023 235777 74051
rect 235811 74023 235839 74051
rect 235625 73961 235653 73989
rect 235687 73961 235715 73989
rect 235749 73961 235777 73989
rect 235811 73961 235839 73989
rect 235625 65147 235653 65175
rect 235687 65147 235715 65175
rect 235749 65147 235777 65175
rect 235811 65147 235839 65175
rect 235625 65085 235653 65113
rect 235687 65085 235715 65113
rect 235749 65085 235777 65113
rect 235811 65085 235839 65113
rect 235625 65023 235653 65051
rect 235687 65023 235715 65051
rect 235749 65023 235777 65051
rect 235811 65023 235839 65051
rect 235625 64961 235653 64989
rect 235687 64961 235715 64989
rect 235749 64961 235777 64989
rect 235811 64961 235839 64989
rect 235625 56147 235653 56175
rect 235687 56147 235715 56175
rect 235749 56147 235777 56175
rect 235811 56147 235839 56175
rect 235625 56085 235653 56113
rect 235687 56085 235715 56113
rect 235749 56085 235777 56113
rect 235811 56085 235839 56113
rect 235625 56023 235653 56051
rect 235687 56023 235715 56051
rect 235749 56023 235777 56051
rect 235811 56023 235839 56051
rect 235625 55961 235653 55989
rect 235687 55961 235715 55989
rect 235749 55961 235777 55989
rect 235811 55961 235839 55989
rect 235625 47147 235653 47175
rect 235687 47147 235715 47175
rect 235749 47147 235777 47175
rect 235811 47147 235839 47175
rect 235625 47085 235653 47113
rect 235687 47085 235715 47113
rect 235749 47085 235777 47113
rect 235811 47085 235839 47113
rect 235625 47023 235653 47051
rect 235687 47023 235715 47051
rect 235749 47023 235777 47051
rect 235811 47023 235839 47051
rect 235625 46961 235653 46989
rect 235687 46961 235715 46989
rect 235749 46961 235777 46989
rect 235811 46961 235839 46989
rect 235625 38147 235653 38175
rect 235687 38147 235715 38175
rect 235749 38147 235777 38175
rect 235811 38147 235839 38175
rect 235625 38085 235653 38113
rect 235687 38085 235715 38113
rect 235749 38085 235777 38113
rect 235811 38085 235839 38113
rect 235625 38023 235653 38051
rect 235687 38023 235715 38051
rect 235749 38023 235777 38051
rect 235811 38023 235839 38051
rect 235625 37961 235653 37989
rect 235687 37961 235715 37989
rect 235749 37961 235777 37989
rect 235811 37961 235839 37989
rect 235625 29147 235653 29175
rect 235687 29147 235715 29175
rect 235749 29147 235777 29175
rect 235811 29147 235839 29175
rect 235625 29085 235653 29113
rect 235687 29085 235715 29113
rect 235749 29085 235777 29113
rect 235811 29085 235839 29113
rect 235625 29023 235653 29051
rect 235687 29023 235715 29051
rect 235749 29023 235777 29051
rect 235811 29023 235839 29051
rect 235625 28961 235653 28989
rect 235687 28961 235715 28989
rect 235749 28961 235777 28989
rect 235811 28961 235839 28989
rect 235625 20147 235653 20175
rect 235687 20147 235715 20175
rect 235749 20147 235777 20175
rect 235811 20147 235839 20175
rect 235625 20085 235653 20113
rect 235687 20085 235715 20113
rect 235749 20085 235777 20113
rect 235811 20085 235839 20113
rect 235625 20023 235653 20051
rect 235687 20023 235715 20051
rect 235749 20023 235777 20051
rect 235811 20023 235839 20051
rect 235625 19961 235653 19989
rect 235687 19961 235715 19989
rect 235749 19961 235777 19989
rect 235811 19961 235839 19989
rect 235625 11147 235653 11175
rect 235687 11147 235715 11175
rect 235749 11147 235777 11175
rect 235811 11147 235839 11175
rect 235625 11085 235653 11113
rect 235687 11085 235715 11113
rect 235749 11085 235777 11113
rect 235811 11085 235839 11113
rect 235625 11023 235653 11051
rect 235687 11023 235715 11051
rect 235749 11023 235777 11051
rect 235811 11023 235839 11051
rect 235625 10961 235653 10989
rect 235687 10961 235715 10989
rect 235749 10961 235777 10989
rect 235811 10961 235839 10989
rect 235625 2147 235653 2175
rect 235687 2147 235715 2175
rect 235749 2147 235777 2175
rect 235811 2147 235839 2175
rect 235625 2085 235653 2113
rect 235687 2085 235715 2113
rect 235749 2085 235777 2113
rect 235811 2085 235839 2113
rect 235625 2023 235653 2051
rect 235687 2023 235715 2051
rect 235749 2023 235777 2051
rect 235811 2023 235839 2051
rect 235625 1961 235653 1989
rect 235687 1961 235715 1989
rect 235749 1961 235777 1989
rect 235811 1961 235839 1989
rect 235625 -108 235653 -80
rect 235687 -108 235715 -80
rect 235749 -108 235777 -80
rect 235811 -108 235839 -80
rect 235625 -170 235653 -142
rect 235687 -170 235715 -142
rect 235749 -170 235777 -142
rect 235811 -170 235839 -142
rect 235625 -232 235653 -204
rect 235687 -232 235715 -204
rect 235749 -232 235777 -204
rect 235811 -232 235839 -204
rect 235625 -294 235653 -266
rect 235687 -294 235715 -266
rect 235749 -294 235777 -266
rect 235811 -294 235839 -266
rect 237485 299058 237513 299086
rect 237547 299058 237575 299086
rect 237609 299058 237637 299086
rect 237671 299058 237699 299086
rect 237485 298996 237513 299024
rect 237547 298996 237575 299024
rect 237609 298996 237637 299024
rect 237671 298996 237699 299024
rect 237485 298934 237513 298962
rect 237547 298934 237575 298962
rect 237609 298934 237637 298962
rect 237671 298934 237699 298962
rect 237485 298872 237513 298900
rect 237547 298872 237575 298900
rect 237609 298872 237637 298900
rect 237671 298872 237699 298900
rect 237485 293147 237513 293175
rect 237547 293147 237575 293175
rect 237609 293147 237637 293175
rect 237671 293147 237699 293175
rect 237485 293085 237513 293113
rect 237547 293085 237575 293113
rect 237609 293085 237637 293113
rect 237671 293085 237699 293113
rect 237485 293023 237513 293051
rect 237547 293023 237575 293051
rect 237609 293023 237637 293051
rect 237671 293023 237699 293051
rect 237485 292961 237513 292989
rect 237547 292961 237575 292989
rect 237609 292961 237637 292989
rect 237671 292961 237699 292989
rect 237485 284147 237513 284175
rect 237547 284147 237575 284175
rect 237609 284147 237637 284175
rect 237671 284147 237699 284175
rect 237485 284085 237513 284113
rect 237547 284085 237575 284113
rect 237609 284085 237637 284113
rect 237671 284085 237699 284113
rect 237485 284023 237513 284051
rect 237547 284023 237575 284051
rect 237609 284023 237637 284051
rect 237671 284023 237699 284051
rect 237485 283961 237513 283989
rect 237547 283961 237575 283989
rect 237609 283961 237637 283989
rect 237671 283961 237699 283989
rect 237485 275147 237513 275175
rect 237547 275147 237575 275175
rect 237609 275147 237637 275175
rect 237671 275147 237699 275175
rect 237485 275085 237513 275113
rect 237547 275085 237575 275113
rect 237609 275085 237637 275113
rect 237671 275085 237699 275113
rect 237485 275023 237513 275051
rect 237547 275023 237575 275051
rect 237609 275023 237637 275051
rect 237671 275023 237699 275051
rect 237485 274961 237513 274989
rect 237547 274961 237575 274989
rect 237609 274961 237637 274989
rect 237671 274961 237699 274989
rect 237485 266147 237513 266175
rect 237547 266147 237575 266175
rect 237609 266147 237637 266175
rect 237671 266147 237699 266175
rect 237485 266085 237513 266113
rect 237547 266085 237575 266113
rect 237609 266085 237637 266113
rect 237671 266085 237699 266113
rect 237485 266023 237513 266051
rect 237547 266023 237575 266051
rect 237609 266023 237637 266051
rect 237671 266023 237699 266051
rect 237485 265961 237513 265989
rect 237547 265961 237575 265989
rect 237609 265961 237637 265989
rect 237671 265961 237699 265989
rect 237485 257147 237513 257175
rect 237547 257147 237575 257175
rect 237609 257147 237637 257175
rect 237671 257147 237699 257175
rect 237485 257085 237513 257113
rect 237547 257085 237575 257113
rect 237609 257085 237637 257113
rect 237671 257085 237699 257113
rect 237485 257023 237513 257051
rect 237547 257023 237575 257051
rect 237609 257023 237637 257051
rect 237671 257023 237699 257051
rect 237485 256961 237513 256989
rect 237547 256961 237575 256989
rect 237609 256961 237637 256989
rect 237671 256961 237699 256989
rect 237485 248147 237513 248175
rect 237547 248147 237575 248175
rect 237609 248147 237637 248175
rect 237671 248147 237699 248175
rect 237485 248085 237513 248113
rect 237547 248085 237575 248113
rect 237609 248085 237637 248113
rect 237671 248085 237699 248113
rect 237485 248023 237513 248051
rect 237547 248023 237575 248051
rect 237609 248023 237637 248051
rect 237671 248023 237699 248051
rect 237485 247961 237513 247989
rect 237547 247961 237575 247989
rect 237609 247961 237637 247989
rect 237671 247961 237699 247989
rect 237485 239147 237513 239175
rect 237547 239147 237575 239175
rect 237609 239147 237637 239175
rect 237671 239147 237699 239175
rect 237485 239085 237513 239113
rect 237547 239085 237575 239113
rect 237609 239085 237637 239113
rect 237671 239085 237699 239113
rect 237485 239023 237513 239051
rect 237547 239023 237575 239051
rect 237609 239023 237637 239051
rect 237671 239023 237699 239051
rect 237485 238961 237513 238989
rect 237547 238961 237575 238989
rect 237609 238961 237637 238989
rect 237671 238961 237699 238989
rect 237485 230147 237513 230175
rect 237547 230147 237575 230175
rect 237609 230147 237637 230175
rect 237671 230147 237699 230175
rect 237485 230085 237513 230113
rect 237547 230085 237575 230113
rect 237609 230085 237637 230113
rect 237671 230085 237699 230113
rect 237485 230023 237513 230051
rect 237547 230023 237575 230051
rect 237609 230023 237637 230051
rect 237671 230023 237699 230051
rect 237485 229961 237513 229989
rect 237547 229961 237575 229989
rect 237609 229961 237637 229989
rect 237671 229961 237699 229989
rect 237485 221147 237513 221175
rect 237547 221147 237575 221175
rect 237609 221147 237637 221175
rect 237671 221147 237699 221175
rect 237485 221085 237513 221113
rect 237547 221085 237575 221113
rect 237609 221085 237637 221113
rect 237671 221085 237699 221113
rect 237485 221023 237513 221051
rect 237547 221023 237575 221051
rect 237609 221023 237637 221051
rect 237671 221023 237699 221051
rect 237485 220961 237513 220989
rect 237547 220961 237575 220989
rect 237609 220961 237637 220989
rect 237671 220961 237699 220989
rect 237485 212147 237513 212175
rect 237547 212147 237575 212175
rect 237609 212147 237637 212175
rect 237671 212147 237699 212175
rect 237485 212085 237513 212113
rect 237547 212085 237575 212113
rect 237609 212085 237637 212113
rect 237671 212085 237699 212113
rect 237485 212023 237513 212051
rect 237547 212023 237575 212051
rect 237609 212023 237637 212051
rect 237671 212023 237699 212051
rect 237485 211961 237513 211989
rect 237547 211961 237575 211989
rect 237609 211961 237637 211989
rect 237671 211961 237699 211989
rect 237485 203147 237513 203175
rect 237547 203147 237575 203175
rect 237609 203147 237637 203175
rect 237671 203147 237699 203175
rect 237485 203085 237513 203113
rect 237547 203085 237575 203113
rect 237609 203085 237637 203113
rect 237671 203085 237699 203113
rect 237485 203023 237513 203051
rect 237547 203023 237575 203051
rect 237609 203023 237637 203051
rect 237671 203023 237699 203051
rect 237485 202961 237513 202989
rect 237547 202961 237575 202989
rect 237609 202961 237637 202989
rect 237671 202961 237699 202989
rect 237485 194147 237513 194175
rect 237547 194147 237575 194175
rect 237609 194147 237637 194175
rect 237671 194147 237699 194175
rect 237485 194085 237513 194113
rect 237547 194085 237575 194113
rect 237609 194085 237637 194113
rect 237671 194085 237699 194113
rect 237485 194023 237513 194051
rect 237547 194023 237575 194051
rect 237609 194023 237637 194051
rect 237671 194023 237699 194051
rect 237485 193961 237513 193989
rect 237547 193961 237575 193989
rect 237609 193961 237637 193989
rect 237671 193961 237699 193989
rect 237485 185147 237513 185175
rect 237547 185147 237575 185175
rect 237609 185147 237637 185175
rect 237671 185147 237699 185175
rect 237485 185085 237513 185113
rect 237547 185085 237575 185113
rect 237609 185085 237637 185113
rect 237671 185085 237699 185113
rect 237485 185023 237513 185051
rect 237547 185023 237575 185051
rect 237609 185023 237637 185051
rect 237671 185023 237699 185051
rect 237485 184961 237513 184989
rect 237547 184961 237575 184989
rect 237609 184961 237637 184989
rect 237671 184961 237699 184989
rect 237485 176147 237513 176175
rect 237547 176147 237575 176175
rect 237609 176147 237637 176175
rect 237671 176147 237699 176175
rect 237485 176085 237513 176113
rect 237547 176085 237575 176113
rect 237609 176085 237637 176113
rect 237671 176085 237699 176113
rect 237485 176023 237513 176051
rect 237547 176023 237575 176051
rect 237609 176023 237637 176051
rect 237671 176023 237699 176051
rect 237485 175961 237513 175989
rect 237547 175961 237575 175989
rect 237609 175961 237637 175989
rect 237671 175961 237699 175989
rect 237485 167147 237513 167175
rect 237547 167147 237575 167175
rect 237609 167147 237637 167175
rect 237671 167147 237699 167175
rect 237485 167085 237513 167113
rect 237547 167085 237575 167113
rect 237609 167085 237637 167113
rect 237671 167085 237699 167113
rect 237485 167023 237513 167051
rect 237547 167023 237575 167051
rect 237609 167023 237637 167051
rect 237671 167023 237699 167051
rect 237485 166961 237513 166989
rect 237547 166961 237575 166989
rect 237609 166961 237637 166989
rect 237671 166961 237699 166989
rect 237485 158147 237513 158175
rect 237547 158147 237575 158175
rect 237609 158147 237637 158175
rect 237671 158147 237699 158175
rect 237485 158085 237513 158113
rect 237547 158085 237575 158113
rect 237609 158085 237637 158113
rect 237671 158085 237699 158113
rect 237485 158023 237513 158051
rect 237547 158023 237575 158051
rect 237609 158023 237637 158051
rect 237671 158023 237699 158051
rect 237485 157961 237513 157989
rect 237547 157961 237575 157989
rect 237609 157961 237637 157989
rect 237671 157961 237699 157989
rect 237485 149147 237513 149175
rect 237547 149147 237575 149175
rect 237609 149147 237637 149175
rect 237671 149147 237699 149175
rect 237485 149085 237513 149113
rect 237547 149085 237575 149113
rect 237609 149085 237637 149113
rect 237671 149085 237699 149113
rect 237485 149023 237513 149051
rect 237547 149023 237575 149051
rect 237609 149023 237637 149051
rect 237671 149023 237699 149051
rect 237485 148961 237513 148989
rect 237547 148961 237575 148989
rect 237609 148961 237637 148989
rect 237671 148961 237699 148989
rect 237485 140147 237513 140175
rect 237547 140147 237575 140175
rect 237609 140147 237637 140175
rect 237671 140147 237699 140175
rect 237485 140085 237513 140113
rect 237547 140085 237575 140113
rect 237609 140085 237637 140113
rect 237671 140085 237699 140113
rect 237485 140023 237513 140051
rect 237547 140023 237575 140051
rect 237609 140023 237637 140051
rect 237671 140023 237699 140051
rect 237485 139961 237513 139989
rect 237547 139961 237575 139989
rect 237609 139961 237637 139989
rect 237671 139961 237699 139989
rect 237485 131147 237513 131175
rect 237547 131147 237575 131175
rect 237609 131147 237637 131175
rect 237671 131147 237699 131175
rect 237485 131085 237513 131113
rect 237547 131085 237575 131113
rect 237609 131085 237637 131113
rect 237671 131085 237699 131113
rect 237485 131023 237513 131051
rect 237547 131023 237575 131051
rect 237609 131023 237637 131051
rect 237671 131023 237699 131051
rect 237485 130961 237513 130989
rect 237547 130961 237575 130989
rect 237609 130961 237637 130989
rect 237671 130961 237699 130989
rect 237485 122147 237513 122175
rect 237547 122147 237575 122175
rect 237609 122147 237637 122175
rect 237671 122147 237699 122175
rect 237485 122085 237513 122113
rect 237547 122085 237575 122113
rect 237609 122085 237637 122113
rect 237671 122085 237699 122113
rect 237485 122023 237513 122051
rect 237547 122023 237575 122051
rect 237609 122023 237637 122051
rect 237671 122023 237699 122051
rect 237485 121961 237513 121989
rect 237547 121961 237575 121989
rect 237609 121961 237637 121989
rect 237671 121961 237699 121989
rect 237485 113147 237513 113175
rect 237547 113147 237575 113175
rect 237609 113147 237637 113175
rect 237671 113147 237699 113175
rect 237485 113085 237513 113113
rect 237547 113085 237575 113113
rect 237609 113085 237637 113113
rect 237671 113085 237699 113113
rect 237485 113023 237513 113051
rect 237547 113023 237575 113051
rect 237609 113023 237637 113051
rect 237671 113023 237699 113051
rect 237485 112961 237513 112989
rect 237547 112961 237575 112989
rect 237609 112961 237637 112989
rect 237671 112961 237699 112989
rect 237485 104147 237513 104175
rect 237547 104147 237575 104175
rect 237609 104147 237637 104175
rect 237671 104147 237699 104175
rect 237485 104085 237513 104113
rect 237547 104085 237575 104113
rect 237609 104085 237637 104113
rect 237671 104085 237699 104113
rect 237485 104023 237513 104051
rect 237547 104023 237575 104051
rect 237609 104023 237637 104051
rect 237671 104023 237699 104051
rect 237485 103961 237513 103989
rect 237547 103961 237575 103989
rect 237609 103961 237637 103989
rect 237671 103961 237699 103989
rect 237485 95147 237513 95175
rect 237547 95147 237575 95175
rect 237609 95147 237637 95175
rect 237671 95147 237699 95175
rect 237485 95085 237513 95113
rect 237547 95085 237575 95113
rect 237609 95085 237637 95113
rect 237671 95085 237699 95113
rect 237485 95023 237513 95051
rect 237547 95023 237575 95051
rect 237609 95023 237637 95051
rect 237671 95023 237699 95051
rect 237485 94961 237513 94989
rect 237547 94961 237575 94989
rect 237609 94961 237637 94989
rect 237671 94961 237699 94989
rect 237485 86147 237513 86175
rect 237547 86147 237575 86175
rect 237609 86147 237637 86175
rect 237671 86147 237699 86175
rect 237485 86085 237513 86113
rect 237547 86085 237575 86113
rect 237609 86085 237637 86113
rect 237671 86085 237699 86113
rect 237485 86023 237513 86051
rect 237547 86023 237575 86051
rect 237609 86023 237637 86051
rect 237671 86023 237699 86051
rect 237485 85961 237513 85989
rect 237547 85961 237575 85989
rect 237609 85961 237637 85989
rect 237671 85961 237699 85989
rect 237485 77147 237513 77175
rect 237547 77147 237575 77175
rect 237609 77147 237637 77175
rect 237671 77147 237699 77175
rect 237485 77085 237513 77113
rect 237547 77085 237575 77113
rect 237609 77085 237637 77113
rect 237671 77085 237699 77113
rect 237485 77023 237513 77051
rect 237547 77023 237575 77051
rect 237609 77023 237637 77051
rect 237671 77023 237699 77051
rect 237485 76961 237513 76989
rect 237547 76961 237575 76989
rect 237609 76961 237637 76989
rect 237671 76961 237699 76989
rect 237485 68147 237513 68175
rect 237547 68147 237575 68175
rect 237609 68147 237637 68175
rect 237671 68147 237699 68175
rect 237485 68085 237513 68113
rect 237547 68085 237575 68113
rect 237609 68085 237637 68113
rect 237671 68085 237699 68113
rect 237485 68023 237513 68051
rect 237547 68023 237575 68051
rect 237609 68023 237637 68051
rect 237671 68023 237699 68051
rect 237485 67961 237513 67989
rect 237547 67961 237575 67989
rect 237609 67961 237637 67989
rect 237671 67961 237699 67989
rect 237485 59147 237513 59175
rect 237547 59147 237575 59175
rect 237609 59147 237637 59175
rect 237671 59147 237699 59175
rect 237485 59085 237513 59113
rect 237547 59085 237575 59113
rect 237609 59085 237637 59113
rect 237671 59085 237699 59113
rect 237485 59023 237513 59051
rect 237547 59023 237575 59051
rect 237609 59023 237637 59051
rect 237671 59023 237699 59051
rect 237485 58961 237513 58989
rect 237547 58961 237575 58989
rect 237609 58961 237637 58989
rect 237671 58961 237699 58989
rect 237485 50147 237513 50175
rect 237547 50147 237575 50175
rect 237609 50147 237637 50175
rect 237671 50147 237699 50175
rect 237485 50085 237513 50113
rect 237547 50085 237575 50113
rect 237609 50085 237637 50113
rect 237671 50085 237699 50113
rect 237485 50023 237513 50051
rect 237547 50023 237575 50051
rect 237609 50023 237637 50051
rect 237671 50023 237699 50051
rect 237485 49961 237513 49989
rect 237547 49961 237575 49989
rect 237609 49961 237637 49989
rect 237671 49961 237699 49989
rect 237485 41147 237513 41175
rect 237547 41147 237575 41175
rect 237609 41147 237637 41175
rect 237671 41147 237699 41175
rect 237485 41085 237513 41113
rect 237547 41085 237575 41113
rect 237609 41085 237637 41113
rect 237671 41085 237699 41113
rect 237485 41023 237513 41051
rect 237547 41023 237575 41051
rect 237609 41023 237637 41051
rect 237671 41023 237699 41051
rect 237485 40961 237513 40989
rect 237547 40961 237575 40989
rect 237609 40961 237637 40989
rect 237671 40961 237699 40989
rect 237485 32147 237513 32175
rect 237547 32147 237575 32175
rect 237609 32147 237637 32175
rect 237671 32147 237699 32175
rect 237485 32085 237513 32113
rect 237547 32085 237575 32113
rect 237609 32085 237637 32113
rect 237671 32085 237699 32113
rect 237485 32023 237513 32051
rect 237547 32023 237575 32051
rect 237609 32023 237637 32051
rect 237671 32023 237699 32051
rect 237485 31961 237513 31989
rect 237547 31961 237575 31989
rect 237609 31961 237637 31989
rect 237671 31961 237699 31989
rect 237485 23147 237513 23175
rect 237547 23147 237575 23175
rect 237609 23147 237637 23175
rect 237671 23147 237699 23175
rect 237485 23085 237513 23113
rect 237547 23085 237575 23113
rect 237609 23085 237637 23113
rect 237671 23085 237699 23113
rect 237485 23023 237513 23051
rect 237547 23023 237575 23051
rect 237609 23023 237637 23051
rect 237671 23023 237699 23051
rect 237485 22961 237513 22989
rect 237547 22961 237575 22989
rect 237609 22961 237637 22989
rect 237671 22961 237699 22989
rect 237485 14147 237513 14175
rect 237547 14147 237575 14175
rect 237609 14147 237637 14175
rect 237671 14147 237699 14175
rect 237485 14085 237513 14113
rect 237547 14085 237575 14113
rect 237609 14085 237637 14113
rect 237671 14085 237699 14113
rect 237485 14023 237513 14051
rect 237547 14023 237575 14051
rect 237609 14023 237637 14051
rect 237671 14023 237699 14051
rect 237485 13961 237513 13989
rect 237547 13961 237575 13989
rect 237609 13961 237637 13989
rect 237671 13961 237699 13989
rect 237485 5147 237513 5175
rect 237547 5147 237575 5175
rect 237609 5147 237637 5175
rect 237671 5147 237699 5175
rect 237485 5085 237513 5113
rect 237547 5085 237575 5113
rect 237609 5085 237637 5113
rect 237671 5085 237699 5113
rect 237485 5023 237513 5051
rect 237547 5023 237575 5051
rect 237609 5023 237637 5051
rect 237671 5023 237699 5051
rect 237485 4961 237513 4989
rect 237547 4961 237575 4989
rect 237609 4961 237637 4989
rect 237671 4961 237699 4989
rect 237485 -588 237513 -560
rect 237547 -588 237575 -560
rect 237609 -588 237637 -560
rect 237671 -588 237699 -560
rect 237485 -650 237513 -622
rect 237547 -650 237575 -622
rect 237609 -650 237637 -622
rect 237671 -650 237699 -622
rect 237485 -712 237513 -684
rect 237547 -712 237575 -684
rect 237609 -712 237637 -684
rect 237671 -712 237699 -684
rect 237485 -774 237513 -746
rect 237547 -774 237575 -746
rect 237609 -774 237637 -746
rect 237671 -774 237699 -746
rect 244625 298578 244653 298606
rect 244687 298578 244715 298606
rect 244749 298578 244777 298606
rect 244811 298578 244839 298606
rect 244625 298516 244653 298544
rect 244687 298516 244715 298544
rect 244749 298516 244777 298544
rect 244811 298516 244839 298544
rect 244625 298454 244653 298482
rect 244687 298454 244715 298482
rect 244749 298454 244777 298482
rect 244811 298454 244839 298482
rect 244625 298392 244653 298420
rect 244687 298392 244715 298420
rect 244749 298392 244777 298420
rect 244811 298392 244839 298420
rect 244625 290147 244653 290175
rect 244687 290147 244715 290175
rect 244749 290147 244777 290175
rect 244811 290147 244839 290175
rect 244625 290085 244653 290113
rect 244687 290085 244715 290113
rect 244749 290085 244777 290113
rect 244811 290085 244839 290113
rect 244625 290023 244653 290051
rect 244687 290023 244715 290051
rect 244749 290023 244777 290051
rect 244811 290023 244839 290051
rect 244625 289961 244653 289989
rect 244687 289961 244715 289989
rect 244749 289961 244777 289989
rect 244811 289961 244839 289989
rect 244625 281147 244653 281175
rect 244687 281147 244715 281175
rect 244749 281147 244777 281175
rect 244811 281147 244839 281175
rect 244625 281085 244653 281113
rect 244687 281085 244715 281113
rect 244749 281085 244777 281113
rect 244811 281085 244839 281113
rect 244625 281023 244653 281051
rect 244687 281023 244715 281051
rect 244749 281023 244777 281051
rect 244811 281023 244839 281051
rect 244625 280961 244653 280989
rect 244687 280961 244715 280989
rect 244749 280961 244777 280989
rect 244811 280961 244839 280989
rect 244625 272147 244653 272175
rect 244687 272147 244715 272175
rect 244749 272147 244777 272175
rect 244811 272147 244839 272175
rect 244625 272085 244653 272113
rect 244687 272085 244715 272113
rect 244749 272085 244777 272113
rect 244811 272085 244839 272113
rect 244625 272023 244653 272051
rect 244687 272023 244715 272051
rect 244749 272023 244777 272051
rect 244811 272023 244839 272051
rect 244625 271961 244653 271989
rect 244687 271961 244715 271989
rect 244749 271961 244777 271989
rect 244811 271961 244839 271989
rect 244625 263147 244653 263175
rect 244687 263147 244715 263175
rect 244749 263147 244777 263175
rect 244811 263147 244839 263175
rect 244625 263085 244653 263113
rect 244687 263085 244715 263113
rect 244749 263085 244777 263113
rect 244811 263085 244839 263113
rect 244625 263023 244653 263051
rect 244687 263023 244715 263051
rect 244749 263023 244777 263051
rect 244811 263023 244839 263051
rect 244625 262961 244653 262989
rect 244687 262961 244715 262989
rect 244749 262961 244777 262989
rect 244811 262961 244839 262989
rect 244625 254147 244653 254175
rect 244687 254147 244715 254175
rect 244749 254147 244777 254175
rect 244811 254147 244839 254175
rect 244625 254085 244653 254113
rect 244687 254085 244715 254113
rect 244749 254085 244777 254113
rect 244811 254085 244839 254113
rect 244625 254023 244653 254051
rect 244687 254023 244715 254051
rect 244749 254023 244777 254051
rect 244811 254023 244839 254051
rect 244625 253961 244653 253989
rect 244687 253961 244715 253989
rect 244749 253961 244777 253989
rect 244811 253961 244839 253989
rect 244625 245147 244653 245175
rect 244687 245147 244715 245175
rect 244749 245147 244777 245175
rect 244811 245147 244839 245175
rect 244625 245085 244653 245113
rect 244687 245085 244715 245113
rect 244749 245085 244777 245113
rect 244811 245085 244839 245113
rect 244625 245023 244653 245051
rect 244687 245023 244715 245051
rect 244749 245023 244777 245051
rect 244811 245023 244839 245051
rect 244625 244961 244653 244989
rect 244687 244961 244715 244989
rect 244749 244961 244777 244989
rect 244811 244961 244839 244989
rect 244625 236147 244653 236175
rect 244687 236147 244715 236175
rect 244749 236147 244777 236175
rect 244811 236147 244839 236175
rect 244625 236085 244653 236113
rect 244687 236085 244715 236113
rect 244749 236085 244777 236113
rect 244811 236085 244839 236113
rect 244625 236023 244653 236051
rect 244687 236023 244715 236051
rect 244749 236023 244777 236051
rect 244811 236023 244839 236051
rect 244625 235961 244653 235989
rect 244687 235961 244715 235989
rect 244749 235961 244777 235989
rect 244811 235961 244839 235989
rect 244625 227147 244653 227175
rect 244687 227147 244715 227175
rect 244749 227147 244777 227175
rect 244811 227147 244839 227175
rect 244625 227085 244653 227113
rect 244687 227085 244715 227113
rect 244749 227085 244777 227113
rect 244811 227085 244839 227113
rect 244625 227023 244653 227051
rect 244687 227023 244715 227051
rect 244749 227023 244777 227051
rect 244811 227023 244839 227051
rect 244625 226961 244653 226989
rect 244687 226961 244715 226989
rect 244749 226961 244777 226989
rect 244811 226961 244839 226989
rect 244625 218147 244653 218175
rect 244687 218147 244715 218175
rect 244749 218147 244777 218175
rect 244811 218147 244839 218175
rect 244625 218085 244653 218113
rect 244687 218085 244715 218113
rect 244749 218085 244777 218113
rect 244811 218085 244839 218113
rect 244625 218023 244653 218051
rect 244687 218023 244715 218051
rect 244749 218023 244777 218051
rect 244811 218023 244839 218051
rect 244625 217961 244653 217989
rect 244687 217961 244715 217989
rect 244749 217961 244777 217989
rect 244811 217961 244839 217989
rect 244625 209147 244653 209175
rect 244687 209147 244715 209175
rect 244749 209147 244777 209175
rect 244811 209147 244839 209175
rect 244625 209085 244653 209113
rect 244687 209085 244715 209113
rect 244749 209085 244777 209113
rect 244811 209085 244839 209113
rect 244625 209023 244653 209051
rect 244687 209023 244715 209051
rect 244749 209023 244777 209051
rect 244811 209023 244839 209051
rect 244625 208961 244653 208989
rect 244687 208961 244715 208989
rect 244749 208961 244777 208989
rect 244811 208961 244839 208989
rect 244625 200147 244653 200175
rect 244687 200147 244715 200175
rect 244749 200147 244777 200175
rect 244811 200147 244839 200175
rect 244625 200085 244653 200113
rect 244687 200085 244715 200113
rect 244749 200085 244777 200113
rect 244811 200085 244839 200113
rect 244625 200023 244653 200051
rect 244687 200023 244715 200051
rect 244749 200023 244777 200051
rect 244811 200023 244839 200051
rect 244625 199961 244653 199989
rect 244687 199961 244715 199989
rect 244749 199961 244777 199989
rect 244811 199961 244839 199989
rect 244625 191147 244653 191175
rect 244687 191147 244715 191175
rect 244749 191147 244777 191175
rect 244811 191147 244839 191175
rect 244625 191085 244653 191113
rect 244687 191085 244715 191113
rect 244749 191085 244777 191113
rect 244811 191085 244839 191113
rect 244625 191023 244653 191051
rect 244687 191023 244715 191051
rect 244749 191023 244777 191051
rect 244811 191023 244839 191051
rect 244625 190961 244653 190989
rect 244687 190961 244715 190989
rect 244749 190961 244777 190989
rect 244811 190961 244839 190989
rect 244625 182147 244653 182175
rect 244687 182147 244715 182175
rect 244749 182147 244777 182175
rect 244811 182147 244839 182175
rect 244625 182085 244653 182113
rect 244687 182085 244715 182113
rect 244749 182085 244777 182113
rect 244811 182085 244839 182113
rect 244625 182023 244653 182051
rect 244687 182023 244715 182051
rect 244749 182023 244777 182051
rect 244811 182023 244839 182051
rect 244625 181961 244653 181989
rect 244687 181961 244715 181989
rect 244749 181961 244777 181989
rect 244811 181961 244839 181989
rect 244625 173147 244653 173175
rect 244687 173147 244715 173175
rect 244749 173147 244777 173175
rect 244811 173147 244839 173175
rect 244625 173085 244653 173113
rect 244687 173085 244715 173113
rect 244749 173085 244777 173113
rect 244811 173085 244839 173113
rect 244625 173023 244653 173051
rect 244687 173023 244715 173051
rect 244749 173023 244777 173051
rect 244811 173023 244839 173051
rect 244625 172961 244653 172989
rect 244687 172961 244715 172989
rect 244749 172961 244777 172989
rect 244811 172961 244839 172989
rect 244625 164147 244653 164175
rect 244687 164147 244715 164175
rect 244749 164147 244777 164175
rect 244811 164147 244839 164175
rect 244625 164085 244653 164113
rect 244687 164085 244715 164113
rect 244749 164085 244777 164113
rect 244811 164085 244839 164113
rect 244625 164023 244653 164051
rect 244687 164023 244715 164051
rect 244749 164023 244777 164051
rect 244811 164023 244839 164051
rect 244625 163961 244653 163989
rect 244687 163961 244715 163989
rect 244749 163961 244777 163989
rect 244811 163961 244839 163989
rect 244625 155147 244653 155175
rect 244687 155147 244715 155175
rect 244749 155147 244777 155175
rect 244811 155147 244839 155175
rect 244625 155085 244653 155113
rect 244687 155085 244715 155113
rect 244749 155085 244777 155113
rect 244811 155085 244839 155113
rect 244625 155023 244653 155051
rect 244687 155023 244715 155051
rect 244749 155023 244777 155051
rect 244811 155023 244839 155051
rect 244625 154961 244653 154989
rect 244687 154961 244715 154989
rect 244749 154961 244777 154989
rect 244811 154961 244839 154989
rect 244625 146147 244653 146175
rect 244687 146147 244715 146175
rect 244749 146147 244777 146175
rect 244811 146147 244839 146175
rect 244625 146085 244653 146113
rect 244687 146085 244715 146113
rect 244749 146085 244777 146113
rect 244811 146085 244839 146113
rect 244625 146023 244653 146051
rect 244687 146023 244715 146051
rect 244749 146023 244777 146051
rect 244811 146023 244839 146051
rect 244625 145961 244653 145989
rect 244687 145961 244715 145989
rect 244749 145961 244777 145989
rect 244811 145961 244839 145989
rect 244625 137147 244653 137175
rect 244687 137147 244715 137175
rect 244749 137147 244777 137175
rect 244811 137147 244839 137175
rect 244625 137085 244653 137113
rect 244687 137085 244715 137113
rect 244749 137085 244777 137113
rect 244811 137085 244839 137113
rect 244625 137023 244653 137051
rect 244687 137023 244715 137051
rect 244749 137023 244777 137051
rect 244811 137023 244839 137051
rect 244625 136961 244653 136989
rect 244687 136961 244715 136989
rect 244749 136961 244777 136989
rect 244811 136961 244839 136989
rect 244625 128147 244653 128175
rect 244687 128147 244715 128175
rect 244749 128147 244777 128175
rect 244811 128147 244839 128175
rect 244625 128085 244653 128113
rect 244687 128085 244715 128113
rect 244749 128085 244777 128113
rect 244811 128085 244839 128113
rect 244625 128023 244653 128051
rect 244687 128023 244715 128051
rect 244749 128023 244777 128051
rect 244811 128023 244839 128051
rect 244625 127961 244653 127989
rect 244687 127961 244715 127989
rect 244749 127961 244777 127989
rect 244811 127961 244839 127989
rect 244625 119147 244653 119175
rect 244687 119147 244715 119175
rect 244749 119147 244777 119175
rect 244811 119147 244839 119175
rect 244625 119085 244653 119113
rect 244687 119085 244715 119113
rect 244749 119085 244777 119113
rect 244811 119085 244839 119113
rect 244625 119023 244653 119051
rect 244687 119023 244715 119051
rect 244749 119023 244777 119051
rect 244811 119023 244839 119051
rect 244625 118961 244653 118989
rect 244687 118961 244715 118989
rect 244749 118961 244777 118989
rect 244811 118961 244839 118989
rect 244625 110147 244653 110175
rect 244687 110147 244715 110175
rect 244749 110147 244777 110175
rect 244811 110147 244839 110175
rect 244625 110085 244653 110113
rect 244687 110085 244715 110113
rect 244749 110085 244777 110113
rect 244811 110085 244839 110113
rect 244625 110023 244653 110051
rect 244687 110023 244715 110051
rect 244749 110023 244777 110051
rect 244811 110023 244839 110051
rect 244625 109961 244653 109989
rect 244687 109961 244715 109989
rect 244749 109961 244777 109989
rect 244811 109961 244839 109989
rect 244625 101147 244653 101175
rect 244687 101147 244715 101175
rect 244749 101147 244777 101175
rect 244811 101147 244839 101175
rect 244625 101085 244653 101113
rect 244687 101085 244715 101113
rect 244749 101085 244777 101113
rect 244811 101085 244839 101113
rect 244625 101023 244653 101051
rect 244687 101023 244715 101051
rect 244749 101023 244777 101051
rect 244811 101023 244839 101051
rect 244625 100961 244653 100989
rect 244687 100961 244715 100989
rect 244749 100961 244777 100989
rect 244811 100961 244839 100989
rect 244625 92147 244653 92175
rect 244687 92147 244715 92175
rect 244749 92147 244777 92175
rect 244811 92147 244839 92175
rect 244625 92085 244653 92113
rect 244687 92085 244715 92113
rect 244749 92085 244777 92113
rect 244811 92085 244839 92113
rect 244625 92023 244653 92051
rect 244687 92023 244715 92051
rect 244749 92023 244777 92051
rect 244811 92023 244839 92051
rect 244625 91961 244653 91989
rect 244687 91961 244715 91989
rect 244749 91961 244777 91989
rect 244811 91961 244839 91989
rect 244625 83147 244653 83175
rect 244687 83147 244715 83175
rect 244749 83147 244777 83175
rect 244811 83147 244839 83175
rect 244625 83085 244653 83113
rect 244687 83085 244715 83113
rect 244749 83085 244777 83113
rect 244811 83085 244839 83113
rect 244625 83023 244653 83051
rect 244687 83023 244715 83051
rect 244749 83023 244777 83051
rect 244811 83023 244839 83051
rect 244625 82961 244653 82989
rect 244687 82961 244715 82989
rect 244749 82961 244777 82989
rect 244811 82961 244839 82989
rect 244625 74147 244653 74175
rect 244687 74147 244715 74175
rect 244749 74147 244777 74175
rect 244811 74147 244839 74175
rect 244625 74085 244653 74113
rect 244687 74085 244715 74113
rect 244749 74085 244777 74113
rect 244811 74085 244839 74113
rect 244625 74023 244653 74051
rect 244687 74023 244715 74051
rect 244749 74023 244777 74051
rect 244811 74023 244839 74051
rect 244625 73961 244653 73989
rect 244687 73961 244715 73989
rect 244749 73961 244777 73989
rect 244811 73961 244839 73989
rect 244625 65147 244653 65175
rect 244687 65147 244715 65175
rect 244749 65147 244777 65175
rect 244811 65147 244839 65175
rect 244625 65085 244653 65113
rect 244687 65085 244715 65113
rect 244749 65085 244777 65113
rect 244811 65085 244839 65113
rect 244625 65023 244653 65051
rect 244687 65023 244715 65051
rect 244749 65023 244777 65051
rect 244811 65023 244839 65051
rect 244625 64961 244653 64989
rect 244687 64961 244715 64989
rect 244749 64961 244777 64989
rect 244811 64961 244839 64989
rect 244625 56147 244653 56175
rect 244687 56147 244715 56175
rect 244749 56147 244777 56175
rect 244811 56147 244839 56175
rect 244625 56085 244653 56113
rect 244687 56085 244715 56113
rect 244749 56085 244777 56113
rect 244811 56085 244839 56113
rect 244625 56023 244653 56051
rect 244687 56023 244715 56051
rect 244749 56023 244777 56051
rect 244811 56023 244839 56051
rect 244625 55961 244653 55989
rect 244687 55961 244715 55989
rect 244749 55961 244777 55989
rect 244811 55961 244839 55989
rect 244625 47147 244653 47175
rect 244687 47147 244715 47175
rect 244749 47147 244777 47175
rect 244811 47147 244839 47175
rect 244625 47085 244653 47113
rect 244687 47085 244715 47113
rect 244749 47085 244777 47113
rect 244811 47085 244839 47113
rect 244625 47023 244653 47051
rect 244687 47023 244715 47051
rect 244749 47023 244777 47051
rect 244811 47023 244839 47051
rect 244625 46961 244653 46989
rect 244687 46961 244715 46989
rect 244749 46961 244777 46989
rect 244811 46961 244839 46989
rect 244625 38147 244653 38175
rect 244687 38147 244715 38175
rect 244749 38147 244777 38175
rect 244811 38147 244839 38175
rect 244625 38085 244653 38113
rect 244687 38085 244715 38113
rect 244749 38085 244777 38113
rect 244811 38085 244839 38113
rect 244625 38023 244653 38051
rect 244687 38023 244715 38051
rect 244749 38023 244777 38051
rect 244811 38023 244839 38051
rect 244625 37961 244653 37989
rect 244687 37961 244715 37989
rect 244749 37961 244777 37989
rect 244811 37961 244839 37989
rect 244625 29147 244653 29175
rect 244687 29147 244715 29175
rect 244749 29147 244777 29175
rect 244811 29147 244839 29175
rect 244625 29085 244653 29113
rect 244687 29085 244715 29113
rect 244749 29085 244777 29113
rect 244811 29085 244839 29113
rect 244625 29023 244653 29051
rect 244687 29023 244715 29051
rect 244749 29023 244777 29051
rect 244811 29023 244839 29051
rect 244625 28961 244653 28989
rect 244687 28961 244715 28989
rect 244749 28961 244777 28989
rect 244811 28961 244839 28989
rect 244625 20147 244653 20175
rect 244687 20147 244715 20175
rect 244749 20147 244777 20175
rect 244811 20147 244839 20175
rect 244625 20085 244653 20113
rect 244687 20085 244715 20113
rect 244749 20085 244777 20113
rect 244811 20085 244839 20113
rect 244625 20023 244653 20051
rect 244687 20023 244715 20051
rect 244749 20023 244777 20051
rect 244811 20023 244839 20051
rect 244625 19961 244653 19989
rect 244687 19961 244715 19989
rect 244749 19961 244777 19989
rect 244811 19961 244839 19989
rect 244625 11147 244653 11175
rect 244687 11147 244715 11175
rect 244749 11147 244777 11175
rect 244811 11147 244839 11175
rect 244625 11085 244653 11113
rect 244687 11085 244715 11113
rect 244749 11085 244777 11113
rect 244811 11085 244839 11113
rect 244625 11023 244653 11051
rect 244687 11023 244715 11051
rect 244749 11023 244777 11051
rect 244811 11023 244839 11051
rect 244625 10961 244653 10989
rect 244687 10961 244715 10989
rect 244749 10961 244777 10989
rect 244811 10961 244839 10989
rect 244625 2147 244653 2175
rect 244687 2147 244715 2175
rect 244749 2147 244777 2175
rect 244811 2147 244839 2175
rect 244625 2085 244653 2113
rect 244687 2085 244715 2113
rect 244749 2085 244777 2113
rect 244811 2085 244839 2113
rect 244625 2023 244653 2051
rect 244687 2023 244715 2051
rect 244749 2023 244777 2051
rect 244811 2023 244839 2051
rect 244625 1961 244653 1989
rect 244687 1961 244715 1989
rect 244749 1961 244777 1989
rect 244811 1961 244839 1989
rect 244625 -108 244653 -80
rect 244687 -108 244715 -80
rect 244749 -108 244777 -80
rect 244811 -108 244839 -80
rect 244625 -170 244653 -142
rect 244687 -170 244715 -142
rect 244749 -170 244777 -142
rect 244811 -170 244839 -142
rect 244625 -232 244653 -204
rect 244687 -232 244715 -204
rect 244749 -232 244777 -204
rect 244811 -232 244839 -204
rect 244625 -294 244653 -266
rect 244687 -294 244715 -266
rect 244749 -294 244777 -266
rect 244811 -294 244839 -266
rect 246485 299058 246513 299086
rect 246547 299058 246575 299086
rect 246609 299058 246637 299086
rect 246671 299058 246699 299086
rect 246485 298996 246513 299024
rect 246547 298996 246575 299024
rect 246609 298996 246637 299024
rect 246671 298996 246699 299024
rect 246485 298934 246513 298962
rect 246547 298934 246575 298962
rect 246609 298934 246637 298962
rect 246671 298934 246699 298962
rect 246485 298872 246513 298900
rect 246547 298872 246575 298900
rect 246609 298872 246637 298900
rect 246671 298872 246699 298900
rect 246485 293147 246513 293175
rect 246547 293147 246575 293175
rect 246609 293147 246637 293175
rect 246671 293147 246699 293175
rect 246485 293085 246513 293113
rect 246547 293085 246575 293113
rect 246609 293085 246637 293113
rect 246671 293085 246699 293113
rect 246485 293023 246513 293051
rect 246547 293023 246575 293051
rect 246609 293023 246637 293051
rect 246671 293023 246699 293051
rect 246485 292961 246513 292989
rect 246547 292961 246575 292989
rect 246609 292961 246637 292989
rect 246671 292961 246699 292989
rect 246485 284147 246513 284175
rect 246547 284147 246575 284175
rect 246609 284147 246637 284175
rect 246671 284147 246699 284175
rect 246485 284085 246513 284113
rect 246547 284085 246575 284113
rect 246609 284085 246637 284113
rect 246671 284085 246699 284113
rect 246485 284023 246513 284051
rect 246547 284023 246575 284051
rect 246609 284023 246637 284051
rect 246671 284023 246699 284051
rect 246485 283961 246513 283989
rect 246547 283961 246575 283989
rect 246609 283961 246637 283989
rect 246671 283961 246699 283989
rect 246485 275147 246513 275175
rect 246547 275147 246575 275175
rect 246609 275147 246637 275175
rect 246671 275147 246699 275175
rect 246485 275085 246513 275113
rect 246547 275085 246575 275113
rect 246609 275085 246637 275113
rect 246671 275085 246699 275113
rect 246485 275023 246513 275051
rect 246547 275023 246575 275051
rect 246609 275023 246637 275051
rect 246671 275023 246699 275051
rect 246485 274961 246513 274989
rect 246547 274961 246575 274989
rect 246609 274961 246637 274989
rect 246671 274961 246699 274989
rect 246485 266147 246513 266175
rect 246547 266147 246575 266175
rect 246609 266147 246637 266175
rect 246671 266147 246699 266175
rect 246485 266085 246513 266113
rect 246547 266085 246575 266113
rect 246609 266085 246637 266113
rect 246671 266085 246699 266113
rect 246485 266023 246513 266051
rect 246547 266023 246575 266051
rect 246609 266023 246637 266051
rect 246671 266023 246699 266051
rect 246485 265961 246513 265989
rect 246547 265961 246575 265989
rect 246609 265961 246637 265989
rect 246671 265961 246699 265989
rect 246485 257147 246513 257175
rect 246547 257147 246575 257175
rect 246609 257147 246637 257175
rect 246671 257147 246699 257175
rect 246485 257085 246513 257113
rect 246547 257085 246575 257113
rect 246609 257085 246637 257113
rect 246671 257085 246699 257113
rect 246485 257023 246513 257051
rect 246547 257023 246575 257051
rect 246609 257023 246637 257051
rect 246671 257023 246699 257051
rect 246485 256961 246513 256989
rect 246547 256961 246575 256989
rect 246609 256961 246637 256989
rect 246671 256961 246699 256989
rect 246485 248147 246513 248175
rect 246547 248147 246575 248175
rect 246609 248147 246637 248175
rect 246671 248147 246699 248175
rect 246485 248085 246513 248113
rect 246547 248085 246575 248113
rect 246609 248085 246637 248113
rect 246671 248085 246699 248113
rect 246485 248023 246513 248051
rect 246547 248023 246575 248051
rect 246609 248023 246637 248051
rect 246671 248023 246699 248051
rect 246485 247961 246513 247989
rect 246547 247961 246575 247989
rect 246609 247961 246637 247989
rect 246671 247961 246699 247989
rect 246485 239147 246513 239175
rect 246547 239147 246575 239175
rect 246609 239147 246637 239175
rect 246671 239147 246699 239175
rect 246485 239085 246513 239113
rect 246547 239085 246575 239113
rect 246609 239085 246637 239113
rect 246671 239085 246699 239113
rect 246485 239023 246513 239051
rect 246547 239023 246575 239051
rect 246609 239023 246637 239051
rect 246671 239023 246699 239051
rect 246485 238961 246513 238989
rect 246547 238961 246575 238989
rect 246609 238961 246637 238989
rect 246671 238961 246699 238989
rect 246485 230147 246513 230175
rect 246547 230147 246575 230175
rect 246609 230147 246637 230175
rect 246671 230147 246699 230175
rect 246485 230085 246513 230113
rect 246547 230085 246575 230113
rect 246609 230085 246637 230113
rect 246671 230085 246699 230113
rect 246485 230023 246513 230051
rect 246547 230023 246575 230051
rect 246609 230023 246637 230051
rect 246671 230023 246699 230051
rect 246485 229961 246513 229989
rect 246547 229961 246575 229989
rect 246609 229961 246637 229989
rect 246671 229961 246699 229989
rect 246485 221147 246513 221175
rect 246547 221147 246575 221175
rect 246609 221147 246637 221175
rect 246671 221147 246699 221175
rect 246485 221085 246513 221113
rect 246547 221085 246575 221113
rect 246609 221085 246637 221113
rect 246671 221085 246699 221113
rect 246485 221023 246513 221051
rect 246547 221023 246575 221051
rect 246609 221023 246637 221051
rect 246671 221023 246699 221051
rect 246485 220961 246513 220989
rect 246547 220961 246575 220989
rect 246609 220961 246637 220989
rect 246671 220961 246699 220989
rect 246485 212147 246513 212175
rect 246547 212147 246575 212175
rect 246609 212147 246637 212175
rect 246671 212147 246699 212175
rect 246485 212085 246513 212113
rect 246547 212085 246575 212113
rect 246609 212085 246637 212113
rect 246671 212085 246699 212113
rect 246485 212023 246513 212051
rect 246547 212023 246575 212051
rect 246609 212023 246637 212051
rect 246671 212023 246699 212051
rect 246485 211961 246513 211989
rect 246547 211961 246575 211989
rect 246609 211961 246637 211989
rect 246671 211961 246699 211989
rect 246485 203147 246513 203175
rect 246547 203147 246575 203175
rect 246609 203147 246637 203175
rect 246671 203147 246699 203175
rect 246485 203085 246513 203113
rect 246547 203085 246575 203113
rect 246609 203085 246637 203113
rect 246671 203085 246699 203113
rect 246485 203023 246513 203051
rect 246547 203023 246575 203051
rect 246609 203023 246637 203051
rect 246671 203023 246699 203051
rect 246485 202961 246513 202989
rect 246547 202961 246575 202989
rect 246609 202961 246637 202989
rect 246671 202961 246699 202989
rect 246485 194147 246513 194175
rect 246547 194147 246575 194175
rect 246609 194147 246637 194175
rect 246671 194147 246699 194175
rect 246485 194085 246513 194113
rect 246547 194085 246575 194113
rect 246609 194085 246637 194113
rect 246671 194085 246699 194113
rect 246485 194023 246513 194051
rect 246547 194023 246575 194051
rect 246609 194023 246637 194051
rect 246671 194023 246699 194051
rect 246485 193961 246513 193989
rect 246547 193961 246575 193989
rect 246609 193961 246637 193989
rect 246671 193961 246699 193989
rect 246485 185147 246513 185175
rect 246547 185147 246575 185175
rect 246609 185147 246637 185175
rect 246671 185147 246699 185175
rect 246485 185085 246513 185113
rect 246547 185085 246575 185113
rect 246609 185085 246637 185113
rect 246671 185085 246699 185113
rect 246485 185023 246513 185051
rect 246547 185023 246575 185051
rect 246609 185023 246637 185051
rect 246671 185023 246699 185051
rect 246485 184961 246513 184989
rect 246547 184961 246575 184989
rect 246609 184961 246637 184989
rect 246671 184961 246699 184989
rect 246485 176147 246513 176175
rect 246547 176147 246575 176175
rect 246609 176147 246637 176175
rect 246671 176147 246699 176175
rect 246485 176085 246513 176113
rect 246547 176085 246575 176113
rect 246609 176085 246637 176113
rect 246671 176085 246699 176113
rect 246485 176023 246513 176051
rect 246547 176023 246575 176051
rect 246609 176023 246637 176051
rect 246671 176023 246699 176051
rect 246485 175961 246513 175989
rect 246547 175961 246575 175989
rect 246609 175961 246637 175989
rect 246671 175961 246699 175989
rect 246485 167147 246513 167175
rect 246547 167147 246575 167175
rect 246609 167147 246637 167175
rect 246671 167147 246699 167175
rect 246485 167085 246513 167113
rect 246547 167085 246575 167113
rect 246609 167085 246637 167113
rect 246671 167085 246699 167113
rect 246485 167023 246513 167051
rect 246547 167023 246575 167051
rect 246609 167023 246637 167051
rect 246671 167023 246699 167051
rect 246485 166961 246513 166989
rect 246547 166961 246575 166989
rect 246609 166961 246637 166989
rect 246671 166961 246699 166989
rect 246485 158147 246513 158175
rect 246547 158147 246575 158175
rect 246609 158147 246637 158175
rect 246671 158147 246699 158175
rect 246485 158085 246513 158113
rect 246547 158085 246575 158113
rect 246609 158085 246637 158113
rect 246671 158085 246699 158113
rect 246485 158023 246513 158051
rect 246547 158023 246575 158051
rect 246609 158023 246637 158051
rect 246671 158023 246699 158051
rect 246485 157961 246513 157989
rect 246547 157961 246575 157989
rect 246609 157961 246637 157989
rect 246671 157961 246699 157989
rect 246485 149147 246513 149175
rect 246547 149147 246575 149175
rect 246609 149147 246637 149175
rect 246671 149147 246699 149175
rect 246485 149085 246513 149113
rect 246547 149085 246575 149113
rect 246609 149085 246637 149113
rect 246671 149085 246699 149113
rect 246485 149023 246513 149051
rect 246547 149023 246575 149051
rect 246609 149023 246637 149051
rect 246671 149023 246699 149051
rect 246485 148961 246513 148989
rect 246547 148961 246575 148989
rect 246609 148961 246637 148989
rect 246671 148961 246699 148989
rect 246485 140147 246513 140175
rect 246547 140147 246575 140175
rect 246609 140147 246637 140175
rect 246671 140147 246699 140175
rect 246485 140085 246513 140113
rect 246547 140085 246575 140113
rect 246609 140085 246637 140113
rect 246671 140085 246699 140113
rect 246485 140023 246513 140051
rect 246547 140023 246575 140051
rect 246609 140023 246637 140051
rect 246671 140023 246699 140051
rect 246485 139961 246513 139989
rect 246547 139961 246575 139989
rect 246609 139961 246637 139989
rect 246671 139961 246699 139989
rect 246485 131147 246513 131175
rect 246547 131147 246575 131175
rect 246609 131147 246637 131175
rect 246671 131147 246699 131175
rect 246485 131085 246513 131113
rect 246547 131085 246575 131113
rect 246609 131085 246637 131113
rect 246671 131085 246699 131113
rect 246485 131023 246513 131051
rect 246547 131023 246575 131051
rect 246609 131023 246637 131051
rect 246671 131023 246699 131051
rect 246485 130961 246513 130989
rect 246547 130961 246575 130989
rect 246609 130961 246637 130989
rect 246671 130961 246699 130989
rect 246485 122147 246513 122175
rect 246547 122147 246575 122175
rect 246609 122147 246637 122175
rect 246671 122147 246699 122175
rect 246485 122085 246513 122113
rect 246547 122085 246575 122113
rect 246609 122085 246637 122113
rect 246671 122085 246699 122113
rect 246485 122023 246513 122051
rect 246547 122023 246575 122051
rect 246609 122023 246637 122051
rect 246671 122023 246699 122051
rect 246485 121961 246513 121989
rect 246547 121961 246575 121989
rect 246609 121961 246637 121989
rect 246671 121961 246699 121989
rect 246485 113147 246513 113175
rect 246547 113147 246575 113175
rect 246609 113147 246637 113175
rect 246671 113147 246699 113175
rect 246485 113085 246513 113113
rect 246547 113085 246575 113113
rect 246609 113085 246637 113113
rect 246671 113085 246699 113113
rect 246485 113023 246513 113051
rect 246547 113023 246575 113051
rect 246609 113023 246637 113051
rect 246671 113023 246699 113051
rect 246485 112961 246513 112989
rect 246547 112961 246575 112989
rect 246609 112961 246637 112989
rect 246671 112961 246699 112989
rect 246485 104147 246513 104175
rect 246547 104147 246575 104175
rect 246609 104147 246637 104175
rect 246671 104147 246699 104175
rect 246485 104085 246513 104113
rect 246547 104085 246575 104113
rect 246609 104085 246637 104113
rect 246671 104085 246699 104113
rect 246485 104023 246513 104051
rect 246547 104023 246575 104051
rect 246609 104023 246637 104051
rect 246671 104023 246699 104051
rect 246485 103961 246513 103989
rect 246547 103961 246575 103989
rect 246609 103961 246637 103989
rect 246671 103961 246699 103989
rect 246485 95147 246513 95175
rect 246547 95147 246575 95175
rect 246609 95147 246637 95175
rect 246671 95147 246699 95175
rect 246485 95085 246513 95113
rect 246547 95085 246575 95113
rect 246609 95085 246637 95113
rect 246671 95085 246699 95113
rect 246485 95023 246513 95051
rect 246547 95023 246575 95051
rect 246609 95023 246637 95051
rect 246671 95023 246699 95051
rect 246485 94961 246513 94989
rect 246547 94961 246575 94989
rect 246609 94961 246637 94989
rect 246671 94961 246699 94989
rect 246485 86147 246513 86175
rect 246547 86147 246575 86175
rect 246609 86147 246637 86175
rect 246671 86147 246699 86175
rect 246485 86085 246513 86113
rect 246547 86085 246575 86113
rect 246609 86085 246637 86113
rect 246671 86085 246699 86113
rect 246485 86023 246513 86051
rect 246547 86023 246575 86051
rect 246609 86023 246637 86051
rect 246671 86023 246699 86051
rect 246485 85961 246513 85989
rect 246547 85961 246575 85989
rect 246609 85961 246637 85989
rect 246671 85961 246699 85989
rect 246485 77147 246513 77175
rect 246547 77147 246575 77175
rect 246609 77147 246637 77175
rect 246671 77147 246699 77175
rect 246485 77085 246513 77113
rect 246547 77085 246575 77113
rect 246609 77085 246637 77113
rect 246671 77085 246699 77113
rect 246485 77023 246513 77051
rect 246547 77023 246575 77051
rect 246609 77023 246637 77051
rect 246671 77023 246699 77051
rect 246485 76961 246513 76989
rect 246547 76961 246575 76989
rect 246609 76961 246637 76989
rect 246671 76961 246699 76989
rect 246485 68147 246513 68175
rect 246547 68147 246575 68175
rect 246609 68147 246637 68175
rect 246671 68147 246699 68175
rect 246485 68085 246513 68113
rect 246547 68085 246575 68113
rect 246609 68085 246637 68113
rect 246671 68085 246699 68113
rect 246485 68023 246513 68051
rect 246547 68023 246575 68051
rect 246609 68023 246637 68051
rect 246671 68023 246699 68051
rect 246485 67961 246513 67989
rect 246547 67961 246575 67989
rect 246609 67961 246637 67989
rect 246671 67961 246699 67989
rect 246485 59147 246513 59175
rect 246547 59147 246575 59175
rect 246609 59147 246637 59175
rect 246671 59147 246699 59175
rect 246485 59085 246513 59113
rect 246547 59085 246575 59113
rect 246609 59085 246637 59113
rect 246671 59085 246699 59113
rect 246485 59023 246513 59051
rect 246547 59023 246575 59051
rect 246609 59023 246637 59051
rect 246671 59023 246699 59051
rect 246485 58961 246513 58989
rect 246547 58961 246575 58989
rect 246609 58961 246637 58989
rect 246671 58961 246699 58989
rect 246485 50147 246513 50175
rect 246547 50147 246575 50175
rect 246609 50147 246637 50175
rect 246671 50147 246699 50175
rect 246485 50085 246513 50113
rect 246547 50085 246575 50113
rect 246609 50085 246637 50113
rect 246671 50085 246699 50113
rect 246485 50023 246513 50051
rect 246547 50023 246575 50051
rect 246609 50023 246637 50051
rect 246671 50023 246699 50051
rect 246485 49961 246513 49989
rect 246547 49961 246575 49989
rect 246609 49961 246637 49989
rect 246671 49961 246699 49989
rect 246485 41147 246513 41175
rect 246547 41147 246575 41175
rect 246609 41147 246637 41175
rect 246671 41147 246699 41175
rect 246485 41085 246513 41113
rect 246547 41085 246575 41113
rect 246609 41085 246637 41113
rect 246671 41085 246699 41113
rect 246485 41023 246513 41051
rect 246547 41023 246575 41051
rect 246609 41023 246637 41051
rect 246671 41023 246699 41051
rect 246485 40961 246513 40989
rect 246547 40961 246575 40989
rect 246609 40961 246637 40989
rect 246671 40961 246699 40989
rect 246485 32147 246513 32175
rect 246547 32147 246575 32175
rect 246609 32147 246637 32175
rect 246671 32147 246699 32175
rect 246485 32085 246513 32113
rect 246547 32085 246575 32113
rect 246609 32085 246637 32113
rect 246671 32085 246699 32113
rect 246485 32023 246513 32051
rect 246547 32023 246575 32051
rect 246609 32023 246637 32051
rect 246671 32023 246699 32051
rect 246485 31961 246513 31989
rect 246547 31961 246575 31989
rect 246609 31961 246637 31989
rect 246671 31961 246699 31989
rect 246485 23147 246513 23175
rect 246547 23147 246575 23175
rect 246609 23147 246637 23175
rect 246671 23147 246699 23175
rect 246485 23085 246513 23113
rect 246547 23085 246575 23113
rect 246609 23085 246637 23113
rect 246671 23085 246699 23113
rect 246485 23023 246513 23051
rect 246547 23023 246575 23051
rect 246609 23023 246637 23051
rect 246671 23023 246699 23051
rect 246485 22961 246513 22989
rect 246547 22961 246575 22989
rect 246609 22961 246637 22989
rect 246671 22961 246699 22989
rect 246485 14147 246513 14175
rect 246547 14147 246575 14175
rect 246609 14147 246637 14175
rect 246671 14147 246699 14175
rect 246485 14085 246513 14113
rect 246547 14085 246575 14113
rect 246609 14085 246637 14113
rect 246671 14085 246699 14113
rect 246485 14023 246513 14051
rect 246547 14023 246575 14051
rect 246609 14023 246637 14051
rect 246671 14023 246699 14051
rect 246485 13961 246513 13989
rect 246547 13961 246575 13989
rect 246609 13961 246637 13989
rect 246671 13961 246699 13989
rect 246485 5147 246513 5175
rect 246547 5147 246575 5175
rect 246609 5147 246637 5175
rect 246671 5147 246699 5175
rect 246485 5085 246513 5113
rect 246547 5085 246575 5113
rect 246609 5085 246637 5113
rect 246671 5085 246699 5113
rect 246485 5023 246513 5051
rect 246547 5023 246575 5051
rect 246609 5023 246637 5051
rect 246671 5023 246699 5051
rect 246485 4961 246513 4989
rect 246547 4961 246575 4989
rect 246609 4961 246637 4989
rect 246671 4961 246699 4989
rect 246485 -588 246513 -560
rect 246547 -588 246575 -560
rect 246609 -588 246637 -560
rect 246671 -588 246699 -560
rect 246485 -650 246513 -622
rect 246547 -650 246575 -622
rect 246609 -650 246637 -622
rect 246671 -650 246699 -622
rect 246485 -712 246513 -684
rect 246547 -712 246575 -684
rect 246609 -712 246637 -684
rect 246671 -712 246699 -684
rect 246485 -774 246513 -746
rect 246547 -774 246575 -746
rect 246609 -774 246637 -746
rect 246671 -774 246699 -746
rect 253625 298578 253653 298606
rect 253687 298578 253715 298606
rect 253749 298578 253777 298606
rect 253811 298578 253839 298606
rect 253625 298516 253653 298544
rect 253687 298516 253715 298544
rect 253749 298516 253777 298544
rect 253811 298516 253839 298544
rect 253625 298454 253653 298482
rect 253687 298454 253715 298482
rect 253749 298454 253777 298482
rect 253811 298454 253839 298482
rect 253625 298392 253653 298420
rect 253687 298392 253715 298420
rect 253749 298392 253777 298420
rect 253811 298392 253839 298420
rect 253625 290147 253653 290175
rect 253687 290147 253715 290175
rect 253749 290147 253777 290175
rect 253811 290147 253839 290175
rect 253625 290085 253653 290113
rect 253687 290085 253715 290113
rect 253749 290085 253777 290113
rect 253811 290085 253839 290113
rect 253625 290023 253653 290051
rect 253687 290023 253715 290051
rect 253749 290023 253777 290051
rect 253811 290023 253839 290051
rect 253625 289961 253653 289989
rect 253687 289961 253715 289989
rect 253749 289961 253777 289989
rect 253811 289961 253839 289989
rect 253625 281147 253653 281175
rect 253687 281147 253715 281175
rect 253749 281147 253777 281175
rect 253811 281147 253839 281175
rect 253625 281085 253653 281113
rect 253687 281085 253715 281113
rect 253749 281085 253777 281113
rect 253811 281085 253839 281113
rect 253625 281023 253653 281051
rect 253687 281023 253715 281051
rect 253749 281023 253777 281051
rect 253811 281023 253839 281051
rect 253625 280961 253653 280989
rect 253687 280961 253715 280989
rect 253749 280961 253777 280989
rect 253811 280961 253839 280989
rect 253625 272147 253653 272175
rect 253687 272147 253715 272175
rect 253749 272147 253777 272175
rect 253811 272147 253839 272175
rect 253625 272085 253653 272113
rect 253687 272085 253715 272113
rect 253749 272085 253777 272113
rect 253811 272085 253839 272113
rect 253625 272023 253653 272051
rect 253687 272023 253715 272051
rect 253749 272023 253777 272051
rect 253811 272023 253839 272051
rect 253625 271961 253653 271989
rect 253687 271961 253715 271989
rect 253749 271961 253777 271989
rect 253811 271961 253839 271989
rect 253625 263147 253653 263175
rect 253687 263147 253715 263175
rect 253749 263147 253777 263175
rect 253811 263147 253839 263175
rect 253625 263085 253653 263113
rect 253687 263085 253715 263113
rect 253749 263085 253777 263113
rect 253811 263085 253839 263113
rect 253625 263023 253653 263051
rect 253687 263023 253715 263051
rect 253749 263023 253777 263051
rect 253811 263023 253839 263051
rect 253625 262961 253653 262989
rect 253687 262961 253715 262989
rect 253749 262961 253777 262989
rect 253811 262961 253839 262989
rect 253625 254147 253653 254175
rect 253687 254147 253715 254175
rect 253749 254147 253777 254175
rect 253811 254147 253839 254175
rect 253625 254085 253653 254113
rect 253687 254085 253715 254113
rect 253749 254085 253777 254113
rect 253811 254085 253839 254113
rect 253625 254023 253653 254051
rect 253687 254023 253715 254051
rect 253749 254023 253777 254051
rect 253811 254023 253839 254051
rect 253625 253961 253653 253989
rect 253687 253961 253715 253989
rect 253749 253961 253777 253989
rect 253811 253961 253839 253989
rect 253625 245147 253653 245175
rect 253687 245147 253715 245175
rect 253749 245147 253777 245175
rect 253811 245147 253839 245175
rect 253625 245085 253653 245113
rect 253687 245085 253715 245113
rect 253749 245085 253777 245113
rect 253811 245085 253839 245113
rect 253625 245023 253653 245051
rect 253687 245023 253715 245051
rect 253749 245023 253777 245051
rect 253811 245023 253839 245051
rect 253625 244961 253653 244989
rect 253687 244961 253715 244989
rect 253749 244961 253777 244989
rect 253811 244961 253839 244989
rect 253625 236147 253653 236175
rect 253687 236147 253715 236175
rect 253749 236147 253777 236175
rect 253811 236147 253839 236175
rect 253625 236085 253653 236113
rect 253687 236085 253715 236113
rect 253749 236085 253777 236113
rect 253811 236085 253839 236113
rect 253625 236023 253653 236051
rect 253687 236023 253715 236051
rect 253749 236023 253777 236051
rect 253811 236023 253839 236051
rect 253625 235961 253653 235989
rect 253687 235961 253715 235989
rect 253749 235961 253777 235989
rect 253811 235961 253839 235989
rect 253625 227147 253653 227175
rect 253687 227147 253715 227175
rect 253749 227147 253777 227175
rect 253811 227147 253839 227175
rect 253625 227085 253653 227113
rect 253687 227085 253715 227113
rect 253749 227085 253777 227113
rect 253811 227085 253839 227113
rect 253625 227023 253653 227051
rect 253687 227023 253715 227051
rect 253749 227023 253777 227051
rect 253811 227023 253839 227051
rect 253625 226961 253653 226989
rect 253687 226961 253715 226989
rect 253749 226961 253777 226989
rect 253811 226961 253839 226989
rect 253625 218147 253653 218175
rect 253687 218147 253715 218175
rect 253749 218147 253777 218175
rect 253811 218147 253839 218175
rect 253625 218085 253653 218113
rect 253687 218085 253715 218113
rect 253749 218085 253777 218113
rect 253811 218085 253839 218113
rect 253625 218023 253653 218051
rect 253687 218023 253715 218051
rect 253749 218023 253777 218051
rect 253811 218023 253839 218051
rect 253625 217961 253653 217989
rect 253687 217961 253715 217989
rect 253749 217961 253777 217989
rect 253811 217961 253839 217989
rect 253625 209147 253653 209175
rect 253687 209147 253715 209175
rect 253749 209147 253777 209175
rect 253811 209147 253839 209175
rect 253625 209085 253653 209113
rect 253687 209085 253715 209113
rect 253749 209085 253777 209113
rect 253811 209085 253839 209113
rect 253625 209023 253653 209051
rect 253687 209023 253715 209051
rect 253749 209023 253777 209051
rect 253811 209023 253839 209051
rect 253625 208961 253653 208989
rect 253687 208961 253715 208989
rect 253749 208961 253777 208989
rect 253811 208961 253839 208989
rect 253625 200147 253653 200175
rect 253687 200147 253715 200175
rect 253749 200147 253777 200175
rect 253811 200147 253839 200175
rect 253625 200085 253653 200113
rect 253687 200085 253715 200113
rect 253749 200085 253777 200113
rect 253811 200085 253839 200113
rect 253625 200023 253653 200051
rect 253687 200023 253715 200051
rect 253749 200023 253777 200051
rect 253811 200023 253839 200051
rect 253625 199961 253653 199989
rect 253687 199961 253715 199989
rect 253749 199961 253777 199989
rect 253811 199961 253839 199989
rect 253625 191147 253653 191175
rect 253687 191147 253715 191175
rect 253749 191147 253777 191175
rect 253811 191147 253839 191175
rect 253625 191085 253653 191113
rect 253687 191085 253715 191113
rect 253749 191085 253777 191113
rect 253811 191085 253839 191113
rect 253625 191023 253653 191051
rect 253687 191023 253715 191051
rect 253749 191023 253777 191051
rect 253811 191023 253839 191051
rect 253625 190961 253653 190989
rect 253687 190961 253715 190989
rect 253749 190961 253777 190989
rect 253811 190961 253839 190989
rect 253625 182147 253653 182175
rect 253687 182147 253715 182175
rect 253749 182147 253777 182175
rect 253811 182147 253839 182175
rect 253625 182085 253653 182113
rect 253687 182085 253715 182113
rect 253749 182085 253777 182113
rect 253811 182085 253839 182113
rect 253625 182023 253653 182051
rect 253687 182023 253715 182051
rect 253749 182023 253777 182051
rect 253811 182023 253839 182051
rect 253625 181961 253653 181989
rect 253687 181961 253715 181989
rect 253749 181961 253777 181989
rect 253811 181961 253839 181989
rect 253625 173147 253653 173175
rect 253687 173147 253715 173175
rect 253749 173147 253777 173175
rect 253811 173147 253839 173175
rect 253625 173085 253653 173113
rect 253687 173085 253715 173113
rect 253749 173085 253777 173113
rect 253811 173085 253839 173113
rect 253625 173023 253653 173051
rect 253687 173023 253715 173051
rect 253749 173023 253777 173051
rect 253811 173023 253839 173051
rect 253625 172961 253653 172989
rect 253687 172961 253715 172989
rect 253749 172961 253777 172989
rect 253811 172961 253839 172989
rect 253625 164147 253653 164175
rect 253687 164147 253715 164175
rect 253749 164147 253777 164175
rect 253811 164147 253839 164175
rect 253625 164085 253653 164113
rect 253687 164085 253715 164113
rect 253749 164085 253777 164113
rect 253811 164085 253839 164113
rect 253625 164023 253653 164051
rect 253687 164023 253715 164051
rect 253749 164023 253777 164051
rect 253811 164023 253839 164051
rect 253625 163961 253653 163989
rect 253687 163961 253715 163989
rect 253749 163961 253777 163989
rect 253811 163961 253839 163989
rect 253625 155147 253653 155175
rect 253687 155147 253715 155175
rect 253749 155147 253777 155175
rect 253811 155147 253839 155175
rect 253625 155085 253653 155113
rect 253687 155085 253715 155113
rect 253749 155085 253777 155113
rect 253811 155085 253839 155113
rect 253625 155023 253653 155051
rect 253687 155023 253715 155051
rect 253749 155023 253777 155051
rect 253811 155023 253839 155051
rect 253625 154961 253653 154989
rect 253687 154961 253715 154989
rect 253749 154961 253777 154989
rect 253811 154961 253839 154989
rect 253625 146147 253653 146175
rect 253687 146147 253715 146175
rect 253749 146147 253777 146175
rect 253811 146147 253839 146175
rect 253625 146085 253653 146113
rect 253687 146085 253715 146113
rect 253749 146085 253777 146113
rect 253811 146085 253839 146113
rect 253625 146023 253653 146051
rect 253687 146023 253715 146051
rect 253749 146023 253777 146051
rect 253811 146023 253839 146051
rect 253625 145961 253653 145989
rect 253687 145961 253715 145989
rect 253749 145961 253777 145989
rect 253811 145961 253839 145989
rect 253625 137147 253653 137175
rect 253687 137147 253715 137175
rect 253749 137147 253777 137175
rect 253811 137147 253839 137175
rect 253625 137085 253653 137113
rect 253687 137085 253715 137113
rect 253749 137085 253777 137113
rect 253811 137085 253839 137113
rect 253625 137023 253653 137051
rect 253687 137023 253715 137051
rect 253749 137023 253777 137051
rect 253811 137023 253839 137051
rect 253625 136961 253653 136989
rect 253687 136961 253715 136989
rect 253749 136961 253777 136989
rect 253811 136961 253839 136989
rect 253625 128147 253653 128175
rect 253687 128147 253715 128175
rect 253749 128147 253777 128175
rect 253811 128147 253839 128175
rect 253625 128085 253653 128113
rect 253687 128085 253715 128113
rect 253749 128085 253777 128113
rect 253811 128085 253839 128113
rect 253625 128023 253653 128051
rect 253687 128023 253715 128051
rect 253749 128023 253777 128051
rect 253811 128023 253839 128051
rect 253625 127961 253653 127989
rect 253687 127961 253715 127989
rect 253749 127961 253777 127989
rect 253811 127961 253839 127989
rect 253625 119147 253653 119175
rect 253687 119147 253715 119175
rect 253749 119147 253777 119175
rect 253811 119147 253839 119175
rect 253625 119085 253653 119113
rect 253687 119085 253715 119113
rect 253749 119085 253777 119113
rect 253811 119085 253839 119113
rect 253625 119023 253653 119051
rect 253687 119023 253715 119051
rect 253749 119023 253777 119051
rect 253811 119023 253839 119051
rect 253625 118961 253653 118989
rect 253687 118961 253715 118989
rect 253749 118961 253777 118989
rect 253811 118961 253839 118989
rect 253625 110147 253653 110175
rect 253687 110147 253715 110175
rect 253749 110147 253777 110175
rect 253811 110147 253839 110175
rect 253625 110085 253653 110113
rect 253687 110085 253715 110113
rect 253749 110085 253777 110113
rect 253811 110085 253839 110113
rect 253625 110023 253653 110051
rect 253687 110023 253715 110051
rect 253749 110023 253777 110051
rect 253811 110023 253839 110051
rect 253625 109961 253653 109989
rect 253687 109961 253715 109989
rect 253749 109961 253777 109989
rect 253811 109961 253839 109989
rect 253625 101147 253653 101175
rect 253687 101147 253715 101175
rect 253749 101147 253777 101175
rect 253811 101147 253839 101175
rect 253625 101085 253653 101113
rect 253687 101085 253715 101113
rect 253749 101085 253777 101113
rect 253811 101085 253839 101113
rect 253625 101023 253653 101051
rect 253687 101023 253715 101051
rect 253749 101023 253777 101051
rect 253811 101023 253839 101051
rect 253625 100961 253653 100989
rect 253687 100961 253715 100989
rect 253749 100961 253777 100989
rect 253811 100961 253839 100989
rect 253625 92147 253653 92175
rect 253687 92147 253715 92175
rect 253749 92147 253777 92175
rect 253811 92147 253839 92175
rect 253625 92085 253653 92113
rect 253687 92085 253715 92113
rect 253749 92085 253777 92113
rect 253811 92085 253839 92113
rect 253625 92023 253653 92051
rect 253687 92023 253715 92051
rect 253749 92023 253777 92051
rect 253811 92023 253839 92051
rect 253625 91961 253653 91989
rect 253687 91961 253715 91989
rect 253749 91961 253777 91989
rect 253811 91961 253839 91989
rect 253625 83147 253653 83175
rect 253687 83147 253715 83175
rect 253749 83147 253777 83175
rect 253811 83147 253839 83175
rect 253625 83085 253653 83113
rect 253687 83085 253715 83113
rect 253749 83085 253777 83113
rect 253811 83085 253839 83113
rect 253625 83023 253653 83051
rect 253687 83023 253715 83051
rect 253749 83023 253777 83051
rect 253811 83023 253839 83051
rect 253625 82961 253653 82989
rect 253687 82961 253715 82989
rect 253749 82961 253777 82989
rect 253811 82961 253839 82989
rect 253625 74147 253653 74175
rect 253687 74147 253715 74175
rect 253749 74147 253777 74175
rect 253811 74147 253839 74175
rect 253625 74085 253653 74113
rect 253687 74085 253715 74113
rect 253749 74085 253777 74113
rect 253811 74085 253839 74113
rect 253625 74023 253653 74051
rect 253687 74023 253715 74051
rect 253749 74023 253777 74051
rect 253811 74023 253839 74051
rect 253625 73961 253653 73989
rect 253687 73961 253715 73989
rect 253749 73961 253777 73989
rect 253811 73961 253839 73989
rect 253625 65147 253653 65175
rect 253687 65147 253715 65175
rect 253749 65147 253777 65175
rect 253811 65147 253839 65175
rect 253625 65085 253653 65113
rect 253687 65085 253715 65113
rect 253749 65085 253777 65113
rect 253811 65085 253839 65113
rect 253625 65023 253653 65051
rect 253687 65023 253715 65051
rect 253749 65023 253777 65051
rect 253811 65023 253839 65051
rect 253625 64961 253653 64989
rect 253687 64961 253715 64989
rect 253749 64961 253777 64989
rect 253811 64961 253839 64989
rect 253625 56147 253653 56175
rect 253687 56147 253715 56175
rect 253749 56147 253777 56175
rect 253811 56147 253839 56175
rect 253625 56085 253653 56113
rect 253687 56085 253715 56113
rect 253749 56085 253777 56113
rect 253811 56085 253839 56113
rect 253625 56023 253653 56051
rect 253687 56023 253715 56051
rect 253749 56023 253777 56051
rect 253811 56023 253839 56051
rect 253625 55961 253653 55989
rect 253687 55961 253715 55989
rect 253749 55961 253777 55989
rect 253811 55961 253839 55989
rect 253625 47147 253653 47175
rect 253687 47147 253715 47175
rect 253749 47147 253777 47175
rect 253811 47147 253839 47175
rect 253625 47085 253653 47113
rect 253687 47085 253715 47113
rect 253749 47085 253777 47113
rect 253811 47085 253839 47113
rect 253625 47023 253653 47051
rect 253687 47023 253715 47051
rect 253749 47023 253777 47051
rect 253811 47023 253839 47051
rect 253625 46961 253653 46989
rect 253687 46961 253715 46989
rect 253749 46961 253777 46989
rect 253811 46961 253839 46989
rect 253625 38147 253653 38175
rect 253687 38147 253715 38175
rect 253749 38147 253777 38175
rect 253811 38147 253839 38175
rect 253625 38085 253653 38113
rect 253687 38085 253715 38113
rect 253749 38085 253777 38113
rect 253811 38085 253839 38113
rect 253625 38023 253653 38051
rect 253687 38023 253715 38051
rect 253749 38023 253777 38051
rect 253811 38023 253839 38051
rect 253625 37961 253653 37989
rect 253687 37961 253715 37989
rect 253749 37961 253777 37989
rect 253811 37961 253839 37989
rect 253625 29147 253653 29175
rect 253687 29147 253715 29175
rect 253749 29147 253777 29175
rect 253811 29147 253839 29175
rect 253625 29085 253653 29113
rect 253687 29085 253715 29113
rect 253749 29085 253777 29113
rect 253811 29085 253839 29113
rect 253625 29023 253653 29051
rect 253687 29023 253715 29051
rect 253749 29023 253777 29051
rect 253811 29023 253839 29051
rect 253625 28961 253653 28989
rect 253687 28961 253715 28989
rect 253749 28961 253777 28989
rect 253811 28961 253839 28989
rect 253625 20147 253653 20175
rect 253687 20147 253715 20175
rect 253749 20147 253777 20175
rect 253811 20147 253839 20175
rect 253625 20085 253653 20113
rect 253687 20085 253715 20113
rect 253749 20085 253777 20113
rect 253811 20085 253839 20113
rect 253625 20023 253653 20051
rect 253687 20023 253715 20051
rect 253749 20023 253777 20051
rect 253811 20023 253839 20051
rect 253625 19961 253653 19989
rect 253687 19961 253715 19989
rect 253749 19961 253777 19989
rect 253811 19961 253839 19989
rect 253625 11147 253653 11175
rect 253687 11147 253715 11175
rect 253749 11147 253777 11175
rect 253811 11147 253839 11175
rect 253625 11085 253653 11113
rect 253687 11085 253715 11113
rect 253749 11085 253777 11113
rect 253811 11085 253839 11113
rect 253625 11023 253653 11051
rect 253687 11023 253715 11051
rect 253749 11023 253777 11051
rect 253811 11023 253839 11051
rect 253625 10961 253653 10989
rect 253687 10961 253715 10989
rect 253749 10961 253777 10989
rect 253811 10961 253839 10989
rect 253625 2147 253653 2175
rect 253687 2147 253715 2175
rect 253749 2147 253777 2175
rect 253811 2147 253839 2175
rect 253625 2085 253653 2113
rect 253687 2085 253715 2113
rect 253749 2085 253777 2113
rect 253811 2085 253839 2113
rect 253625 2023 253653 2051
rect 253687 2023 253715 2051
rect 253749 2023 253777 2051
rect 253811 2023 253839 2051
rect 253625 1961 253653 1989
rect 253687 1961 253715 1989
rect 253749 1961 253777 1989
rect 253811 1961 253839 1989
rect 253625 -108 253653 -80
rect 253687 -108 253715 -80
rect 253749 -108 253777 -80
rect 253811 -108 253839 -80
rect 253625 -170 253653 -142
rect 253687 -170 253715 -142
rect 253749 -170 253777 -142
rect 253811 -170 253839 -142
rect 253625 -232 253653 -204
rect 253687 -232 253715 -204
rect 253749 -232 253777 -204
rect 253811 -232 253839 -204
rect 253625 -294 253653 -266
rect 253687 -294 253715 -266
rect 253749 -294 253777 -266
rect 253811 -294 253839 -266
rect 255485 299058 255513 299086
rect 255547 299058 255575 299086
rect 255609 299058 255637 299086
rect 255671 299058 255699 299086
rect 255485 298996 255513 299024
rect 255547 298996 255575 299024
rect 255609 298996 255637 299024
rect 255671 298996 255699 299024
rect 255485 298934 255513 298962
rect 255547 298934 255575 298962
rect 255609 298934 255637 298962
rect 255671 298934 255699 298962
rect 255485 298872 255513 298900
rect 255547 298872 255575 298900
rect 255609 298872 255637 298900
rect 255671 298872 255699 298900
rect 255485 293147 255513 293175
rect 255547 293147 255575 293175
rect 255609 293147 255637 293175
rect 255671 293147 255699 293175
rect 255485 293085 255513 293113
rect 255547 293085 255575 293113
rect 255609 293085 255637 293113
rect 255671 293085 255699 293113
rect 255485 293023 255513 293051
rect 255547 293023 255575 293051
rect 255609 293023 255637 293051
rect 255671 293023 255699 293051
rect 255485 292961 255513 292989
rect 255547 292961 255575 292989
rect 255609 292961 255637 292989
rect 255671 292961 255699 292989
rect 255485 284147 255513 284175
rect 255547 284147 255575 284175
rect 255609 284147 255637 284175
rect 255671 284147 255699 284175
rect 255485 284085 255513 284113
rect 255547 284085 255575 284113
rect 255609 284085 255637 284113
rect 255671 284085 255699 284113
rect 255485 284023 255513 284051
rect 255547 284023 255575 284051
rect 255609 284023 255637 284051
rect 255671 284023 255699 284051
rect 255485 283961 255513 283989
rect 255547 283961 255575 283989
rect 255609 283961 255637 283989
rect 255671 283961 255699 283989
rect 255485 275147 255513 275175
rect 255547 275147 255575 275175
rect 255609 275147 255637 275175
rect 255671 275147 255699 275175
rect 255485 275085 255513 275113
rect 255547 275085 255575 275113
rect 255609 275085 255637 275113
rect 255671 275085 255699 275113
rect 255485 275023 255513 275051
rect 255547 275023 255575 275051
rect 255609 275023 255637 275051
rect 255671 275023 255699 275051
rect 255485 274961 255513 274989
rect 255547 274961 255575 274989
rect 255609 274961 255637 274989
rect 255671 274961 255699 274989
rect 255485 266147 255513 266175
rect 255547 266147 255575 266175
rect 255609 266147 255637 266175
rect 255671 266147 255699 266175
rect 255485 266085 255513 266113
rect 255547 266085 255575 266113
rect 255609 266085 255637 266113
rect 255671 266085 255699 266113
rect 255485 266023 255513 266051
rect 255547 266023 255575 266051
rect 255609 266023 255637 266051
rect 255671 266023 255699 266051
rect 255485 265961 255513 265989
rect 255547 265961 255575 265989
rect 255609 265961 255637 265989
rect 255671 265961 255699 265989
rect 255485 257147 255513 257175
rect 255547 257147 255575 257175
rect 255609 257147 255637 257175
rect 255671 257147 255699 257175
rect 255485 257085 255513 257113
rect 255547 257085 255575 257113
rect 255609 257085 255637 257113
rect 255671 257085 255699 257113
rect 255485 257023 255513 257051
rect 255547 257023 255575 257051
rect 255609 257023 255637 257051
rect 255671 257023 255699 257051
rect 255485 256961 255513 256989
rect 255547 256961 255575 256989
rect 255609 256961 255637 256989
rect 255671 256961 255699 256989
rect 255485 248147 255513 248175
rect 255547 248147 255575 248175
rect 255609 248147 255637 248175
rect 255671 248147 255699 248175
rect 255485 248085 255513 248113
rect 255547 248085 255575 248113
rect 255609 248085 255637 248113
rect 255671 248085 255699 248113
rect 255485 248023 255513 248051
rect 255547 248023 255575 248051
rect 255609 248023 255637 248051
rect 255671 248023 255699 248051
rect 255485 247961 255513 247989
rect 255547 247961 255575 247989
rect 255609 247961 255637 247989
rect 255671 247961 255699 247989
rect 255485 239147 255513 239175
rect 255547 239147 255575 239175
rect 255609 239147 255637 239175
rect 255671 239147 255699 239175
rect 255485 239085 255513 239113
rect 255547 239085 255575 239113
rect 255609 239085 255637 239113
rect 255671 239085 255699 239113
rect 255485 239023 255513 239051
rect 255547 239023 255575 239051
rect 255609 239023 255637 239051
rect 255671 239023 255699 239051
rect 255485 238961 255513 238989
rect 255547 238961 255575 238989
rect 255609 238961 255637 238989
rect 255671 238961 255699 238989
rect 255485 230147 255513 230175
rect 255547 230147 255575 230175
rect 255609 230147 255637 230175
rect 255671 230147 255699 230175
rect 255485 230085 255513 230113
rect 255547 230085 255575 230113
rect 255609 230085 255637 230113
rect 255671 230085 255699 230113
rect 255485 230023 255513 230051
rect 255547 230023 255575 230051
rect 255609 230023 255637 230051
rect 255671 230023 255699 230051
rect 255485 229961 255513 229989
rect 255547 229961 255575 229989
rect 255609 229961 255637 229989
rect 255671 229961 255699 229989
rect 255485 221147 255513 221175
rect 255547 221147 255575 221175
rect 255609 221147 255637 221175
rect 255671 221147 255699 221175
rect 255485 221085 255513 221113
rect 255547 221085 255575 221113
rect 255609 221085 255637 221113
rect 255671 221085 255699 221113
rect 255485 221023 255513 221051
rect 255547 221023 255575 221051
rect 255609 221023 255637 221051
rect 255671 221023 255699 221051
rect 255485 220961 255513 220989
rect 255547 220961 255575 220989
rect 255609 220961 255637 220989
rect 255671 220961 255699 220989
rect 255485 212147 255513 212175
rect 255547 212147 255575 212175
rect 255609 212147 255637 212175
rect 255671 212147 255699 212175
rect 255485 212085 255513 212113
rect 255547 212085 255575 212113
rect 255609 212085 255637 212113
rect 255671 212085 255699 212113
rect 255485 212023 255513 212051
rect 255547 212023 255575 212051
rect 255609 212023 255637 212051
rect 255671 212023 255699 212051
rect 255485 211961 255513 211989
rect 255547 211961 255575 211989
rect 255609 211961 255637 211989
rect 255671 211961 255699 211989
rect 255485 203147 255513 203175
rect 255547 203147 255575 203175
rect 255609 203147 255637 203175
rect 255671 203147 255699 203175
rect 255485 203085 255513 203113
rect 255547 203085 255575 203113
rect 255609 203085 255637 203113
rect 255671 203085 255699 203113
rect 255485 203023 255513 203051
rect 255547 203023 255575 203051
rect 255609 203023 255637 203051
rect 255671 203023 255699 203051
rect 255485 202961 255513 202989
rect 255547 202961 255575 202989
rect 255609 202961 255637 202989
rect 255671 202961 255699 202989
rect 255485 194147 255513 194175
rect 255547 194147 255575 194175
rect 255609 194147 255637 194175
rect 255671 194147 255699 194175
rect 255485 194085 255513 194113
rect 255547 194085 255575 194113
rect 255609 194085 255637 194113
rect 255671 194085 255699 194113
rect 255485 194023 255513 194051
rect 255547 194023 255575 194051
rect 255609 194023 255637 194051
rect 255671 194023 255699 194051
rect 255485 193961 255513 193989
rect 255547 193961 255575 193989
rect 255609 193961 255637 193989
rect 255671 193961 255699 193989
rect 255485 185147 255513 185175
rect 255547 185147 255575 185175
rect 255609 185147 255637 185175
rect 255671 185147 255699 185175
rect 255485 185085 255513 185113
rect 255547 185085 255575 185113
rect 255609 185085 255637 185113
rect 255671 185085 255699 185113
rect 255485 185023 255513 185051
rect 255547 185023 255575 185051
rect 255609 185023 255637 185051
rect 255671 185023 255699 185051
rect 255485 184961 255513 184989
rect 255547 184961 255575 184989
rect 255609 184961 255637 184989
rect 255671 184961 255699 184989
rect 255485 176147 255513 176175
rect 255547 176147 255575 176175
rect 255609 176147 255637 176175
rect 255671 176147 255699 176175
rect 255485 176085 255513 176113
rect 255547 176085 255575 176113
rect 255609 176085 255637 176113
rect 255671 176085 255699 176113
rect 255485 176023 255513 176051
rect 255547 176023 255575 176051
rect 255609 176023 255637 176051
rect 255671 176023 255699 176051
rect 255485 175961 255513 175989
rect 255547 175961 255575 175989
rect 255609 175961 255637 175989
rect 255671 175961 255699 175989
rect 255485 167147 255513 167175
rect 255547 167147 255575 167175
rect 255609 167147 255637 167175
rect 255671 167147 255699 167175
rect 255485 167085 255513 167113
rect 255547 167085 255575 167113
rect 255609 167085 255637 167113
rect 255671 167085 255699 167113
rect 255485 167023 255513 167051
rect 255547 167023 255575 167051
rect 255609 167023 255637 167051
rect 255671 167023 255699 167051
rect 255485 166961 255513 166989
rect 255547 166961 255575 166989
rect 255609 166961 255637 166989
rect 255671 166961 255699 166989
rect 255485 158147 255513 158175
rect 255547 158147 255575 158175
rect 255609 158147 255637 158175
rect 255671 158147 255699 158175
rect 255485 158085 255513 158113
rect 255547 158085 255575 158113
rect 255609 158085 255637 158113
rect 255671 158085 255699 158113
rect 255485 158023 255513 158051
rect 255547 158023 255575 158051
rect 255609 158023 255637 158051
rect 255671 158023 255699 158051
rect 255485 157961 255513 157989
rect 255547 157961 255575 157989
rect 255609 157961 255637 157989
rect 255671 157961 255699 157989
rect 255485 149147 255513 149175
rect 255547 149147 255575 149175
rect 255609 149147 255637 149175
rect 255671 149147 255699 149175
rect 255485 149085 255513 149113
rect 255547 149085 255575 149113
rect 255609 149085 255637 149113
rect 255671 149085 255699 149113
rect 255485 149023 255513 149051
rect 255547 149023 255575 149051
rect 255609 149023 255637 149051
rect 255671 149023 255699 149051
rect 255485 148961 255513 148989
rect 255547 148961 255575 148989
rect 255609 148961 255637 148989
rect 255671 148961 255699 148989
rect 255485 140147 255513 140175
rect 255547 140147 255575 140175
rect 255609 140147 255637 140175
rect 255671 140147 255699 140175
rect 255485 140085 255513 140113
rect 255547 140085 255575 140113
rect 255609 140085 255637 140113
rect 255671 140085 255699 140113
rect 255485 140023 255513 140051
rect 255547 140023 255575 140051
rect 255609 140023 255637 140051
rect 255671 140023 255699 140051
rect 255485 139961 255513 139989
rect 255547 139961 255575 139989
rect 255609 139961 255637 139989
rect 255671 139961 255699 139989
rect 255485 131147 255513 131175
rect 255547 131147 255575 131175
rect 255609 131147 255637 131175
rect 255671 131147 255699 131175
rect 255485 131085 255513 131113
rect 255547 131085 255575 131113
rect 255609 131085 255637 131113
rect 255671 131085 255699 131113
rect 255485 131023 255513 131051
rect 255547 131023 255575 131051
rect 255609 131023 255637 131051
rect 255671 131023 255699 131051
rect 255485 130961 255513 130989
rect 255547 130961 255575 130989
rect 255609 130961 255637 130989
rect 255671 130961 255699 130989
rect 255485 122147 255513 122175
rect 255547 122147 255575 122175
rect 255609 122147 255637 122175
rect 255671 122147 255699 122175
rect 255485 122085 255513 122113
rect 255547 122085 255575 122113
rect 255609 122085 255637 122113
rect 255671 122085 255699 122113
rect 255485 122023 255513 122051
rect 255547 122023 255575 122051
rect 255609 122023 255637 122051
rect 255671 122023 255699 122051
rect 255485 121961 255513 121989
rect 255547 121961 255575 121989
rect 255609 121961 255637 121989
rect 255671 121961 255699 121989
rect 255485 113147 255513 113175
rect 255547 113147 255575 113175
rect 255609 113147 255637 113175
rect 255671 113147 255699 113175
rect 255485 113085 255513 113113
rect 255547 113085 255575 113113
rect 255609 113085 255637 113113
rect 255671 113085 255699 113113
rect 255485 113023 255513 113051
rect 255547 113023 255575 113051
rect 255609 113023 255637 113051
rect 255671 113023 255699 113051
rect 255485 112961 255513 112989
rect 255547 112961 255575 112989
rect 255609 112961 255637 112989
rect 255671 112961 255699 112989
rect 255485 104147 255513 104175
rect 255547 104147 255575 104175
rect 255609 104147 255637 104175
rect 255671 104147 255699 104175
rect 255485 104085 255513 104113
rect 255547 104085 255575 104113
rect 255609 104085 255637 104113
rect 255671 104085 255699 104113
rect 255485 104023 255513 104051
rect 255547 104023 255575 104051
rect 255609 104023 255637 104051
rect 255671 104023 255699 104051
rect 255485 103961 255513 103989
rect 255547 103961 255575 103989
rect 255609 103961 255637 103989
rect 255671 103961 255699 103989
rect 255485 95147 255513 95175
rect 255547 95147 255575 95175
rect 255609 95147 255637 95175
rect 255671 95147 255699 95175
rect 255485 95085 255513 95113
rect 255547 95085 255575 95113
rect 255609 95085 255637 95113
rect 255671 95085 255699 95113
rect 255485 95023 255513 95051
rect 255547 95023 255575 95051
rect 255609 95023 255637 95051
rect 255671 95023 255699 95051
rect 255485 94961 255513 94989
rect 255547 94961 255575 94989
rect 255609 94961 255637 94989
rect 255671 94961 255699 94989
rect 255485 86147 255513 86175
rect 255547 86147 255575 86175
rect 255609 86147 255637 86175
rect 255671 86147 255699 86175
rect 255485 86085 255513 86113
rect 255547 86085 255575 86113
rect 255609 86085 255637 86113
rect 255671 86085 255699 86113
rect 255485 86023 255513 86051
rect 255547 86023 255575 86051
rect 255609 86023 255637 86051
rect 255671 86023 255699 86051
rect 255485 85961 255513 85989
rect 255547 85961 255575 85989
rect 255609 85961 255637 85989
rect 255671 85961 255699 85989
rect 255485 77147 255513 77175
rect 255547 77147 255575 77175
rect 255609 77147 255637 77175
rect 255671 77147 255699 77175
rect 255485 77085 255513 77113
rect 255547 77085 255575 77113
rect 255609 77085 255637 77113
rect 255671 77085 255699 77113
rect 255485 77023 255513 77051
rect 255547 77023 255575 77051
rect 255609 77023 255637 77051
rect 255671 77023 255699 77051
rect 255485 76961 255513 76989
rect 255547 76961 255575 76989
rect 255609 76961 255637 76989
rect 255671 76961 255699 76989
rect 255485 68147 255513 68175
rect 255547 68147 255575 68175
rect 255609 68147 255637 68175
rect 255671 68147 255699 68175
rect 255485 68085 255513 68113
rect 255547 68085 255575 68113
rect 255609 68085 255637 68113
rect 255671 68085 255699 68113
rect 255485 68023 255513 68051
rect 255547 68023 255575 68051
rect 255609 68023 255637 68051
rect 255671 68023 255699 68051
rect 255485 67961 255513 67989
rect 255547 67961 255575 67989
rect 255609 67961 255637 67989
rect 255671 67961 255699 67989
rect 255485 59147 255513 59175
rect 255547 59147 255575 59175
rect 255609 59147 255637 59175
rect 255671 59147 255699 59175
rect 255485 59085 255513 59113
rect 255547 59085 255575 59113
rect 255609 59085 255637 59113
rect 255671 59085 255699 59113
rect 255485 59023 255513 59051
rect 255547 59023 255575 59051
rect 255609 59023 255637 59051
rect 255671 59023 255699 59051
rect 255485 58961 255513 58989
rect 255547 58961 255575 58989
rect 255609 58961 255637 58989
rect 255671 58961 255699 58989
rect 255485 50147 255513 50175
rect 255547 50147 255575 50175
rect 255609 50147 255637 50175
rect 255671 50147 255699 50175
rect 255485 50085 255513 50113
rect 255547 50085 255575 50113
rect 255609 50085 255637 50113
rect 255671 50085 255699 50113
rect 255485 50023 255513 50051
rect 255547 50023 255575 50051
rect 255609 50023 255637 50051
rect 255671 50023 255699 50051
rect 255485 49961 255513 49989
rect 255547 49961 255575 49989
rect 255609 49961 255637 49989
rect 255671 49961 255699 49989
rect 255485 41147 255513 41175
rect 255547 41147 255575 41175
rect 255609 41147 255637 41175
rect 255671 41147 255699 41175
rect 255485 41085 255513 41113
rect 255547 41085 255575 41113
rect 255609 41085 255637 41113
rect 255671 41085 255699 41113
rect 255485 41023 255513 41051
rect 255547 41023 255575 41051
rect 255609 41023 255637 41051
rect 255671 41023 255699 41051
rect 255485 40961 255513 40989
rect 255547 40961 255575 40989
rect 255609 40961 255637 40989
rect 255671 40961 255699 40989
rect 255485 32147 255513 32175
rect 255547 32147 255575 32175
rect 255609 32147 255637 32175
rect 255671 32147 255699 32175
rect 255485 32085 255513 32113
rect 255547 32085 255575 32113
rect 255609 32085 255637 32113
rect 255671 32085 255699 32113
rect 255485 32023 255513 32051
rect 255547 32023 255575 32051
rect 255609 32023 255637 32051
rect 255671 32023 255699 32051
rect 255485 31961 255513 31989
rect 255547 31961 255575 31989
rect 255609 31961 255637 31989
rect 255671 31961 255699 31989
rect 255485 23147 255513 23175
rect 255547 23147 255575 23175
rect 255609 23147 255637 23175
rect 255671 23147 255699 23175
rect 255485 23085 255513 23113
rect 255547 23085 255575 23113
rect 255609 23085 255637 23113
rect 255671 23085 255699 23113
rect 255485 23023 255513 23051
rect 255547 23023 255575 23051
rect 255609 23023 255637 23051
rect 255671 23023 255699 23051
rect 255485 22961 255513 22989
rect 255547 22961 255575 22989
rect 255609 22961 255637 22989
rect 255671 22961 255699 22989
rect 255485 14147 255513 14175
rect 255547 14147 255575 14175
rect 255609 14147 255637 14175
rect 255671 14147 255699 14175
rect 255485 14085 255513 14113
rect 255547 14085 255575 14113
rect 255609 14085 255637 14113
rect 255671 14085 255699 14113
rect 255485 14023 255513 14051
rect 255547 14023 255575 14051
rect 255609 14023 255637 14051
rect 255671 14023 255699 14051
rect 255485 13961 255513 13989
rect 255547 13961 255575 13989
rect 255609 13961 255637 13989
rect 255671 13961 255699 13989
rect 255485 5147 255513 5175
rect 255547 5147 255575 5175
rect 255609 5147 255637 5175
rect 255671 5147 255699 5175
rect 255485 5085 255513 5113
rect 255547 5085 255575 5113
rect 255609 5085 255637 5113
rect 255671 5085 255699 5113
rect 255485 5023 255513 5051
rect 255547 5023 255575 5051
rect 255609 5023 255637 5051
rect 255671 5023 255699 5051
rect 255485 4961 255513 4989
rect 255547 4961 255575 4989
rect 255609 4961 255637 4989
rect 255671 4961 255699 4989
rect 255485 -588 255513 -560
rect 255547 -588 255575 -560
rect 255609 -588 255637 -560
rect 255671 -588 255699 -560
rect 255485 -650 255513 -622
rect 255547 -650 255575 -622
rect 255609 -650 255637 -622
rect 255671 -650 255699 -622
rect 255485 -712 255513 -684
rect 255547 -712 255575 -684
rect 255609 -712 255637 -684
rect 255671 -712 255699 -684
rect 255485 -774 255513 -746
rect 255547 -774 255575 -746
rect 255609 -774 255637 -746
rect 255671 -774 255699 -746
rect 262625 298578 262653 298606
rect 262687 298578 262715 298606
rect 262749 298578 262777 298606
rect 262811 298578 262839 298606
rect 262625 298516 262653 298544
rect 262687 298516 262715 298544
rect 262749 298516 262777 298544
rect 262811 298516 262839 298544
rect 262625 298454 262653 298482
rect 262687 298454 262715 298482
rect 262749 298454 262777 298482
rect 262811 298454 262839 298482
rect 262625 298392 262653 298420
rect 262687 298392 262715 298420
rect 262749 298392 262777 298420
rect 262811 298392 262839 298420
rect 262625 290147 262653 290175
rect 262687 290147 262715 290175
rect 262749 290147 262777 290175
rect 262811 290147 262839 290175
rect 262625 290085 262653 290113
rect 262687 290085 262715 290113
rect 262749 290085 262777 290113
rect 262811 290085 262839 290113
rect 262625 290023 262653 290051
rect 262687 290023 262715 290051
rect 262749 290023 262777 290051
rect 262811 290023 262839 290051
rect 262625 289961 262653 289989
rect 262687 289961 262715 289989
rect 262749 289961 262777 289989
rect 262811 289961 262839 289989
rect 262625 281147 262653 281175
rect 262687 281147 262715 281175
rect 262749 281147 262777 281175
rect 262811 281147 262839 281175
rect 262625 281085 262653 281113
rect 262687 281085 262715 281113
rect 262749 281085 262777 281113
rect 262811 281085 262839 281113
rect 262625 281023 262653 281051
rect 262687 281023 262715 281051
rect 262749 281023 262777 281051
rect 262811 281023 262839 281051
rect 262625 280961 262653 280989
rect 262687 280961 262715 280989
rect 262749 280961 262777 280989
rect 262811 280961 262839 280989
rect 262625 272147 262653 272175
rect 262687 272147 262715 272175
rect 262749 272147 262777 272175
rect 262811 272147 262839 272175
rect 262625 272085 262653 272113
rect 262687 272085 262715 272113
rect 262749 272085 262777 272113
rect 262811 272085 262839 272113
rect 262625 272023 262653 272051
rect 262687 272023 262715 272051
rect 262749 272023 262777 272051
rect 262811 272023 262839 272051
rect 262625 271961 262653 271989
rect 262687 271961 262715 271989
rect 262749 271961 262777 271989
rect 262811 271961 262839 271989
rect 262625 263147 262653 263175
rect 262687 263147 262715 263175
rect 262749 263147 262777 263175
rect 262811 263147 262839 263175
rect 262625 263085 262653 263113
rect 262687 263085 262715 263113
rect 262749 263085 262777 263113
rect 262811 263085 262839 263113
rect 262625 263023 262653 263051
rect 262687 263023 262715 263051
rect 262749 263023 262777 263051
rect 262811 263023 262839 263051
rect 262625 262961 262653 262989
rect 262687 262961 262715 262989
rect 262749 262961 262777 262989
rect 262811 262961 262839 262989
rect 262625 254147 262653 254175
rect 262687 254147 262715 254175
rect 262749 254147 262777 254175
rect 262811 254147 262839 254175
rect 262625 254085 262653 254113
rect 262687 254085 262715 254113
rect 262749 254085 262777 254113
rect 262811 254085 262839 254113
rect 262625 254023 262653 254051
rect 262687 254023 262715 254051
rect 262749 254023 262777 254051
rect 262811 254023 262839 254051
rect 262625 253961 262653 253989
rect 262687 253961 262715 253989
rect 262749 253961 262777 253989
rect 262811 253961 262839 253989
rect 262625 245147 262653 245175
rect 262687 245147 262715 245175
rect 262749 245147 262777 245175
rect 262811 245147 262839 245175
rect 262625 245085 262653 245113
rect 262687 245085 262715 245113
rect 262749 245085 262777 245113
rect 262811 245085 262839 245113
rect 262625 245023 262653 245051
rect 262687 245023 262715 245051
rect 262749 245023 262777 245051
rect 262811 245023 262839 245051
rect 262625 244961 262653 244989
rect 262687 244961 262715 244989
rect 262749 244961 262777 244989
rect 262811 244961 262839 244989
rect 262625 236147 262653 236175
rect 262687 236147 262715 236175
rect 262749 236147 262777 236175
rect 262811 236147 262839 236175
rect 262625 236085 262653 236113
rect 262687 236085 262715 236113
rect 262749 236085 262777 236113
rect 262811 236085 262839 236113
rect 262625 236023 262653 236051
rect 262687 236023 262715 236051
rect 262749 236023 262777 236051
rect 262811 236023 262839 236051
rect 262625 235961 262653 235989
rect 262687 235961 262715 235989
rect 262749 235961 262777 235989
rect 262811 235961 262839 235989
rect 262625 227147 262653 227175
rect 262687 227147 262715 227175
rect 262749 227147 262777 227175
rect 262811 227147 262839 227175
rect 262625 227085 262653 227113
rect 262687 227085 262715 227113
rect 262749 227085 262777 227113
rect 262811 227085 262839 227113
rect 262625 227023 262653 227051
rect 262687 227023 262715 227051
rect 262749 227023 262777 227051
rect 262811 227023 262839 227051
rect 262625 226961 262653 226989
rect 262687 226961 262715 226989
rect 262749 226961 262777 226989
rect 262811 226961 262839 226989
rect 262625 218147 262653 218175
rect 262687 218147 262715 218175
rect 262749 218147 262777 218175
rect 262811 218147 262839 218175
rect 262625 218085 262653 218113
rect 262687 218085 262715 218113
rect 262749 218085 262777 218113
rect 262811 218085 262839 218113
rect 262625 218023 262653 218051
rect 262687 218023 262715 218051
rect 262749 218023 262777 218051
rect 262811 218023 262839 218051
rect 262625 217961 262653 217989
rect 262687 217961 262715 217989
rect 262749 217961 262777 217989
rect 262811 217961 262839 217989
rect 262625 209147 262653 209175
rect 262687 209147 262715 209175
rect 262749 209147 262777 209175
rect 262811 209147 262839 209175
rect 262625 209085 262653 209113
rect 262687 209085 262715 209113
rect 262749 209085 262777 209113
rect 262811 209085 262839 209113
rect 262625 209023 262653 209051
rect 262687 209023 262715 209051
rect 262749 209023 262777 209051
rect 262811 209023 262839 209051
rect 262625 208961 262653 208989
rect 262687 208961 262715 208989
rect 262749 208961 262777 208989
rect 262811 208961 262839 208989
rect 262625 200147 262653 200175
rect 262687 200147 262715 200175
rect 262749 200147 262777 200175
rect 262811 200147 262839 200175
rect 262625 200085 262653 200113
rect 262687 200085 262715 200113
rect 262749 200085 262777 200113
rect 262811 200085 262839 200113
rect 262625 200023 262653 200051
rect 262687 200023 262715 200051
rect 262749 200023 262777 200051
rect 262811 200023 262839 200051
rect 262625 199961 262653 199989
rect 262687 199961 262715 199989
rect 262749 199961 262777 199989
rect 262811 199961 262839 199989
rect 262625 191147 262653 191175
rect 262687 191147 262715 191175
rect 262749 191147 262777 191175
rect 262811 191147 262839 191175
rect 262625 191085 262653 191113
rect 262687 191085 262715 191113
rect 262749 191085 262777 191113
rect 262811 191085 262839 191113
rect 262625 191023 262653 191051
rect 262687 191023 262715 191051
rect 262749 191023 262777 191051
rect 262811 191023 262839 191051
rect 262625 190961 262653 190989
rect 262687 190961 262715 190989
rect 262749 190961 262777 190989
rect 262811 190961 262839 190989
rect 262625 182147 262653 182175
rect 262687 182147 262715 182175
rect 262749 182147 262777 182175
rect 262811 182147 262839 182175
rect 262625 182085 262653 182113
rect 262687 182085 262715 182113
rect 262749 182085 262777 182113
rect 262811 182085 262839 182113
rect 262625 182023 262653 182051
rect 262687 182023 262715 182051
rect 262749 182023 262777 182051
rect 262811 182023 262839 182051
rect 262625 181961 262653 181989
rect 262687 181961 262715 181989
rect 262749 181961 262777 181989
rect 262811 181961 262839 181989
rect 262625 173147 262653 173175
rect 262687 173147 262715 173175
rect 262749 173147 262777 173175
rect 262811 173147 262839 173175
rect 262625 173085 262653 173113
rect 262687 173085 262715 173113
rect 262749 173085 262777 173113
rect 262811 173085 262839 173113
rect 262625 173023 262653 173051
rect 262687 173023 262715 173051
rect 262749 173023 262777 173051
rect 262811 173023 262839 173051
rect 262625 172961 262653 172989
rect 262687 172961 262715 172989
rect 262749 172961 262777 172989
rect 262811 172961 262839 172989
rect 262625 164147 262653 164175
rect 262687 164147 262715 164175
rect 262749 164147 262777 164175
rect 262811 164147 262839 164175
rect 262625 164085 262653 164113
rect 262687 164085 262715 164113
rect 262749 164085 262777 164113
rect 262811 164085 262839 164113
rect 262625 164023 262653 164051
rect 262687 164023 262715 164051
rect 262749 164023 262777 164051
rect 262811 164023 262839 164051
rect 262625 163961 262653 163989
rect 262687 163961 262715 163989
rect 262749 163961 262777 163989
rect 262811 163961 262839 163989
rect 262625 155147 262653 155175
rect 262687 155147 262715 155175
rect 262749 155147 262777 155175
rect 262811 155147 262839 155175
rect 262625 155085 262653 155113
rect 262687 155085 262715 155113
rect 262749 155085 262777 155113
rect 262811 155085 262839 155113
rect 262625 155023 262653 155051
rect 262687 155023 262715 155051
rect 262749 155023 262777 155051
rect 262811 155023 262839 155051
rect 262625 154961 262653 154989
rect 262687 154961 262715 154989
rect 262749 154961 262777 154989
rect 262811 154961 262839 154989
rect 262625 146147 262653 146175
rect 262687 146147 262715 146175
rect 262749 146147 262777 146175
rect 262811 146147 262839 146175
rect 262625 146085 262653 146113
rect 262687 146085 262715 146113
rect 262749 146085 262777 146113
rect 262811 146085 262839 146113
rect 262625 146023 262653 146051
rect 262687 146023 262715 146051
rect 262749 146023 262777 146051
rect 262811 146023 262839 146051
rect 262625 145961 262653 145989
rect 262687 145961 262715 145989
rect 262749 145961 262777 145989
rect 262811 145961 262839 145989
rect 262625 137147 262653 137175
rect 262687 137147 262715 137175
rect 262749 137147 262777 137175
rect 262811 137147 262839 137175
rect 262625 137085 262653 137113
rect 262687 137085 262715 137113
rect 262749 137085 262777 137113
rect 262811 137085 262839 137113
rect 262625 137023 262653 137051
rect 262687 137023 262715 137051
rect 262749 137023 262777 137051
rect 262811 137023 262839 137051
rect 262625 136961 262653 136989
rect 262687 136961 262715 136989
rect 262749 136961 262777 136989
rect 262811 136961 262839 136989
rect 262625 128147 262653 128175
rect 262687 128147 262715 128175
rect 262749 128147 262777 128175
rect 262811 128147 262839 128175
rect 262625 128085 262653 128113
rect 262687 128085 262715 128113
rect 262749 128085 262777 128113
rect 262811 128085 262839 128113
rect 262625 128023 262653 128051
rect 262687 128023 262715 128051
rect 262749 128023 262777 128051
rect 262811 128023 262839 128051
rect 262625 127961 262653 127989
rect 262687 127961 262715 127989
rect 262749 127961 262777 127989
rect 262811 127961 262839 127989
rect 262625 119147 262653 119175
rect 262687 119147 262715 119175
rect 262749 119147 262777 119175
rect 262811 119147 262839 119175
rect 262625 119085 262653 119113
rect 262687 119085 262715 119113
rect 262749 119085 262777 119113
rect 262811 119085 262839 119113
rect 262625 119023 262653 119051
rect 262687 119023 262715 119051
rect 262749 119023 262777 119051
rect 262811 119023 262839 119051
rect 262625 118961 262653 118989
rect 262687 118961 262715 118989
rect 262749 118961 262777 118989
rect 262811 118961 262839 118989
rect 262625 110147 262653 110175
rect 262687 110147 262715 110175
rect 262749 110147 262777 110175
rect 262811 110147 262839 110175
rect 262625 110085 262653 110113
rect 262687 110085 262715 110113
rect 262749 110085 262777 110113
rect 262811 110085 262839 110113
rect 262625 110023 262653 110051
rect 262687 110023 262715 110051
rect 262749 110023 262777 110051
rect 262811 110023 262839 110051
rect 262625 109961 262653 109989
rect 262687 109961 262715 109989
rect 262749 109961 262777 109989
rect 262811 109961 262839 109989
rect 262625 101147 262653 101175
rect 262687 101147 262715 101175
rect 262749 101147 262777 101175
rect 262811 101147 262839 101175
rect 262625 101085 262653 101113
rect 262687 101085 262715 101113
rect 262749 101085 262777 101113
rect 262811 101085 262839 101113
rect 262625 101023 262653 101051
rect 262687 101023 262715 101051
rect 262749 101023 262777 101051
rect 262811 101023 262839 101051
rect 262625 100961 262653 100989
rect 262687 100961 262715 100989
rect 262749 100961 262777 100989
rect 262811 100961 262839 100989
rect 262625 92147 262653 92175
rect 262687 92147 262715 92175
rect 262749 92147 262777 92175
rect 262811 92147 262839 92175
rect 262625 92085 262653 92113
rect 262687 92085 262715 92113
rect 262749 92085 262777 92113
rect 262811 92085 262839 92113
rect 262625 92023 262653 92051
rect 262687 92023 262715 92051
rect 262749 92023 262777 92051
rect 262811 92023 262839 92051
rect 262625 91961 262653 91989
rect 262687 91961 262715 91989
rect 262749 91961 262777 91989
rect 262811 91961 262839 91989
rect 262625 83147 262653 83175
rect 262687 83147 262715 83175
rect 262749 83147 262777 83175
rect 262811 83147 262839 83175
rect 262625 83085 262653 83113
rect 262687 83085 262715 83113
rect 262749 83085 262777 83113
rect 262811 83085 262839 83113
rect 262625 83023 262653 83051
rect 262687 83023 262715 83051
rect 262749 83023 262777 83051
rect 262811 83023 262839 83051
rect 262625 82961 262653 82989
rect 262687 82961 262715 82989
rect 262749 82961 262777 82989
rect 262811 82961 262839 82989
rect 262625 74147 262653 74175
rect 262687 74147 262715 74175
rect 262749 74147 262777 74175
rect 262811 74147 262839 74175
rect 262625 74085 262653 74113
rect 262687 74085 262715 74113
rect 262749 74085 262777 74113
rect 262811 74085 262839 74113
rect 262625 74023 262653 74051
rect 262687 74023 262715 74051
rect 262749 74023 262777 74051
rect 262811 74023 262839 74051
rect 262625 73961 262653 73989
rect 262687 73961 262715 73989
rect 262749 73961 262777 73989
rect 262811 73961 262839 73989
rect 262625 65147 262653 65175
rect 262687 65147 262715 65175
rect 262749 65147 262777 65175
rect 262811 65147 262839 65175
rect 262625 65085 262653 65113
rect 262687 65085 262715 65113
rect 262749 65085 262777 65113
rect 262811 65085 262839 65113
rect 262625 65023 262653 65051
rect 262687 65023 262715 65051
rect 262749 65023 262777 65051
rect 262811 65023 262839 65051
rect 262625 64961 262653 64989
rect 262687 64961 262715 64989
rect 262749 64961 262777 64989
rect 262811 64961 262839 64989
rect 262625 56147 262653 56175
rect 262687 56147 262715 56175
rect 262749 56147 262777 56175
rect 262811 56147 262839 56175
rect 262625 56085 262653 56113
rect 262687 56085 262715 56113
rect 262749 56085 262777 56113
rect 262811 56085 262839 56113
rect 262625 56023 262653 56051
rect 262687 56023 262715 56051
rect 262749 56023 262777 56051
rect 262811 56023 262839 56051
rect 262625 55961 262653 55989
rect 262687 55961 262715 55989
rect 262749 55961 262777 55989
rect 262811 55961 262839 55989
rect 262625 47147 262653 47175
rect 262687 47147 262715 47175
rect 262749 47147 262777 47175
rect 262811 47147 262839 47175
rect 262625 47085 262653 47113
rect 262687 47085 262715 47113
rect 262749 47085 262777 47113
rect 262811 47085 262839 47113
rect 262625 47023 262653 47051
rect 262687 47023 262715 47051
rect 262749 47023 262777 47051
rect 262811 47023 262839 47051
rect 262625 46961 262653 46989
rect 262687 46961 262715 46989
rect 262749 46961 262777 46989
rect 262811 46961 262839 46989
rect 262625 38147 262653 38175
rect 262687 38147 262715 38175
rect 262749 38147 262777 38175
rect 262811 38147 262839 38175
rect 262625 38085 262653 38113
rect 262687 38085 262715 38113
rect 262749 38085 262777 38113
rect 262811 38085 262839 38113
rect 262625 38023 262653 38051
rect 262687 38023 262715 38051
rect 262749 38023 262777 38051
rect 262811 38023 262839 38051
rect 262625 37961 262653 37989
rect 262687 37961 262715 37989
rect 262749 37961 262777 37989
rect 262811 37961 262839 37989
rect 262625 29147 262653 29175
rect 262687 29147 262715 29175
rect 262749 29147 262777 29175
rect 262811 29147 262839 29175
rect 262625 29085 262653 29113
rect 262687 29085 262715 29113
rect 262749 29085 262777 29113
rect 262811 29085 262839 29113
rect 262625 29023 262653 29051
rect 262687 29023 262715 29051
rect 262749 29023 262777 29051
rect 262811 29023 262839 29051
rect 262625 28961 262653 28989
rect 262687 28961 262715 28989
rect 262749 28961 262777 28989
rect 262811 28961 262839 28989
rect 262625 20147 262653 20175
rect 262687 20147 262715 20175
rect 262749 20147 262777 20175
rect 262811 20147 262839 20175
rect 262625 20085 262653 20113
rect 262687 20085 262715 20113
rect 262749 20085 262777 20113
rect 262811 20085 262839 20113
rect 262625 20023 262653 20051
rect 262687 20023 262715 20051
rect 262749 20023 262777 20051
rect 262811 20023 262839 20051
rect 262625 19961 262653 19989
rect 262687 19961 262715 19989
rect 262749 19961 262777 19989
rect 262811 19961 262839 19989
rect 262625 11147 262653 11175
rect 262687 11147 262715 11175
rect 262749 11147 262777 11175
rect 262811 11147 262839 11175
rect 262625 11085 262653 11113
rect 262687 11085 262715 11113
rect 262749 11085 262777 11113
rect 262811 11085 262839 11113
rect 262625 11023 262653 11051
rect 262687 11023 262715 11051
rect 262749 11023 262777 11051
rect 262811 11023 262839 11051
rect 262625 10961 262653 10989
rect 262687 10961 262715 10989
rect 262749 10961 262777 10989
rect 262811 10961 262839 10989
rect 262625 2147 262653 2175
rect 262687 2147 262715 2175
rect 262749 2147 262777 2175
rect 262811 2147 262839 2175
rect 262625 2085 262653 2113
rect 262687 2085 262715 2113
rect 262749 2085 262777 2113
rect 262811 2085 262839 2113
rect 262625 2023 262653 2051
rect 262687 2023 262715 2051
rect 262749 2023 262777 2051
rect 262811 2023 262839 2051
rect 262625 1961 262653 1989
rect 262687 1961 262715 1989
rect 262749 1961 262777 1989
rect 262811 1961 262839 1989
rect 262625 -108 262653 -80
rect 262687 -108 262715 -80
rect 262749 -108 262777 -80
rect 262811 -108 262839 -80
rect 262625 -170 262653 -142
rect 262687 -170 262715 -142
rect 262749 -170 262777 -142
rect 262811 -170 262839 -142
rect 262625 -232 262653 -204
rect 262687 -232 262715 -204
rect 262749 -232 262777 -204
rect 262811 -232 262839 -204
rect 262625 -294 262653 -266
rect 262687 -294 262715 -266
rect 262749 -294 262777 -266
rect 262811 -294 262839 -266
rect 264485 299058 264513 299086
rect 264547 299058 264575 299086
rect 264609 299058 264637 299086
rect 264671 299058 264699 299086
rect 264485 298996 264513 299024
rect 264547 298996 264575 299024
rect 264609 298996 264637 299024
rect 264671 298996 264699 299024
rect 264485 298934 264513 298962
rect 264547 298934 264575 298962
rect 264609 298934 264637 298962
rect 264671 298934 264699 298962
rect 264485 298872 264513 298900
rect 264547 298872 264575 298900
rect 264609 298872 264637 298900
rect 264671 298872 264699 298900
rect 264485 293147 264513 293175
rect 264547 293147 264575 293175
rect 264609 293147 264637 293175
rect 264671 293147 264699 293175
rect 264485 293085 264513 293113
rect 264547 293085 264575 293113
rect 264609 293085 264637 293113
rect 264671 293085 264699 293113
rect 264485 293023 264513 293051
rect 264547 293023 264575 293051
rect 264609 293023 264637 293051
rect 264671 293023 264699 293051
rect 264485 292961 264513 292989
rect 264547 292961 264575 292989
rect 264609 292961 264637 292989
rect 264671 292961 264699 292989
rect 264485 284147 264513 284175
rect 264547 284147 264575 284175
rect 264609 284147 264637 284175
rect 264671 284147 264699 284175
rect 264485 284085 264513 284113
rect 264547 284085 264575 284113
rect 264609 284085 264637 284113
rect 264671 284085 264699 284113
rect 264485 284023 264513 284051
rect 264547 284023 264575 284051
rect 264609 284023 264637 284051
rect 264671 284023 264699 284051
rect 264485 283961 264513 283989
rect 264547 283961 264575 283989
rect 264609 283961 264637 283989
rect 264671 283961 264699 283989
rect 264485 275147 264513 275175
rect 264547 275147 264575 275175
rect 264609 275147 264637 275175
rect 264671 275147 264699 275175
rect 264485 275085 264513 275113
rect 264547 275085 264575 275113
rect 264609 275085 264637 275113
rect 264671 275085 264699 275113
rect 264485 275023 264513 275051
rect 264547 275023 264575 275051
rect 264609 275023 264637 275051
rect 264671 275023 264699 275051
rect 264485 274961 264513 274989
rect 264547 274961 264575 274989
rect 264609 274961 264637 274989
rect 264671 274961 264699 274989
rect 264485 266147 264513 266175
rect 264547 266147 264575 266175
rect 264609 266147 264637 266175
rect 264671 266147 264699 266175
rect 264485 266085 264513 266113
rect 264547 266085 264575 266113
rect 264609 266085 264637 266113
rect 264671 266085 264699 266113
rect 264485 266023 264513 266051
rect 264547 266023 264575 266051
rect 264609 266023 264637 266051
rect 264671 266023 264699 266051
rect 264485 265961 264513 265989
rect 264547 265961 264575 265989
rect 264609 265961 264637 265989
rect 264671 265961 264699 265989
rect 264485 257147 264513 257175
rect 264547 257147 264575 257175
rect 264609 257147 264637 257175
rect 264671 257147 264699 257175
rect 264485 257085 264513 257113
rect 264547 257085 264575 257113
rect 264609 257085 264637 257113
rect 264671 257085 264699 257113
rect 264485 257023 264513 257051
rect 264547 257023 264575 257051
rect 264609 257023 264637 257051
rect 264671 257023 264699 257051
rect 264485 256961 264513 256989
rect 264547 256961 264575 256989
rect 264609 256961 264637 256989
rect 264671 256961 264699 256989
rect 264485 248147 264513 248175
rect 264547 248147 264575 248175
rect 264609 248147 264637 248175
rect 264671 248147 264699 248175
rect 264485 248085 264513 248113
rect 264547 248085 264575 248113
rect 264609 248085 264637 248113
rect 264671 248085 264699 248113
rect 264485 248023 264513 248051
rect 264547 248023 264575 248051
rect 264609 248023 264637 248051
rect 264671 248023 264699 248051
rect 264485 247961 264513 247989
rect 264547 247961 264575 247989
rect 264609 247961 264637 247989
rect 264671 247961 264699 247989
rect 264485 239147 264513 239175
rect 264547 239147 264575 239175
rect 264609 239147 264637 239175
rect 264671 239147 264699 239175
rect 264485 239085 264513 239113
rect 264547 239085 264575 239113
rect 264609 239085 264637 239113
rect 264671 239085 264699 239113
rect 264485 239023 264513 239051
rect 264547 239023 264575 239051
rect 264609 239023 264637 239051
rect 264671 239023 264699 239051
rect 264485 238961 264513 238989
rect 264547 238961 264575 238989
rect 264609 238961 264637 238989
rect 264671 238961 264699 238989
rect 264485 230147 264513 230175
rect 264547 230147 264575 230175
rect 264609 230147 264637 230175
rect 264671 230147 264699 230175
rect 264485 230085 264513 230113
rect 264547 230085 264575 230113
rect 264609 230085 264637 230113
rect 264671 230085 264699 230113
rect 264485 230023 264513 230051
rect 264547 230023 264575 230051
rect 264609 230023 264637 230051
rect 264671 230023 264699 230051
rect 264485 229961 264513 229989
rect 264547 229961 264575 229989
rect 264609 229961 264637 229989
rect 264671 229961 264699 229989
rect 264485 221147 264513 221175
rect 264547 221147 264575 221175
rect 264609 221147 264637 221175
rect 264671 221147 264699 221175
rect 264485 221085 264513 221113
rect 264547 221085 264575 221113
rect 264609 221085 264637 221113
rect 264671 221085 264699 221113
rect 264485 221023 264513 221051
rect 264547 221023 264575 221051
rect 264609 221023 264637 221051
rect 264671 221023 264699 221051
rect 264485 220961 264513 220989
rect 264547 220961 264575 220989
rect 264609 220961 264637 220989
rect 264671 220961 264699 220989
rect 264485 212147 264513 212175
rect 264547 212147 264575 212175
rect 264609 212147 264637 212175
rect 264671 212147 264699 212175
rect 264485 212085 264513 212113
rect 264547 212085 264575 212113
rect 264609 212085 264637 212113
rect 264671 212085 264699 212113
rect 264485 212023 264513 212051
rect 264547 212023 264575 212051
rect 264609 212023 264637 212051
rect 264671 212023 264699 212051
rect 264485 211961 264513 211989
rect 264547 211961 264575 211989
rect 264609 211961 264637 211989
rect 264671 211961 264699 211989
rect 264485 203147 264513 203175
rect 264547 203147 264575 203175
rect 264609 203147 264637 203175
rect 264671 203147 264699 203175
rect 264485 203085 264513 203113
rect 264547 203085 264575 203113
rect 264609 203085 264637 203113
rect 264671 203085 264699 203113
rect 264485 203023 264513 203051
rect 264547 203023 264575 203051
rect 264609 203023 264637 203051
rect 264671 203023 264699 203051
rect 264485 202961 264513 202989
rect 264547 202961 264575 202989
rect 264609 202961 264637 202989
rect 264671 202961 264699 202989
rect 264485 194147 264513 194175
rect 264547 194147 264575 194175
rect 264609 194147 264637 194175
rect 264671 194147 264699 194175
rect 264485 194085 264513 194113
rect 264547 194085 264575 194113
rect 264609 194085 264637 194113
rect 264671 194085 264699 194113
rect 264485 194023 264513 194051
rect 264547 194023 264575 194051
rect 264609 194023 264637 194051
rect 264671 194023 264699 194051
rect 264485 193961 264513 193989
rect 264547 193961 264575 193989
rect 264609 193961 264637 193989
rect 264671 193961 264699 193989
rect 264485 185147 264513 185175
rect 264547 185147 264575 185175
rect 264609 185147 264637 185175
rect 264671 185147 264699 185175
rect 264485 185085 264513 185113
rect 264547 185085 264575 185113
rect 264609 185085 264637 185113
rect 264671 185085 264699 185113
rect 264485 185023 264513 185051
rect 264547 185023 264575 185051
rect 264609 185023 264637 185051
rect 264671 185023 264699 185051
rect 264485 184961 264513 184989
rect 264547 184961 264575 184989
rect 264609 184961 264637 184989
rect 264671 184961 264699 184989
rect 264485 176147 264513 176175
rect 264547 176147 264575 176175
rect 264609 176147 264637 176175
rect 264671 176147 264699 176175
rect 264485 176085 264513 176113
rect 264547 176085 264575 176113
rect 264609 176085 264637 176113
rect 264671 176085 264699 176113
rect 264485 176023 264513 176051
rect 264547 176023 264575 176051
rect 264609 176023 264637 176051
rect 264671 176023 264699 176051
rect 264485 175961 264513 175989
rect 264547 175961 264575 175989
rect 264609 175961 264637 175989
rect 264671 175961 264699 175989
rect 264485 167147 264513 167175
rect 264547 167147 264575 167175
rect 264609 167147 264637 167175
rect 264671 167147 264699 167175
rect 264485 167085 264513 167113
rect 264547 167085 264575 167113
rect 264609 167085 264637 167113
rect 264671 167085 264699 167113
rect 264485 167023 264513 167051
rect 264547 167023 264575 167051
rect 264609 167023 264637 167051
rect 264671 167023 264699 167051
rect 264485 166961 264513 166989
rect 264547 166961 264575 166989
rect 264609 166961 264637 166989
rect 264671 166961 264699 166989
rect 264485 158147 264513 158175
rect 264547 158147 264575 158175
rect 264609 158147 264637 158175
rect 264671 158147 264699 158175
rect 264485 158085 264513 158113
rect 264547 158085 264575 158113
rect 264609 158085 264637 158113
rect 264671 158085 264699 158113
rect 264485 158023 264513 158051
rect 264547 158023 264575 158051
rect 264609 158023 264637 158051
rect 264671 158023 264699 158051
rect 264485 157961 264513 157989
rect 264547 157961 264575 157989
rect 264609 157961 264637 157989
rect 264671 157961 264699 157989
rect 264485 149147 264513 149175
rect 264547 149147 264575 149175
rect 264609 149147 264637 149175
rect 264671 149147 264699 149175
rect 264485 149085 264513 149113
rect 264547 149085 264575 149113
rect 264609 149085 264637 149113
rect 264671 149085 264699 149113
rect 264485 149023 264513 149051
rect 264547 149023 264575 149051
rect 264609 149023 264637 149051
rect 264671 149023 264699 149051
rect 264485 148961 264513 148989
rect 264547 148961 264575 148989
rect 264609 148961 264637 148989
rect 264671 148961 264699 148989
rect 264485 140147 264513 140175
rect 264547 140147 264575 140175
rect 264609 140147 264637 140175
rect 264671 140147 264699 140175
rect 264485 140085 264513 140113
rect 264547 140085 264575 140113
rect 264609 140085 264637 140113
rect 264671 140085 264699 140113
rect 264485 140023 264513 140051
rect 264547 140023 264575 140051
rect 264609 140023 264637 140051
rect 264671 140023 264699 140051
rect 264485 139961 264513 139989
rect 264547 139961 264575 139989
rect 264609 139961 264637 139989
rect 264671 139961 264699 139989
rect 264485 131147 264513 131175
rect 264547 131147 264575 131175
rect 264609 131147 264637 131175
rect 264671 131147 264699 131175
rect 264485 131085 264513 131113
rect 264547 131085 264575 131113
rect 264609 131085 264637 131113
rect 264671 131085 264699 131113
rect 264485 131023 264513 131051
rect 264547 131023 264575 131051
rect 264609 131023 264637 131051
rect 264671 131023 264699 131051
rect 264485 130961 264513 130989
rect 264547 130961 264575 130989
rect 264609 130961 264637 130989
rect 264671 130961 264699 130989
rect 264485 122147 264513 122175
rect 264547 122147 264575 122175
rect 264609 122147 264637 122175
rect 264671 122147 264699 122175
rect 264485 122085 264513 122113
rect 264547 122085 264575 122113
rect 264609 122085 264637 122113
rect 264671 122085 264699 122113
rect 264485 122023 264513 122051
rect 264547 122023 264575 122051
rect 264609 122023 264637 122051
rect 264671 122023 264699 122051
rect 264485 121961 264513 121989
rect 264547 121961 264575 121989
rect 264609 121961 264637 121989
rect 264671 121961 264699 121989
rect 264485 113147 264513 113175
rect 264547 113147 264575 113175
rect 264609 113147 264637 113175
rect 264671 113147 264699 113175
rect 264485 113085 264513 113113
rect 264547 113085 264575 113113
rect 264609 113085 264637 113113
rect 264671 113085 264699 113113
rect 264485 113023 264513 113051
rect 264547 113023 264575 113051
rect 264609 113023 264637 113051
rect 264671 113023 264699 113051
rect 264485 112961 264513 112989
rect 264547 112961 264575 112989
rect 264609 112961 264637 112989
rect 264671 112961 264699 112989
rect 264485 104147 264513 104175
rect 264547 104147 264575 104175
rect 264609 104147 264637 104175
rect 264671 104147 264699 104175
rect 264485 104085 264513 104113
rect 264547 104085 264575 104113
rect 264609 104085 264637 104113
rect 264671 104085 264699 104113
rect 264485 104023 264513 104051
rect 264547 104023 264575 104051
rect 264609 104023 264637 104051
rect 264671 104023 264699 104051
rect 264485 103961 264513 103989
rect 264547 103961 264575 103989
rect 264609 103961 264637 103989
rect 264671 103961 264699 103989
rect 264485 95147 264513 95175
rect 264547 95147 264575 95175
rect 264609 95147 264637 95175
rect 264671 95147 264699 95175
rect 264485 95085 264513 95113
rect 264547 95085 264575 95113
rect 264609 95085 264637 95113
rect 264671 95085 264699 95113
rect 264485 95023 264513 95051
rect 264547 95023 264575 95051
rect 264609 95023 264637 95051
rect 264671 95023 264699 95051
rect 264485 94961 264513 94989
rect 264547 94961 264575 94989
rect 264609 94961 264637 94989
rect 264671 94961 264699 94989
rect 264485 86147 264513 86175
rect 264547 86147 264575 86175
rect 264609 86147 264637 86175
rect 264671 86147 264699 86175
rect 264485 86085 264513 86113
rect 264547 86085 264575 86113
rect 264609 86085 264637 86113
rect 264671 86085 264699 86113
rect 264485 86023 264513 86051
rect 264547 86023 264575 86051
rect 264609 86023 264637 86051
rect 264671 86023 264699 86051
rect 264485 85961 264513 85989
rect 264547 85961 264575 85989
rect 264609 85961 264637 85989
rect 264671 85961 264699 85989
rect 264485 77147 264513 77175
rect 264547 77147 264575 77175
rect 264609 77147 264637 77175
rect 264671 77147 264699 77175
rect 264485 77085 264513 77113
rect 264547 77085 264575 77113
rect 264609 77085 264637 77113
rect 264671 77085 264699 77113
rect 264485 77023 264513 77051
rect 264547 77023 264575 77051
rect 264609 77023 264637 77051
rect 264671 77023 264699 77051
rect 264485 76961 264513 76989
rect 264547 76961 264575 76989
rect 264609 76961 264637 76989
rect 264671 76961 264699 76989
rect 264485 68147 264513 68175
rect 264547 68147 264575 68175
rect 264609 68147 264637 68175
rect 264671 68147 264699 68175
rect 264485 68085 264513 68113
rect 264547 68085 264575 68113
rect 264609 68085 264637 68113
rect 264671 68085 264699 68113
rect 264485 68023 264513 68051
rect 264547 68023 264575 68051
rect 264609 68023 264637 68051
rect 264671 68023 264699 68051
rect 264485 67961 264513 67989
rect 264547 67961 264575 67989
rect 264609 67961 264637 67989
rect 264671 67961 264699 67989
rect 264485 59147 264513 59175
rect 264547 59147 264575 59175
rect 264609 59147 264637 59175
rect 264671 59147 264699 59175
rect 264485 59085 264513 59113
rect 264547 59085 264575 59113
rect 264609 59085 264637 59113
rect 264671 59085 264699 59113
rect 264485 59023 264513 59051
rect 264547 59023 264575 59051
rect 264609 59023 264637 59051
rect 264671 59023 264699 59051
rect 264485 58961 264513 58989
rect 264547 58961 264575 58989
rect 264609 58961 264637 58989
rect 264671 58961 264699 58989
rect 264485 50147 264513 50175
rect 264547 50147 264575 50175
rect 264609 50147 264637 50175
rect 264671 50147 264699 50175
rect 264485 50085 264513 50113
rect 264547 50085 264575 50113
rect 264609 50085 264637 50113
rect 264671 50085 264699 50113
rect 264485 50023 264513 50051
rect 264547 50023 264575 50051
rect 264609 50023 264637 50051
rect 264671 50023 264699 50051
rect 264485 49961 264513 49989
rect 264547 49961 264575 49989
rect 264609 49961 264637 49989
rect 264671 49961 264699 49989
rect 264485 41147 264513 41175
rect 264547 41147 264575 41175
rect 264609 41147 264637 41175
rect 264671 41147 264699 41175
rect 264485 41085 264513 41113
rect 264547 41085 264575 41113
rect 264609 41085 264637 41113
rect 264671 41085 264699 41113
rect 264485 41023 264513 41051
rect 264547 41023 264575 41051
rect 264609 41023 264637 41051
rect 264671 41023 264699 41051
rect 264485 40961 264513 40989
rect 264547 40961 264575 40989
rect 264609 40961 264637 40989
rect 264671 40961 264699 40989
rect 264485 32147 264513 32175
rect 264547 32147 264575 32175
rect 264609 32147 264637 32175
rect 264671 32147 264699 32175
rect 264485 32085 264513 32113
rect 264547 32085 264575 32113
rect 264609 32085 264637 32113
rect 264671 32085 264699 32113
rect 264485 32023 264513 32051
rect 264547 32023 264575 32051
rect 264609 32023 264637 32051
rect 264671 32023 264699 32051
rect 264485 31961 264513 31989
rect 264547 31961 264575 31989
rect 264609 31961 264637 31989
rect 264671 31961 264699 31989
rect 264485 23147 264513 23175
rect 264547 23147 264575 23175
rect 264609 23147 264637 23175
rect 264671 23147 264699 23175
rect 264485 23085 264513 23113
rect 264547 23085 264575 23113
rect 264609 23085 264637 23113
rect 264671 23085 264699 23113
rect 264485 23023 264513 23051
rect 264547 23023 264575 23051
rect 264609 23023 264637 23051
rect 264671 23023 264699 23051
rect 264485 22961 264513 22989
rect 264547 22961 264575 22989
rect 264609 22961 264637 22989
rect 264671 22961 264699 22989
rect 264485 14147 264513 14175
rect 264547 14147 264575 14175
rect 264609 14147 264637 14175
rect 264671 14147 264699 14175
rect 264485 14085 264513 14113
rect 264547 14085 264575 14113
rect 264609 14085 264637 14113
rect 264671 14085 264699 14113
rect 264485 14023 264513 14051
rect 264547 14023 264575 14051
rect 264609 14023 264637 14051
rect 264671 14023 264699 14051
rect 264485 13961 264513 13989
rect 264547 13961 264575 13989
rect 264609 13961 264637 13989
rect 264671 13961 264699 13989
rect 264485 5147 264513 5175
rect 264547 5147 264575 5175
rect 264609 5147 264637 5175
rect 264671 5147 264699 5175
rect 264485 5085 264513 5113
rect 264547 5085 264575 5113
rect 264609 5085 264637 5113
rect 264671 5085 264699 5113
rect 264485 5023 264513 5051
rect 264547 5023 264575 5051
rect 264609 5023 264637 5051
rect 264671 5023 264699 5051
rect 264485 4961 264513 4989
rect 264547 4961 264575 4989
rect 264609 4961 264637 4989
rect 264671 4961 264699 4989
rect 264485 -588 264513 -560
rect 264547 -588 264575 -560
rect 264609 -588 264637 -560
rect 264671 -588 264699 -560
rect 264485 -650 264513 -622
rect 264547 -650 264575 -622
rect 264609 -650 264637 -622
rect 264671 -650 264699 -622
rect 264485 -712 264513 -684
rect 264547 -712 264575 -684
rect 264609 -712 264637 -684
rect 264671 -712 264699 -684
rect 264485 -774 264513 -746
rect 264547 -774 264575 -746
rect 264609 -774 264637 -746
rect 264671 -774 264699 -746
rect 271625 298578 271653 298606
rect 271687 298578 271715 298606
rect 271749 298578 271777 298606
rect 271811 298578 271839 298606
rect 271625 298516 271653 298544
rect 271687 298516 271715 298544
rect 271749 298516 271777 298544
rect 271811 298516 271839 298544
rect 271625 298454 271653 298482
rect 271687 298454 271715 298482
rect 271749 298454 271777 298482
rect 271811 298454 271839 298482
rect 271625 298392 271653 298420
rect 271687 298392 271715 298420
rect 271749 298392 271777 298420
rect 271811 298392 271839 298420
rect 271625 290147 271653 290175
rect 271687 290147 271715 290175
rect 271749 290147 271777 290175
rect 271811 290147 271839 290175
rect 271625 290085 271653 290113
rect 271687 290085 271715 290113
rect 271749 290085 271777 290113
rect 271811 290085 271839 290113
rect 271625 290023 271653 290051
rect 271687 290023 271715 290051
rect 271749 290023 271777 290051
rect 271811 290023 271839 290051
rect 271625 289961 271653 289989
rect 271687 289961 271715 289989
rect 271749 289961 271777 289989
rect 271811 289961 271839 289989
rect 271625 281147 271653 281175
rect 271687 281147 271715 281175
rect 271749 281147 271777 281175
rect 271811 281147 271839 281175
rect 271625 281085 271653 281113
rect 271687 281085 271715 281113
rect 271749 281085 271777 281113
rect 271811 281085 271839 281113
rect 271625 281023 271653 281051
rect 271687 281023 271715 281051
rect 271749 281023 271777 281051
rect 271811 281023 271839 281051
rect 271625 280961 271653 280989
rect 271687 280961 271715 280989
rect 271749 280961 271777 280989
rect 271811 280961 271839 280989
rect 271625 272147 271653 272175
rect 271687 272147 271715 272175
rect 271749 272147 271777 272175
rect 271811 272147 271839 272175
rect 271625 272085 271653 272113
rect 271687 272085 271715 272113
rect 271749 272085 271777 272113
rect 271811 272085 271839 272113
rect 271625 272023 271653 272051
rect 271687 272023 271715 272051
rect 271749 272023 271777 272051
rect 271811 272023 271839 272051
rect 271625 271961 271653 271989
rect 271687 271961 271715 271989
rect 271749 271961 271777 271989
rect 271811 271961 271839 271989
rect 271625 263147 271653 263175
rect 271687 263147 271715 263175
rect 271749 263147 271777 263175
rect 271811 263147 271839 263175
rect 271625 263085 271653 263113
rect 271687 263085 271715 263113
rect 271749 263085 271777 263113
rect 271811 263085 271839 263113
rect 271625 263023 271653 263051
rect 271687 263023 271715 263051
rect 271749 263023 271777 263051
rect 271811 263023 271839 263051
rect 271625 262961 271653 262989
rect 271687 262961 271715 262989
rect 271749 262961 271777 262989
rect 271811 262961 271839 262989
rect 271625 254147 271653 254175
rect 271687 254147 271715 254175
rect 271749 254147 271777 254175
rect 271811 254147 271839 254175
rect 271625 254085 271653 254113
rect 271687 254085 271715 254113
rect 271749 254085 271777 254113
rect 271811 254085 271839 254113
rect 271625 254023 271653 254051
rect 271687 254023 271715 254051
rect 271749 254023 271777 254051
rect 271811 254023 271839 254051
rect 271625 253961 271653 253989
rect 271687 253961 271715 253989
rect 271749 253961 271777 253989
rect 271811 253961 271839 253989
rect 271625 245147 271653 245175
rect 271687 245147 271715 245175
rect 271749 245147 271777 245175
rect 271811 245147 271839 245175
rect 271625 245085 271653 245113
rect 271687 245085 271715 245113
rect 271749 245085 271777 245113
rect 271811 245085 271839 245113
rect 271625 245023 271653 245051
rect 271687 245023 271715 245051
rect 271749 245023 271777 245051
rect 271811 245023 271839 245051
rect 271625 244961 271653 244989
rect 271687 244961 271715 244989
rect 271749 244961 271777 244989
rect 271811 244961 271839 244989
rect 271625 236147 271653 236175
rect 271687 236147 271715 236175
rect 271749 236147 271777 236175
rect 271811 236147 271839 236175
rect 271625 236085 271653 236113
rect 271687 236085 271715 236113
rect 271749 236085 271777 236113
rect 271811 236085 271839 236113
rect 271625 236023 271653 236051
rect 271687 236023 271715 236051
rect 271749 236023 271777 236051
rect 271811 236023 271839 236051
rect 271625 235961 271653 235989
rect 271687 235961 271715 235989
rect 271749 235961 271777 235989
rect 271811 235961 271839 235989
rect 271625 227147 271653 227175
rect 271687 227147 271715 227175
rect 271749 227147 271777 227175
rect 271811 227147 271839 227175
rect 271625 227085 271653 227113
rect 271687 227085 271715 227113
rect 271749 227085 271777 227113
rect 271811 227085 271839 227113
rect 271625 227023 271653 227051
rect 271687 227023 271715 227051
rect 271749 227023 271777 227051
rect 271811 227023 271839 227051
rect 271625 226961 271653 226989
rect 271687 226961 271715 226989
rect 271749 226961 271777 226989
rect 271811 226961 271839 226989
rect 271625 218147 271653 218175
rect 271687 218147 271715 218175
rect 271749 218147 271777 218175
rect 271811 218147 271839 218175
rect 271625 218085 271653 218113
rect 271687 218085 271715 218113
rect 271749 218085 271777 218113
rect 271811 218085 271839 218113
rect 271625 218023 271653 218051
rect 271687 218023 271715 218051
rect 271749 218023 271777 218051
rect 271811 218023 271839 218051
rect 271625 217961 271653 217989
rect 271687 217961 271715 217989
rect 271749 217961 271777 217989
rect 271811 217961 271839 217989
rect 271625 209147 271653 209175
rect 271687 209147 271715 209175
rect 271749 209147 271777 209175
rect 271811 209147 271839 209175
rect 271625 209085 271653 209113
rect 271687 209085 271715 209113
rect 271749 209085 271777 209113
rect 271811 209085 271839 209113
rect 271625 209023 271653 209051
rect 271687 209023 271715 209051
rect 271749 209023 271777 209051
rect 271811 209023 271839 209051
rect 271625 208961 271653 208989
rect 271687 208961 271715 208989
rect 271749 208961 271777 208989
rect 271811 208961 271839 208989
rect 271625 200147 271653 200175
rect 271687 200147 271715 200175
rect 271749 200147 271777 200175
rect 271811 200147 271839 200175
rect 271625 200085 271653 200113
rect 271687 200085 271715 200113
rect 271749 200085 271777 200113
rect 271811 200085 271839 200113
rect 271625 200023 271653 200051
rect 271687 200023 271715 200051
rect 271749 200023 271777 200051
rect 271811 200023 271839 200051
rect 271625 199961 271653 199989
rect 271687 199961 271715 199989
rect 271749 199961 271777 199989
rect 271811 199961 271839 199989
rect 271625 191147 271653 191175
rect 271687 191147 271715 191175
rect 271749 191147 271777 191175
rect 271811 191147 271839 191175
rect 271625 191085 271653 191113
rect 271687 191085 271715 191113
rect 271749 191085 271777 191113
rect 271811 191085 271839 191113
rect 271625 191023 271653 191051
rect 271687 191023 271715 191051
rect 271749 191023 271777 191051
rect 271811 191023 271839 191051
rect 271625 190961 271653 190989
rect 271687 190961 271715 190989
rect 271749 190961 271777 190989
rect 271811 190961 271839 190989
rect 271625 182147 271653 182175
rect 271687 182147 271715 182175
rect 271749 182147 271777 182175
rect 271811 182147 271839 182175
rect 271625 182085 271653 182113
rect 271687 182085 271715 182113
rect 271749 182085 271777 182113
rect 271811 182085 271839 182113
rect 271625 182023 271653 182051
rect 271687 182023 271715 182051
rect 271749 182023 271777 182051
rect 271811 182023 271839 182051
rect 271625 181961 271653 181989
rect 271687 181961 271715 181989
rect 271749 181961 271777 181989
rect 271811 181961 271839 181989
rect 271625 173147 271653 173175
rect 271687 173147 271715 173175
rect 271749 173147 271777 173175
rect 271811 173147 271839 173175
rect 271625 173085 271653 173113
rect 271687 173085 271715 173113
rect 271749 173085 271777 173113
rect 271811 173085 271839 173113
rect 271625 173023 271653 173051
rect 271687 173023 271715 173051
rect 271749 173023 271777 173051
rect 271811 173023 271839 173051
rect 271625 172961 271653 172989
rect 271687 172961 271715 172989
rect 271749 172961 271777 172989
rect 271811 172961 271839 172989
rect 271625 164147 271653 164175
rect 271687 164147 271715 164175
rect 271749 164147 271777 164175
rect 271811 164147 271839 164175
rect 271625 164085 271653 164113
rect 271687 164085 271715 164113
rect 271749 164085 271777 164113
rect 271811 164085 271839 164113
rect 271625 164023 271653 164051
rect 271687 164023 271715 164051
rect 271749 164023 271777 164051
rect 271811 164023 271839 164051
rect 271625 163961 271653 163989
rect 271687 163961 271715 163989
rect 271749 163961 271777 163989
rect 271811 163961 271839 163989
rect 271625 155147 271653 155175
rect 271687 155147 271715 155175
rect 271749 155147 271777 155175
rect 271811 155147 271839 155175
rect 271625 155085 271653 155113
rect 271687 155085 271715 155113
rect 271749 155085 271777 155113
rect 271811 155085 271839 155113
rect 271625 155023 271653 155051
rect 271687 155023 271715 155051
rect 271749 155023 271777 155051
rect 271811 155023 271839 155051
rect 271625 154961 271653 154989
rect 271687 154961 271715 154989
rect 271749 154961 271777 154989
rect 271811 154961 271839 154989
rect 271625 146147 271653 146175
rect 271687 146147 271715 146175
rect 271749 146147 271777 146175
rect 271811 146147 271839 146175
rect 271625 146085 271653 146113
rect 271687 146085 271715 146113
rect 271749 146085 271777 146113
rect 271811 146085 271839 146113
rect 271625 146023 271653 146051
rect 271687 146023 271715 146051
rect 271749 146023 271777 146051
rect 271811 146023 271839 146051
rect 271625 145961 271653 145989
rect 271687 145961 271715 145989
rect 271749 145961 271777 145989
rect 271811 145961 271839 145989
rect 271625 137147 271653 137175
rect 271687 137147 271715 137175
rect 271749 137147 271777 137175
rect 271811 137147 271839 137175
rect 271625 137085 271653 137113
rect 271687 137085 271715 137113
rect 271749 137085 271777 137113
rect 271811 137085 271839 137113
rect 271625 137023 271653 137051
rect 271687 137023 271715 137051
rect 271749 137023 271777 137051
rect 271811 137023 271839 137051
rect 271625 136961 271653 136989
rect 271687 136961 271715 136989
rect 271749 136961 271777 136989
rect 271811 136961 271839 136989
rect 271625 128147 271653 128175
rect 271687 128147 271715 128175
rect 271749 128147 271777 128175
rect 271811 128147 271839 128175
rect 271625 128085 271653 128113
rect 271687 128085 271715 128113
rect 271749 128085 271777 128113
rect 271811 128085 271839 128113
rect 271625 128023 271653 128051
rect 271687 128023 271715 128051
rect 271749 128023 271777 128051
rect 271811 128023 271839 128051
rect 271625 127961 271653 127989
rect 271687 127961 271715 127989
rect 271749 127961 271777 127989
rect 271811 127961 271839 127989
rect 271625 119147 271653 119175
rect 271687 119147 271715 119175
rect 271749 119147 271777 119175
rect 271811 119147 271839 119175
rect 271625 119085 271653 119113
rect 271687 119085 271715 119113
rect 271749 119085 271777 119113
rect 271811 119085 271839 119113
rect 271625 119023 271653 119051
rect 271687 119023 271715 119051
rect 271749 119023 271777 119051
rect 271811 119023 271839 119051
rect 271625 118961 271653 118989
rect 271687 118961 271715 118989
rect 271749 118961 271777 118989
rect 271811 118961 271839 118989
rect 271625 110147 271653 110175
rect 271687 110147 271715 110175
rect 271749 110147 271777 110175
rect 271811 110147 271839 110175
rect 271625 110085 271653 110113
rect 271687 110085 271715 110113
rect 271749 110085 271777 110113
rect 271811 110085 271839 110113
rect 271625 110023 271653 110051
rect 271687 110023 271715 110051
rect 271749 110023 271777 110051
rect 271811 110023 271839 110051
rect 271625 109961 271653 109989
rect 271687 109961 271715 109989
rect 271749 109961 271777 109989
rect 271811 109961 271839 109989
rect 271625 101147 271653 101175
rect 271687 101147 271715 101175
rect 271749 101147 271777 101175
rect 271811 101147 271839 101175
rect 271625 101085 271653 101113
rect 271687 101085 271715 101113
rect 271749 101085 271777 101113
rect 271811 101085 271839 101113
rect 271625 101023 271653 101051
rect 271687 101023 271715 101051
rect 271749 101023 271777 101051
rect 271811 101023 271839 101051
rect 271625 100961 271653 100989
rect 271687 100961 271715 100989
rect 271749 100961 271777 100989
rect 271811 100961 271839 100989
rect 271625 92147 271653 92175
rect 271687 92147 271715 92175
rect 271749 92147 271777 92175
rect 271811 92147 271839 92175
rect 271625 92085 271653 92113
rect 271687 92085 271715 92113
rect 271749 92085 271777 92113
rect 271811 92085 271839 92113
rect 271625 92023 271653 92051
rect 271687 92023 271715 92051
rect 271749 92023 271777 92051
rect 271811 92023 271839 92051
rect 271625 91961 271653 91989
rect 271687 91961 271715 91989
rect 271749 91961 271777 91989
rect 271811 91961 271839 91989
rect 271625 83147 271653 83175
rect 271687 83147 271715 83175
rect 271749 83147 271777 83175
rect 271811 83147 271839 83175
rect 271625 83085 271653 83113
rect 271687 83085 271715 83113
rect 271749 83085 271777 83113
rect 271811 83085 271839 83113
rect 271625 83023 271653 83051
rect 271687 83023 271715 83051
rect 271749 83023 271777 83051
rect 271811 83023 271839 83051
rect 271625 82961 271653 82989
rect 271687 82961 271715 82989
rect 271749 82961 271777 82989
rect 271811 82961 271839 82989
rect 271625 74147 271653 74175
rect 271687 74147 271715 74175
rect 271749 74147 271777 74175
rect 271811 74147 271839 74175
rect 271625 74085 271653 74113
rect 271687 74085 271715 74113
rect 271749 74085 271777 74113
rect 271811 74085 271839 74113
rect 271625 74023 271653 74051
rect 271687 74023 271715 74051
rect 271749 74023 271777 74051
rect 271811 74023 271839 74051
rect 271625 73961 271653 73989
rect 271687 73961 271715 73989
rect 271749 73961 271777 73989
rect 271811 73961 271839 73989
rect 271625 65147 271653 65175
rect 271687 65147 271715 65175
rect 271749 65147 271777 65175
rect 271811 65147 271839 65175
rect 271625 65085 271653 65113
rect 271687 65085 271715 65113
rect 271749 65085 271777 65113
rect 271811 65085 271839 65113
rect 271625 65023 271653 65051
rect 271687 65023 271715 65051
rect 271749 65023 271777 65051
rect 271811 65023 271839 65051
rect 271625 64961 271653 64989
rect 271687 64961 271715 64989
rect 271749 64961 271777 64989
rect 271811 64961 271839 64989
rect 271625 56147 271653 56175
rect 271687 56147 271715 56175
rect 271749 56147 271777 56175
rect 271811 56147 271839 56175
rect 271625 56085 271653 56113
rect 271687 56085 271715 56113
rect 271749 56085 271777 56113
rect 271811 56085 271839 56113
rect 271625 56023 271653 56051
rect 271687 56023 271715 56051
rect 271749 56023 271777 56051
rect 271811 56023 271839 56051
rect 271625 55961 271653 55989
rect 271687 55961 271715 55989
rect 271749 55961 271777 55989
rect 271811 55961 271839 55989
rect 271625 47147 271653 47175
rect 271687 47147 271715 47175
rect 271749 47147 271777 47175
rect 271811 47147 271839 47175
rect 271625 47085 271653 47113
rect 271687 47085 271715 47113
rect 271749 47085 271777 47113
rect 271811 47085 271839 47113
rect 271625 47023 271653 47051
rect 271687 47023 271715 47051
rect 271749 47023 271777 47051
rect 271811 47023 271839 47051
rect 271625 46961 271653 46989
rect 271687 46961 271715 46989
rect 271749 46961 271777 46989
rect 271811 46961 271839 46989
rect 271625 38147 271653 38175
rect 271687 38147 271715 38175
rect 271749 38147 271777 38175
rect 271811 38147 271839 38175
rect 271625 38085 271653 38113
rect 271687 38085 271715 38113
rect 271749 38085 271777 38113
rect 271811 38085 271839 38113
rect 271625 38023 271653 38051
rect 271687 38023 271715 38051
rect 271749 38023 271777 38051
rect 271811 38023 271839 38051
rect 271625 37961 271653 37989
rect 271687 37961 271715 37989
rect 271749 37961 271777 37989
rect 271811 37961 271839 37989
rect 271625 29147 271653 29175
rect 271687 29147 271715 29175
rect 271749 29147 271777 29175
rect 271811 29147 271839 29175
rect 271625 29085 271653 29113
rect 271687 29085 271715 29113
rect 271749 29085 271777 29113
rect 271811 29085 271839 29113
rect 271625 29023 271653 29051
rect 271687 29023 271715 29051
rect 271749 29023 271777 29051
rect 271811 29023 271839 29051
rect 271625 28961 271653 28989
rect 271687 28961 271715 28989
rect 271749 28961 271777 28989
rect 271811 28961 271839 28989
rect 271625 20147 271653 20175
rect 271687 20147 271715 20175
rect 271749 20147 271777 20175
rect 271811 20147 271839 20175
rect 271625 20085 271653 20113
rect 271687 20085 271715 20113
rect 271749 20085 271777 20113
rect 271811 20085 271839 20113
rect 271625 20023 271653 20051
rect 271687 20023 271715 20051
rect 271749 20023 271777 20051
rect 271811 20023 271839 20051
rect 271625 19961 271653 19989
rect 271687 19961 271715 19989
rect 271749 19961 271777 19989
rect 271811 19961 271839 19989
rect 271625 11147 271653 11175
rect 271687 11147 271715 11175
rect 271749 11147 271777 11175
rect 271811 11147 271839 11175
rect 271625 11085 271653 11113
rect 271687 11085 271715 11113
rect 271749 11085 271777 11113
rect 271811 11085 271839 11113
rect 271625 11023 271653 11051
rect 271687 11023 271715 11051
rect 271749 11023 271777 11051
rect 271811 11023 271839 11051
rect 271625 10961 271653 10989
rect 271687 10961 271715 10989
rect 271749 10961 271777 10989
rect 271811 10961 271839 10989
rect 271625 2147 271653 2175
rect 271687 2147 271715 2175
rect 271749 2147 271777 2175
rect 271811 2147 271839 2175
rect 271625 2085 271653 2113
rect 271687 2085 271715 2113
rect 271749 2085 271777 2113
rect 271811 2085 271839 2113
rect 271625 2023 271653 2051
rect 271687 2023 271715 2051
rect 271749 2023 271777 2051
rect 271811 2023 271839 2051
rect 271625 1961 271653 1989
rect 271687 1961 271715 1989
rect 271749 1961 271777 1989
rect 271811 1961 271839 1989
rect 271625 -108 271653 -80
rect 271687 -108 271715 -80
rect 271749 -108 271777 -80
rect 271811 -108 271839 -80
rect 271625 -170 271653 -142
rect 271687 -170 271715 -142
rect 271749 -170 271777 -142
rect 271811 -170 271839 -142
rect 271625 -232 271653 -204
rect 271687 -232 271715 -204
rect 271749 -232 271777 -204
rect 271811 -232 271839 -204
rect 271625 -294 271653 -266
rect 271687 -294 271715 -266
rect 271749 -294 271777 -266
rect 271811 -294 271839 -266
rect 273485 299058 273513 299086
rect 273547 299058 273575 299086
rect 273609 299058 273637 299086
rect 273671 299058 273699 299086
rect 273485 298996 273513 299024
rect 273547 298996 273575 299024
rect 273609 298996 273637 299024
rect 273671 298996 273699 299024
rect 273485 298934 273513 298962
rect 273547 298934 273575 298962
rect 273609 298934 273637 298962
rect 273671 298934 273699 298962
rect 273485 298872 273513 298900
rect 273547 298872 273575 298900
rect 273609 298872 273637 298900
rect 273671 298872 273699 298900
rect 273485 293147 273513 293175
rect 273547 293147 273575 293175
rect 273609 293147 273637 293175
rect 273671 293147 273699 293175
rect 273485 293085 273513 293113
rect 273547 293085 273575 293113
rect 273609 293085 273637 293113
rect 273671 293085 273699 293113
rect 273485 293023 273513 293051
rect 273547 293023 273575 293051
rect 273609 293023 273637 293051
rect 273671 293023 273699 293051
rect 273485 292961 273513 292989
rect 273547 292961 273575 292989
rect 273609 292961 273637 292989
rect 273671 292961 273699 292989
rect 273485 284147 273513 284175
rect 273547 284147 273575 284175
rect 273609 284147 273637 284175
rect 273671 284147 273699 284175
rect 273485 284085 273513 284113
rect 273547 284085 273575 284113
rect 273609 284085 273637 284113
rect 273671 284085 273699 284113
rect 273485 284023 273513 284051
rect 273547 284023 273575 284051
rect 273609 284023 273637 284051
rect 273671 284023 273699 284051
rect 273485 283961 273513 283989
rect 273547 283961 273575 283989
rect 273609 283961 273637 283989
rect 273671 283961 273699 283989
rect 273485 275147 273513 275175
rect 273547 275147 273575 275175
rect 273609 275147 273637 275175
rect 273671 275147 273699 275175
rect 273485 275085 273513 275113
rect 273547 275085 273575 275113
rect 273609 275085 273637 275113
rect 273671 275085 273699 275113
rect 273485 275023 273513 275051
rect 273547 275023 273575 275051
rect 273609 275023 273637 275051
rect 273671 275023 273699 275051
rect 273485 274961 273513 274989
rect 273547 274961 273575 274989
rect 273609 274961 273637 274989
rect 273671 274961 273699 274989
rect 273485 266147 273513 266175
rect 273547 266147 273575 266175
rect 273609 266147 273637 266175
rect 273671 266147 273699 266175
rect 273485 266085 273513 266113
rect 273547 266085 273575 266113
rect 273609 266085 273637 266113
rect 273671 266085 273699 266113
rect 273485 266023 273513 266051
rect 273547 266023 273575 266051
rect 273609 266023 273637 266051
rect 273671 266023 273699 266051
rect 273485 265961 273513 265989
rect 273547 265961 273575 265989
rect 273609 265961 273637 265989
rect 273671 265961 273699 265989
rect 273485 257147 273513 257175
rect 273547 257147 273575 257175
rect 273609 257147 273637 257175
rect 273671 257147 273699 257175
rect 273485 257085 273513 257113
rect 273547 257085 273575 257113
rect 273609 257085 273637 257113
rect 273671 257085 273699 257113
rect 273485 257023 273513 257051
rect 273547 257023 273575 257051
rect 273609 257023 273637 257051
rect 273671 257023 273699 257051
rect 273485 256961 273513 256989
rect 273547 256961 273575 256989
rect 273609 256961 273637 256989
rect 273671 256961 273699 256989
rect 273485 248147 273513 248175
rect 273547 248147 273575 248175
rect 273609 248147 273637 248175
rect 273671 248147 273699 248175
rect 273485 248085 273513 248113
rect 273547 248085 273575 248113
rect 273609 248085 273637 248113
rect 273671 248085 273699 248113
rect 273485 248023 273513 248051
rect 273547 248023 273575 248051
rect 273609 248023 273637 248051
rect 273671 248023 273699 248051
rect 273485 247961 273513 247989
rect 273547 247961 273575 247989
rect 273609 247961 273637 247989
rect 273671 247961 273699 247989
rect 273485 239147 273513 239175
rect 273547 239147 273575 239175
rect 273609 239147 273637 239175
rect 273671 239147 273699 239175
rect 273485 239085 273513 239113
rect 273547 239085 273575 239113
rect 273609 239085 273637 239113
rect 273671 239085 273699 239113
rect 273485 239023 273513 239051
rect 273547 239023 273575 239051
rect 273609 239023 273637 239051
rect 273671 239023 273699 239051
rect 273485 238961 273513 238989
rect 273547 238961 273575 238989
rect 273609 238961 273637 238989
rect 273671 238961 273699 238989
rect 273485 230147 273513 230175
rect 273547 230147 273575 230175
rect 273609 230147 273637 230175
rect 273671 230147 273699 230175
rect 273485 230085 273513 230113
rect 273547 230085 273575 230113
rect 273609 230085 273637 230113
rect 273671 230085 273699 230113
rect 273485 230023 273513 230051
rect 273547 230023 273575 230051
rect 273609 230023 273637 230051
rect 273671 230023 273699 230051
rect 273485 229961 273513 229989
rect 273547 229961 273575 229989
rect 273609 229961 273637 229989
rect 273671 229961 273699 229989
rect 273485 221147 273513 221175
rect 273547 221147 273575 221175
rect 273609 221147 273637 221175
rect 273671 221147 273699 221175
rect 273485 221085 273513 221113
rect 273547 221085 273575 221113
rect 273609 221085 273637 221113
rect 273671 221085 273699 221113
rect 273485 221023 273513 221051
rect 273547 221023 273575 221051
rect 273609 221023 273637 221051
rect 273671 221023 273699 221051
rect 273485 220961 273513 220989
rect 273547 220961 273575 220989
rect 273609 220961 273637 220989
rect 273671 220961 273699 220989
rect 273485 212147 273513 212175
rect 273547 212147 273575 212175
rect 273609 212147 273637 212175
rect 273671 212147 273699 212175
rect 273485 212085 273513 212113
rect 273547 212085 273575 212113
rect 273609 212085 273637 212113
rect 273671 212085 273699 212113
rect 273485 212023 273513 212051
rect 273547 212023 273575 212051
rect 273609 212023 273637 212051
rect 273671 212023 273699 212051
rect 273485 211961 273513 211989
rect 273547 211961 273575 211989
rect 273609 211961 273637 211989
rect 273671 211961 273699 211989
rect 273485 203147 273513 203175
rect 273547 203147 273575 203175
rect 273609 203147 273637 203175
rect 273671 203147 273699 203175
rect 273485 203085 273513 203113
rect 273547 203085 273575 203113
rect 273609 203085 273637 203113
rect 273671 203085 273699 203113
rect 273485 203023 273513 203051
rect 273547 203023 273575 203051
rect 273609 203023 273637 203051
rect 273671 203023 273699 203051
rect 273485 202961 273513 202989
rect 273547 202961 273575 202989
rect 273609 202961 273637 202989
rect 273671 202961 273699 202989
rect 273485 194147 273513 194175
rect 273547 194147 273575 194175
rect 273609 194147 273637 194175
rect 273671 194147 273699 194175
rect 273485 194085 273513 194113
rect 273547 194085 273575 194113
rect 273609 194085 273637 194113
rect 273671 194085 273699 194113
rect 273485 194023 273513 194051
rect 273547 194023 273575 194051
rect 273609 194023 273637 194051
rect 273671 194023 273699 194051
rect 273485 193961 273513 193989
rect 273547 193961 273575 193989
rect 273609 193961 273637 193989
rect 273671 193961 273699 193989
rect 273485 185147 273513 185175
rect 273547 185147 273575 185175
rect 273609 185147 273637 185175
rect 273671 185147 273699 185175
rect 273485 185085 273513 185113
rect 273547 185085 273575 185113
rect 273609 185085 273637 185113
rect 273671 185085 273699 185113
rect 273485 185023 273513 185051
rect 273547 185023 273575 185051
rect 273609 185023 273637 185051
rect 273671 185023 273699 185051
rect 273485 184961 273513 184989
rect 273547 184961 273575 184989
rect 273609 184961 273637 184989
rect 273671 184961 273699 184989
rect 273485 176147 273513 176175
rect 273547 176147 273575 176175
rect 273609 176147 273637 176175
rect 273671 176147 273699 176175
rect 273485 176085 273513 176113
rect 273547 176085 273575 176113
rect 273609 176085 273637 176113
rect 273671 176085 273699 176113
rect 273485 176023 273513 176051
rect 273547 176023 273575 176051
rect 273609 176023 273637 176051
rect 273671 176023 273699 176051
rect 273485 175961 273513 175989
rect 273547 175961 273575 175989
rect 273609 175961 273637 175989
rect 273671 175961 273699 175989
rect 273485 167147 273513 167175
rect 273547 167147 273575 167175
rect 273609 167147 273637 167175
rect 273671 167147 273699 167175
rect 273485 167085 273513 167113
rect 273547 167085 273575 167113
rect 273609 167085 273637 167113
rect 273671 167085 273699 167113
rect 273485 167023 273513 167051
rect 273547 167023 273575 167051
rect 273609 167023 273637 167051
rect 273671 167023 273699 167051
rect 273485 166961 273513 166989
rect 273547 166961 273575 166989
rect 273609 166961 273637 166989
rect 273671 166961 273699 166989
rect 273485 158147 273513 158175
rect 273547 158147 273575 158175
rect 273609 158147 273637 158175
rect 273671 158147 273699 158175
rect 273485 158085 273513 158113
rect 273547 158085 273575 158113
rect 273609 158085 273637 158113
rect 273671 158085 273699 158113
rect 273485 158023 273513 158051
rect 273547 158023 273575 158051
rect 273609 158023 273637 158051
rect 273671 158023 273699 158051
rect 273485 157961 273513 157989
rect 273547 157961 273575 157989
rect 273609 157961 273637 157989
rect 273671 157961 273699 157989
rect 273485 149147 273513 149175
rect 273547 149147 273575 149175
rect 273609 149147 273637 149175
rect 273671 149147 273699 149175
rect 273485 149085 273513 149113
rect 273547 149085 273575 149113
rect 273609 149085 273637 149113
rect 273671 149085 273699 149113
rect 273485 149023 273513 149051
rect 273547 149023 273575 149051
rect 273609 149023 273637 149051
rect 273671 149023 273699 149051
rect 273485 148961 273513 148989
rect 273547 148961 273575 148989
rect 273609 148961 273637 148989
rect 273671 148961 273699 148989
rect 273485 140147 273513 140175
rect 273547 140147 273575 140175
rect 273609 140147 273637 140175
rect 273671 140147 273699 140175
rect 273485 140085 273513 140113
rect 273547 140085 273575 140113
rect 273609 140085 273637 140113
rect 273671 140085 273699 140113
rect 273485 140023 273513 140051
rect 273547 140023 273575 140051
rect 273609 140023 273637 140051
rect 273671 140023 273699 140051
rect 273485 139961 273513 139989
rect 273547 139961 273575 139989
rect 273609 139961 273637 139989
rect 273671 139961 273699 139989
rect 273485 131147 273513 131175
rect 273547 131147 273575 131175
rect 273609 131147 273637 131175
rect 273671 131147 273699 131175
rect 273485 131085 273513 131113
rect 273547 131085 273575 131113
rect 273609 131085 273637 131113
rect 273671 131085 273699 131113
rect 273485 131023 273513 131051
rect 273547 131023 273575 131051
rect 273609 131023 273637 131051
rect 273671 131023 273699 131051
rect 273485 130961 273513 130989
rect 273547 130961 273575 130989
rect 273609 130961 273637 130989
rect 273671 130961 273699 130989
rect 273485 122147 273513 122175
rect 273547 122147 273575 122175
rect 273609 122147 273637 122175
rect 273671 122147 273699 122175
rect 273485 122085 273513 122113
rect 273547 122085 273575 122113
rect 273609 122085 273637 122113
rect 273671 122085 273699 122113
rect 273485 122023 273513 122051
rect 273547 122023 273575 122051
rect 273609 122023 273637 122051
rect 273671 122023 273699 122051
rect 273485 121961 273513 121989
rect 273547 121961 273575 121989
rect 273609 121961 273637 121989
rect 273671 121961 273699 121989
rect 273485 113147 273513 113175
rect 273547 113147 273575 113175
rect 273609 113147 273637 113175
rect 273671 113147 273699 113175
rect 273485 113085 273513 113113
rect 273547 113085 273575 113113
rect 273609 113085 273637 113113
rect 273671 113085 273699 113113
rect 273485 113023 273513 113051
rect 273547 113023 273575 113051
rect 273609 113023 273637 113051
rect 273671 113023 273699 113051
rect 273485 112961 273513 112989
rect 273547 112961 273575 112989
rect 273609 112961 273637 112989
rect 273671 112961 273699 112989
rect 273485 104147 273513 104175
rect 273547 104147 273575 104175
rect 273609 104147 273637 104175
rect 273671 104147 273699 104175
rect 273485 104085 273513 104113
rect 273547 104085 273575 104113
rect 273609 104085 273637 104113
rect 273671 104085 273699 104113
rect 273485 104023 273513 104051
rect 273547 104023 273575 104051
rect 273609 104023 273637 104051
rect 273671 104023 273699 104051
rect 273485 103961 273513 103989
rect 273547 103961 273575 103989
rect 273609 103961 273637 103989
rect 273671 103961 273699 103989
rect 273485 95147 273513 95175
rect 273547 95147 273575 95175
rect 273609 95147 273637 95175
rect 273671 95147 273699 95175
rect 273485 95085 273513 95113
rect 273547 95085 273575 95113
rect 273609 95085 273637 95113
rect 273671 95085 273699 95113
rect 273485 95023 273513 95051
rect 273547 95023 273575 95051
rect 273609 95023 273637 95051
rect 273671 95023 273699 95051
rect 273485 94961 273513 94989
rect 273547 94961 273575 94989
rect 273609 94961 273637 94989
rect 273671 94961 273699 94989
rect 273485 86147 273513 86175
rect 273547 86147 273575 86175
rect 273609 86147 273637 86175
rect 273671 86147 273699 86175
rect 273485 86085 273513 86113
rect 273547 86085 273575 86113
rect 273609 86085 273637 86113
rect 273671 86085 273699 86113
rect 273485 86023 273513 86051
rect 273547 86023 273575 86051
rect 273609 86023 273637 86051
rect 273671 86023 273699 86051
rect 273485 85961 273513 85989
rect 273547 85961 273575 85989
rect 273609 85961 273637 85989
rect 273671 85961 273699 85989
rect 273485 77147 273513 77175
rect 273547 77147 273575 77175
rect 273609 77147 273637 77175
rect 273671 77147 273699 77175
rect 273485 77085 273513 77113
rect 273547 77085 273575 77113
rect 273609 77085 273637 77113
rect 273671 77085 273699 77113
rect 273485 77023 273513 77051
rect 273547 77023 273575 77051
rect 273609 77023 273637 77051
rect 273671 77023 273699 77051
rect 273485 76961 273513 76989
rect 273547 76961 273575 76989
rect 273609 76961 273637 76989
rect 273671 76961 273699 76989
rect 273485 68147 273513 68175
rect 273547 68147 273575 68175
rect 273609 68147 273637 68175
rect 273671 68147 273699 68175
rect 273485 68085 273513 68113
rect 273547 68085 273575 68113
rect 273609 68085 273637 68113
rect 273671 68085 273699 68113
rect 273485 68023 273513 68051
rect 273547 68023 273575 68051
rect 273609 68023 273637 68051
rect 273671 68023 273699 68051
rect 273485 67961 273513 67989
rect 273547 67961 273575 67989
rect 273609 67961 273637 67989
rect 273671 67961 273699 67989
rect 273485 59147 273513 59175
rect 273547 59147 273575 59175
rect 273609 59147 273637 59175
rect 273671 59147 273699 59175
rect 273485 59085 273513 59113
rect 273547 59085 273575 59113
rect 273609 59085 273637 59113
rect 273671 59085 273699 59113
rect 273485 59023 273513 59051
rect 273547 59023 273575 59051
rect 273609 59023 273637 59051
rect 273671 59023 273699 59051
rect 273485 58961 273513 58989
rect 273547 58961 273575 58989
rect 273609 58961 273637 58989
rect 273671 58961 273699 58989
rect 273485 50147 273513 50175
rect 273547 50147 273575 50175
rect 273609 50147 273637 50175
rect 273671 50147 273699 50175
rect 273485 50085 273513 50113
rect 273547 50085 273575 50113
rect 273609 50085 273637 50113
rect 273671 50085 273699 50113
rect 273485 50023 273513 50051
rect 273547 50023 273575 50051
rect 273609 50023 273637 50051
rect 273671 50023 273699 50051
rect 273485 49961 273513 49989
rect 273547 49961 273575 49989
rect 273609 49961 273637 49989
rect 273671 49961 273699 49989
rect 273485 41147 273513 41175
rect 273547 41147 273575 41175
rect 273609 41147 273637 41175
rect 273671 41147 273699 41175
rect 273485 41085 273513 41113
rect 273547 41085 273575 41113
rect 273609 41085 273637 41113
rect 273671 41085 273699 41113
rect 273485 41023 273513 41051
rect 273547 41023 273575 41051
rect 273609 41023 273637 41051
rect 273671 41023 273699 41051
rect 273485 40961 273513 40989
rect 273547 40961 273575 40989
rect 273609 40961 273637 40989
rect 273671 40961 273699 40989
rect 273485 32147 273513 32175
rect 273547 32147 273575 32175
rect 273609 32147 273637 32175
rect 273671 32147 273699 32175
rect 273485 32085 273513 32113
rect 273547 32085 273575 32113
rect 273609 32085 273637 32113
rect 273671 32085 273699 32113
rect 273485 32023 273513 32051
rect 273547 32023 273575 32051
rect 273609 32023 273637 32051
rect 273671 32023 273699 32051
rect 273485 31961 273513 31989
rect 273547 31961 273575 31989
rect 273609 31961 273637 31989
rect 273671 31961 273699 31989
rect 273485 23147 273513 23175
rect 273547 23147 273575 23175
rect 273609 23147 273637 23175
rect 273671 23147 273699 23175
rect 273485 23085 273513 23113
rect 273547 23085 273575 23113
rect 273609 23085 273637 23113
rect 273671 23085 273699 23113
rect 273485 23023 273513 23051
rect 273547 23023 273575 23051
rect 273609 23023 273637 23051
rect 273671 23023 273699 23051
rect 273485 22961 273513 22989
rect 273547 22961 273575 22989
rect 273609 22961 273637 22989
rect 273671 22961 273699 22989
rect 273485 14147 273513 14175
rect 273547 14147 273575 14175
rect 273609 14147 273637 14175
rect 273671 14147 273699 14175
rect 273485 14085 273513 14113
rect 273547 14085 273575 14113
rect 273609 14085 273637 14113
rect 273671 14085 273699 14113
rect 273485 14023 273513 14051
rect 273547 14023 273575 14051
rect 273609 14023 273637 14051
rect 273671 14023 273699 14051
rect 273485 13961 273513 13989
rect 273547 13961 273575 13989
rect 273609 13961 273637 13989
rect 273671 13961 273699 13989
rect 273485 5147 273513 5175
rect 273547 5147 273575 5175
rect 273609 5147 273637 5175
rect 273671 5147 273699 5175
rect 273485 5085 273513 5113
rect 273547 5085 273575 5113
rect 273609 5085 273637 5113
rect 273671 5085 273699 5113
rect 273485 5023 273513 5051
rect 273547 5023 273575 5051
rect 273609 5023 273637 5051
rect 273671 5023 273699 5051
rect 273485 4961 273513 4989
rect 273547 4961 273575 4989
rect 273609 4961 273637 4989
rect 273671 4961 273699 4989
rect 273485 -588 273513 -560
rect 273547 -588 273575 -560
rect 273609 -588 273637 -560
rect 273671 -588 273699 -560
rect 273485 -650 273513 -622
rect 273547 -650 273575 -622
rect 273609 -650 273637 -622
rect 273671 -650 273699 -622
rect 273485 -712 273513 -684
rect 273547 -712 273575 -684
rect 273609 -712 273637 -684
rect 273671 -712 273699 -684
rect 273485 -774 273513 -746
rect 273547 -774 273575 -746
rect 273609 -774 273637 -746
rect 273671 -774 273699 -746
rect 280625 298578 280653 298606
rect 280687 298578 280715 298606
rect 280749 298578 280777 298606
rect 280811 298578 280839 298606
rect 280625 298516 280653 298544
rect 280687 298516 280715 298544
rect 280749 298516 280777 298544
rect 280811 298516 280839 298544
rect 280625 298454 280653 298482
rect 280687 298454 280715 298482
rect 280749 298454 280777 298482
rect 280811 298454 280839 298482
rect 280625 298392 280653 298420
rect 280687 298392 280715 298420
rect 280749 298392 280777 298420
rect 280811 298392 280839 298420
rect 280625 290147 280653 290175
rect 280687 290147 280715 290175
rect 280749 290147 280777 290175
rect 280811 290147 280839 290175
rect 280625 290085 280653 290113
rect 280687 290085 280715 290113
rect 280749 290085 280777 290113
rect 280811 290085 280839 290113
rect 280625 290023 280653 290051
rect 280687 290023 280715 290051
rect 280749 290023 280777 290051
rect 280811 290023 280839 290051
rect 280625 289961 280653 289989
rect 280687 289961 280715 289989
rect 280749 289961 280777 289989
rect 280811 289961 280839 289989
rect 280625 281147 280653 281175
rect 280687 281147 280715 281175
rect 280749 281147 280777 281175
rect 280811 281147 280839 281175
rect 280625 281085 280653 281113
rect 280687 281085 280715 281113
rect 280749 281085 280777 281113
rect 280811 281085 280839 281113
rect 280625 281023 280653 281051
rect 280687 281023 280715 281051
rect 280749 281023 280777 281051
rect 280811 281023 280839 281051
rect 280625 280961 280653 280989
rect 280687 280961 280715 280989
rect 280749 280961 280777 280989
rect 280811 280961 280839 280989
rect 280625 272147 280653 272175
rect 280687 272147 280715 272175
rect 280749 272147 280777 272175
rect 280811 272147 280839 272175
rect 280625 272085 280653 272113
rect 280687 272085 280715 272113
rect 280749 272085 280777 272113
rect 280811 272085 280839 272113
rect 280625 272023 280653 272051
rect 280687 272023 280715 272051
rect 280749 272023 280777 272051
rect 280811 272023 280839 272051
rect 280625 271961 280653 271989
rect 280687 271961 280715 271989
rect 280749 271961 280777 271989
rect 280811 271961 280839 271989
rect 280625 263147 280653 263175
rect 280687 263147 280715 263175
rect 280749 263147 280777 263175
rect 280811 263147 280839 263175
rect 280625 263085 280653 263113
rect 280687 263085 280715 263113
rect 280749 263085 280777 263113
rect 280811 263085 280839 263113
rect 280625 263023 280653 263051
rect 280687 263023 280715 263051
rect 280749 263023 280777 263051
rect 280811 263023 280839 263051
rect 280625 262961 280653 262989
rect 280687 262961 280715 262989
rect 280749 262961 280777 262989
rect 280811 262961 280839 262989
rect 280625 254147 280653 254175
rect 280687 254147 280715 254175
rect 280749 254147 280777 254175
rect 280811 254147 280839 254175
rect 280625 254085 280653 254113
rect 280687 254085 280715 254113
rect 280749 254085 280777 254113
rect 280811 254085 280839 254113
rect 280625 254023 280653 254051
rect 280687 254023 280715 254051
rect 280749 254023 280777 254051
rect 280811 254023 280839 254051
rect 280625 253961 280653 253989
rect 280687 253961 280715 253989
rect 280749 253961 280777 253989
rect 280811 253961 280839 253989
rect 280625 245147 280653 245175
rect 280687 245147 280715 245175
rect 280749 245147 280777 245175
rect 280811 245147 280839 245175
rect 280625 245085 280653 245113
rect 280687 245085 280715 245113
rect 280749 245085 280777 245113
rect 280811 245085 280839 245113
rect 280625 245023 280653 245051
rect 280687 245023 280715 245051
rect 280749 245023 280777 245051
rect 280811 245023 280839 245051
rect 280625 244961 280653 244989
rect 280687 244961 280715 244989
rect 280749 244961 280777 244989
rect 280811 244961 280839 244989
rect 280625 236147 280653 236175
rect 280687 236147 280715 236175
rect 280749 236147 280777 236175
rect 280811 236147 280839 236175
rect 280625 236085 280653 236113
rect 280687 236085 280715 236113
rect 280749 236085 280777 236113
rect 280811 236085 280839 236113
rect 280625 236023 280653 236051
rect 280687 236023 280715 236051
rect 280749 236023 280777 236051
rect 280811 236023 280839 236051
rect 280625 235961 280653 235989
rect 280687 235961 280715 235989
rect 280749 235961 280777 235989
rect 280811 235961 280839 235989
rect 280625 227147 280653 227175
rect 280687 227147 280715 227175
rect 280749 227147 280777 227175
rect 280811 227147 280839 227175
rect 280625 227085 280653 227113
rect 280687 227085 280715 227113
rect 280749 227085 280777 227113
rect 280811 227085 280839 227113
rect 280625 227023 280653 227051
rect 280687 227023 280715 227051
rect 280749 227023 280777 227051
rect 280811 227023 280839 227051
rect 280625 226961 280653 226989
rect 280687 226961 280715 226989
rect 280749 226961 280777 226989
rect 280811 226961 280839 226989
rect 280625 218147 280653 218175
rect 280687 218147 280715 218175
rect 280749 218147 280777 218175
rect 280811 218147 280839 218175
rect 280625 218085 280653 218113
rect 280687 218085 280715 218113
rect 280749 218085 280777 218113
rect 280811 218085 280839 218113
rect 280625 218023 280653 218051
rect 280687 218023 280715 218051
rect 280749 218023 280777 218051
rect 280811 218023 280839 218051
rect 280625 217961 280653 217989
rect 280687 217961 280715 217989
rect 280749 217961 280777 217989
rect 280811 217961 280839 217989
rect 280625 209147 280653 209175
rect 280687 209147 280715 209175
rect 280749 209147 280777 209175
rect 280811 209147 280839 209175
rect 280625 209085 280653 209113
rect 280687 209085 280715 209113
rect 280749 209085 280777 209113
rect 280811 209085 280839 209113
rect 280625 209023 280653 209051
rect 280687 209023 280715 209051
rect 280749 209023 280777 209051
rect 280811 209023 280839 209051
rect 280625 208961 280653 208989
rect 280687 208961 280715 208989
rect 280749 208961 280777 208989
rect 280811 208961 280839 208989
rect 280625 200147 280653 200175
rect 280687 200147 280715 200175
rect 280749 200147 280777 200175
rect 280811 200147 280839 200175
rect 280625 200085 280653 200113
rect 280687 200085 280715 200113
rect 280749 200085 280777 200113
rect 280811 200085 280839 200113
rect 280625 200023 280653 200051
rect 280687 200023 280715 200051
rect 280749 200023 280777 200051
rect 280811 200023 280839 200051
rect 280625 199961 280653 199989
rect 280687 199961 280715 199989
rect 280749 199961 280777 199989
rect 280811 199961 280839 199989
rect 280625 191147 280653 191175
rect 280687 191147 280715 191175
rect 280749 191147 280777 191175
rect 280811 191147 280839 191175
rect 280625 191085 280653 191113
rect 280687 191085 280715 191113
rect 280749 191085 280777 191113
rect 280811 191085 280839 191113
rect 280625 191023 280653 191051
rect 280687 191023 280715 191051
rect 280749 191023 280777 191051
rect 280811 191023 280839 191051
rect 280625 190961 280653 190989
rect 280687 190961 280715 190989
rect 280749 190961 280777 190989
rect 280811 190961 280839 190989
rect 280625 182147 280653 182175
rect 280687 182147 280715 182175
rect 280749 182147 280777 182175
rect 280811 182147 280839 182175
rect 280625 182085 280653 182113
rect 280687 182085 280715 182113
rect 280749 182085 280777 182113
rect 280811 182085 280839 182113
rect 280625 182023 280653 182051
rect 280687 182023 280715 182051
rect 280749 182023 280777 182051
rect 280811 182023 280839 182051
rect 280625 181961 280653 181989
rect 280687 181961 280715 181989
rect 280749 181961 280777 181989
rect 280811 181961 280839 181989
rect 280625 173147 280653 173175
rect 280687 173147 280715 173175
rect 280749 173147 280777 173175
rect 280811 173147 280839 173175
rect 280625 173085 280653 173113
rect 280687 173085 280715 173113
rect 280749 173085 280777 173113
rect 280811 173085 280839 173113
rect 280625 173023 280653 173051
rect 280687 173023 280715 173051
rect 280749 173023 280777 173051
rect 280811 173023 280839 173051
rect 280625 172961 280653 172989
rect 280687 172961 280715 172989
rect 280749 172961 280777 172989
rect 280811 172961 280839 172989
rect 280625 164147 280653 164175
rect 280687 164147 280715 164175
rect 280749 164147 280777 164175
rect 280811 164147 280839 164175
rect 280625 164085 280653 164113
rect 280687 164085 280715 164113
rect 280749 164085 280777 164113
rect 280811 164085 280839 164113
rect 280625 164023 280653 164051
rect 280687 164023 280715 164051
rect 280749 164023 280777 164051
rect 280811 164023 280839 164051
rect 280625 163961 280653 163989
rect 280687 163961 280715 163989
rect 280749 163961 280777 163989
rect 280811 163961 280839 163989
rect 280625 155147 280653 155175
rect 280687 155147 280715 155175
rect 280749 155147 280777 155175
rect 280811 155147 280839 155175
rect 280625 155085 280653 155113
rect 280687 155085 280715 155113
rect 280749 155085 280777 155113
rect 280811 155085 280839 155113
rect 280625 155023 280653 155051
rect 280687 155023 280715 155051
rect 280749 155023 280777 155051
rect 280811 155023 280839 155051
rect 280625 154961 280653 154989
rect 280687 154961 280715 154989
rect 280749 154961 280777 154989
rect 280811 154961 280839 154989
rect 280625 146147 280653 146175
rect 280687 146147 280715 146175
rect 280749 146147 280777 146175
rect 280811 146147 280839 146175
rect 280625 146085 280653 146113
rect 280687 146085 280715 146113
rect 280749 146085 280777 146113
rect 280811 146085 280839 146113
rect 280625 146023 280653 146051
rect 280687 146023 280715 146051
rect 280749 146023 280777 146051
rect 280811 146023 280839 146051
rect 280625 145961 280653 145989
rect 280687 145961 280715 145989
rect 280749 145961 280777 145989
rect 280811 145961 280839 145989
rect 280625 137147 280653 137175
rect 280687 137147 280715 137175
rect 280749 137147 280777 137175
rect 280811 137147 280839 137175
rect 280625 137085 280653 137113
rect 280687 137085 280715 137113
rect 280749 137085 280777 137113
rect 280811 137085 280839 137113
rect 280625 137023 280653 137051
rect 280687 137023 280715 137051
rect 280749 137023 280777 137051
rect 280811 137023 280839 137051
rect 280625 136961 280653 136989
rect 280687 136961 280715 136989
rect 280749 136961 280777 136989
rect 280811 136961 280839 136989
rect 280625 128147 280653 128175
rect 280687 128147 280715 128175
rect 280749 128147 280777 128175
rect 280811 128147 280839 128175
rect 280625 128085 280653 128113
rect 280687 128085 280715 128113
rect 280749 128085 280777 128113
rect 280811 128085 280839 128113
rect 280625 128023 280653 128051
rect 280687 128023 280715 128051
rect 280749 128023 280777 128051
rect 280811 128023 280839 128051
rect 280625 127961 280653 127989
rect 280687 127961 280715 127989
rect 280749 127961 280777 127989
rect 280811 127961 280839 127989
rect 280625 119147 280653 119175
rect 280687 119147 280715 119175
rect 280749 119147 280777 119175
rect 280811 119147 280839 119175
rect 280625 119085 280653 119113
rect 280687 119085 280715 119113
rect 280749 119085 280777 119113
rect 280811 119085 280839 119113
rect 280625 119023 280653 119051
rect 280687 119023 280715 119051
rect 280749 119023 280777 119051
rect 280811 119023 280839 119051
rect 280625 118961 280653 118989
rect 280687 118961 280715 118989
rect 280749 118961 280777 118989
rect 280811 118961 280839 118989
rect 280625 110147 280653 110175
rect 280687 110147 280715 110175
rect 280749 110147 280777 110175
rect 280811 110147 280839 110175
rect 280625 110085 280653 110113
rect 280687 110085 280715 110113
rect 280749 110085 280777 110113
rect 280811 110085 280839 110113
rect 280625 110023 280653 110051
rect 280687 110023 280715 110051
rect 280749 110023 280777 110051
rect 280811 110023 280839 110051
rect 280625 109961 280653 109989
rect 280687 109961 280715 109989
rect 280749 109961 280777 109989
rect 280811 109961 280839 109989
rect 280625 101147 280653 101175
rect 280687 101147 280715 101175
rect 280749 101147 280777 101175
rect 280811 101147 280839 101175
rect 280625 101085 280653 101113
rect 280687 101085 280715 101113
rect 280749 101085 280777 101113
rect 280811 101085 280839 101113
rect 280625 101023 280653 101051
rect 280687 101023 280715 101051
rect 280749 101023 280777 101051
rect 280811 101023 280839 101051
rect 280625 100961 280653 100989
rect 280687 100961 280715 100989
rect 280749 100961 280777 100989
rect 280811 100961 280839 100989
rect 280625 92147 280653 92175
rect 280687 92147 280715 92175
rect 280749 92147 280777 92175
rect 280811 92147 280839 92175
rect 280625 92085 280653 92113
rect 280687 92085 280715 92113
rect 280749 92085 280777 92113
rect 280811 92085 280839 92113
rect 280625 92023 280653 92051
rect 280687 92023 280715 92051
rect 280749 92023 280777 92051
rect 280811 92023 280839 92051
rect 280625 91961 280653 91989
rect 280687 91961 280715 91989
rect 280749 91961 280777 91989
rect 280811 91961 280839 91989
rect 280625 83147 280653 83175
rect 280687 83147 280715 83175
rect 280749 83147 280777 83175
rect 280811 83147 280839 83175
rect 280625 83085 280653 83113
rect 280687 83085 280715 83113
rect 280749 83085 280777 83113
rect 280811 83085 280839 83113
rect 280625 83023 280653 83051
rect 280687 83023 280715 83051
rect 280749 83023 280777 83051
rect 280811 83023 280839 83051
rect 280625 82961 280653 82989
rect 280687 82961 280715 82989
rect 280749 82961 280777 82989
rect 280811 82961 280839 82989
rect 280625 74147 280653 74175
rect 280687 74147 280715 74175
rect 280749 74147 280777 74175
rect 280811 74147 280839 74175
rect 280625 74085 280653 74113
rect 280687 74085 280715 74113
rect 280749 74085 280777 74113
rect 280811 74085 280839 74113
rect 280625 74023 280653 74051
rect 280687 74023 280715 74051
rect 280749 74023 280777 74051
rect 280811 74023 280839 74051
rect 280625 73961 280653 73989
rect 280687 73961 280715 73989
rect 280749 73961 280777 73989
rect 280811 73961 280839 73989
rect 280625 65147 280653 65175
rect 280687 65147 280715 65175
rect 280749 65147 280777 65175
rect 280811 65147 280839 65175
rect 280625 65085 280653 65113
rect 280687 65085 280715 65113
rect 280749 65085 280777 65113
rect 280811 65085 280839 65113
rect 280625 65023 280653 65051
rect 280687 65023 280715 65051
rect 280749 65023 280777 65051
rect 280811 65023 280839 65051
rect 280625 64961 280653 64989
rect 280687 64961 280715 64989
rect 280749 64961 280777 64989
rect 280811 64961 280839 64989
rect 280625 56147 280653 56175
rect 280687 56147 280715 56175
rect 280749 56147 280777 56175
rect 280811 56147 280839 56175
rect 280625 56085 280653 56113
rect 280687 56085 280715 56113
rect 280749 56085 280777 56113
rect 280811 56085 280839 56113
rect 280625 56023 280653 56051
rect 280687 56023 280715 56051
rect 280749 56023 280777 56051
rect 280811 56023 280839 56051
rect 280625 55961 280653 55989
rect 280687 55961 280715 55989
rect 280749 55961 280777 55989
rect 280811 55961 280839 55989
rect 280625 47147 280653 47175
rect 280687 47147 280715 47175
rect 280749 47147 280777 47175
rect 280811 47147 280839 47175
rect 280625 47085 280653 47113
rect 280687 47085 280715 47113
rect 280749 47085 280777 47113
rect 280811 47085 280839 47113
rect 280625 47023 280653 47051
rect 280687 47023 280715 47051
rect 280749 47023 280777 47051
rect 280811 47023 280839 47051
rect 280625 46961 280653 46989
rect 280687 46961 280715 46989
rect 280749 46961 280777 46989
rect 280811 46961 280839 46989
rect 280625 38147 280653 38175
rect 280687 38147 280715 38175
rect 280749 38147 280777 38175
rect 280811 38147 280839 38175
rect 280625 38085 280653 38113
rect 280687 38085 280715 38113
rect 280749 38085 280777 38113
rect 280811 38085 280839 38113
rect 280625 38023 280653 38051
rect 280687 38023 280715 38051
rect 280749 38023 280777 38051
rect 280811 38023 280839 38051
rect 280625 37961 280653 37989
rect 280687 37961 280715 37989
rect 280749 37961 280777 37989
rect 280811 37961 280839 37989
rect 280625 29147 280653 29175
rect 280687 29147 280715 29175
rect 280749 29147 280777 29175
rect 280811 29147 280839 29175
rect 280625 29085 280653 29113
rect 280687 29085 280715 29113
rect 280749 29085 280777 29113
rect 280811 29085 280839 29113
rect 280625 29023 280653 29051
rect 280687 29023 280715 29051
rect 280749 29023 280777 29051
rect 280811 29023 280839 29051
rect 280625 28961 280653 28989
rect 280687 28961 280715 28989
rect 280749 28961 280777 28989
rect 280811 28961 280839 28989
rect 280625 20147 280653 20175
rect 280687 20147 280715 20175
rect 280749 20147 280777 20175
rect 280811 20147 280839 20175
rect 280625 20085 280653 20113
rect 280687 20085 280715 20113
rect 280749 20085 280777 20113
rect 280811 20085 280839 20113
rect 280625 20023 280653 20051
rect 280687 20023 280715 20051
rect 280749 20023 280777 20051
rect 280811 20023 280839 20051
rect 280625 19961 280653 19989
rect 280687 19961 280715 19989
rect 280749 19961 280777 19989
rect 280811 19961 280839 19989
rect 280625 11147 280653 11175
rect 280687 11147 280715 11175
rect 280749 11147 280777 11175
rect 280811 11147 280839 11175
rect 280625 11085 280653 11113
rect 280687 11085 280715 11113
rect 280749 11085 280777 11113
rect 280811 11085 280839 11113
rect 280625 11023 280653 11051
rect 280687 11023 280715 11051
rect 280749 11023 280777 11051
rect 280811 11023 280839 11051
rect 280625 10961 280653 10989
rect 280687 10961 280715 10989
rect 280749 10961 280777 10989
rect 280811 10961 280839 10989
rect 280625 2147 280653 2175
rect 280687 2147 280715 2175
rect 280749 2147 280777 2175
rect 280811 2147 280839 2175
rect 280625 2085 280653 2113
rect 280687 2085 280715 2113
rect 280749 2085 280777 2113
rect 280811 2085 280839 2113
rect 280625 2023 280653 2051
rect 280687 2023 280715 2051
rect 280749 2023 280777 2051
rect 280811 2023 280839 2051
rect 280625 1961 280653 1989
rect 280687 1961 280715 1989
rect 280749 1961 280777 1989
rect 280811 1961 280839 1989
rect 280625 -108 280653 -80
rect 280687 -108 280715 -80
rect 280749 -108 280777 -80
rect 280811 -108 280839 -80
rect 280625 -170 280653 -142
rect 280687 -170 280715 -142
rect 280749 -170 280777 -142
rect 280811 -170 280839 -142
rect 280625 -232 280653 -204
rect 280687 -232 280715 -204
rect 280749 -232 280777 -204
rect 280811 -232 280839 -204
rect 280625 -294 280653 -266
rect 280687 -294 280715 -266
rect 280749 -294 280777 -266
rect 280811 -294 280839 -266
rect 282485 299058 282513 299086
rect 282547 299058 282575 299086
rect 282609 299058 282637 299086
rect 282671 299058 282699 299086
rect 282485 298996 282513 299024
rect 282547 298996 282575 299024
rect 282609 298996 282637 299024
rect 282671 298996 282699 299024
rect 282485 298934 282513 298962
rect 282547 298934 282575 298962
rect 282609 298934 282637 298962
rect 282671 298934 282699 298962
rect 282485 298872 282513 298900
rect 282547 298872 282575 298900
rect 282609 298872 282637 298900
rect 282671 298872 282699 298900
rect 282485 293147 282513 293175
rect 282547 293147 282575 293175
rect 282609 293147 282637 293175
rect 282671 293147 282699 293175
rect 282485 293085 282513 293113
rect 282547 293085 282575 293113
rect 282609 293085 282637 293113
rect 282671 293085 282699 293113
rect 282485 293023 282513 293051
rect 282547 293023 282575 293051
rect 282609 293023 282637 293051
rect 282671 293023 282699 293051
rect 282485 292961 282513 292989
rect 282547 292961 282575 292989
rect 282609 292961 282637 292989
rect 282671 292961 282699 292989
rect 282485 284147 282513 284175
rect 282547 284147 282575 284175
rect 282609 284147 282637 284175
rect 282671 284147 282699 284175
rect 282485 284085 282513 284113
rect 282547 284085 282575 284113
rect 282609 284085 282637 284113
rect 282671 284085 282699 284113
rect 282485 284023 282513 284051
rect 282547 284023 282575 284051
rect 282609 284023 282637 284051
rect 282671 284023 282699 284051
rect 282485 283961 282513 283989
rect 282547 283961 282575 283989
rect 282609 283961 282637 283989
rect 282671 283961 282699 283989
rect 282485 275147 282513 275175
rect 282547 275147 282575 275175
rect 282609 275147 282637 275175
rect 282671 275147 282699 275175
rect 282485 275085 282513 275113
rect 282547 275085 282575 275113
rect 282609 275085 282637 275113
rect 282671 275085 282699 275113
rect 282485 275023 282513 275051
rect 282547 275023 282575 275051
rect 282609 275023 282637 275051
rect 282671 275023 282699 275051
rect 282485 274961 282513 274989
rect 282547 274961 282575 274989
rect 282609 274961 282637 274989
rect 282671 274961 282699 274989
rect 282485 266147 282513 266175
rect 282547 266147 282575 266175
rect 282609 266147 282637 266175
rect 282671 266147 282699 266175
rect 282485 266085 282513 266113
rect 282547 266085 282575 266113
rect 282609 266085 282637 266113
rect 282671 266085 282699 266113
rect 282485 266023 282513 266051
rect 282547 266023 282575 266051
rect 282609 266023 282637 266051
rect 282671 266023 282699 266051
rect 282485 265961 282513 265989
rect 282547 265961 282575 265989
rect 282609 265961 282637 265989
rect 282671 265961 282699 265989
rect 282485 257147 282513 257175
rect 282547 257147 282575 257175
rect 282609 257147 282637 257175
rect 282671 257147 282699 257175
rect 282485 257085 282513 257113
rect 282547 257085 282575 257113
rect 282609 257085 282637 257113
rect 282671 257085 282699 257113
rect 282485 257023 282513 257051
rect 282547 257023 282575 257051
rect 282609 257023 282637 257051
rect 282671 257023 282699 257051
rect 282485 256961 282513 256989
rect 282547 256961 282575 256989
rect 282609 256961 282637 256989
rect 282671 256961 282699 256989
rect 282485 248147 282513 248175
rect 282547 248147 282575 248175
rect 282609 248147 282637 248175
rect 282671 248147 282699 248175
rect 282485 248085 282513 248113
rect 282547 248085 282575 248113
rect 282609 248085 282637 248113
rect 282671 248085 282699 248113
rect 282485 248023 282513 248051
rect 282547 248023 282575 248051
rect 282609 248023 282637 248051
rect 282671 248023 282699 248051
rect 282485 247961 282513 247989
rect 282547 247961 282575 247989
rect 282609 247961 282637 247989
rect 282671 247961 282699 247989
rect 282485 239147 282513 239175
rect 282547 239147 282575 239175
rect 282609 239147 282637 239175
rect 282671 239147 282699 239175
rect 282485 239085 282513 239113
rect 282547 239085 282575 239113
rect 282609 239085 282637 239113
rect 282671 239085 282699 239113
rect 282485 239023 282513 239051
rect 282547 239023 282575 239051
rect 282609 239023 282637 239051
rect 282671 239023 282699 239051
rect 282485 238961 282513 238989
rect 282547 238961 282575 238989
rect 282609 238961 282637 238989
rect 282671 238961 282699 238989
rect 282485 230147 282513 230175
rect 282547 230147 282575 230175
rect 282609 230147 282637 230175
rect 282671 230147 282699 230175
rect 282485 230085 282513 230113
rect 282547 230085 282575 230113
rect 282609 230085 282637 230113
rect 282671 230085 282699 230113
rect 282485 230023 282513 230051
rect 282547 230023 282575 230051
rect 282609 230023 282637 230051
rect 282671 230023 282699 230051
rect 282485 229961 282513 229989
rect 282547 229961 282575 229989
rect 282609 229961 282637 229989
rect 282671 229961 282699 229989
rect 282485 221147 282513 221175
rect 282547 221147 282575 221175
rect 282609 221147 282637 221175
rect 282671 221147 282699 221175
rect 282485 221085 282513 221113
rect 282547 221085 282575 221113
rect 282609 221085 282637 221113
rect 282671 221085 282699 221113
rect 282485 221023 282513 221051
rect 282547 221023 282575 221051
rect 282609 221023 282637 221051
rect 282671 221023 282699 221051
rect 282485 220961 282513 220989
rect 282547 220961 282575 220989
rect 282609 220961 282637 220989
rect 282671 220961 282699 220989
rect 282485 212147 282513 212175
rect 282547 212147 282575 212175
rect 282609 212147 282637 212175
rect 282671 212147 282699 212175
rect 282485 212085 282513 212113
rect 282547 212085 282575 212113
rect 282609 212085 282637 212113
rect 282671 212085 282699 212113
rect 282485 212023 282513 212051
rect 282547 212023 282575 212051
rect 282609 212023 282637 212051
rect 282671 212023 282699 212051
rect 282485 211961 282513 211989
rect 282547 211961 282575 211989
rect 282609 211961 282637 211989
rect 282671 211961 282699 211989
rect 282485 203147 282513 203175
rect 282547 203147 282575 203175
rect 282609 203147 282637 203175
rect 282671 203147 282699 203175
rect 282485 203085 282513 203113
rect 282547 203085 282575 203113
rect 282609 203085 282637 203113
rect 282671 203085 282699 203113
rect 282485 203023 282513 203051
rect 282547 203023 282575 203051
rect 282609 203023 282637 203051
rect 282671 203023 282699 203051
rect 282485 202961 282513 202989
rect 282547 202961 282575 202989
rect 282609 202961 282637 202989
rect 282671 202961 282699 202989
rect 282485 194147 282513 194175
rect 282547 194147 282575 194175
rect 282609 194147 282637 194175
rect 282671 194147 282699 194175
rect 282485 194085 282513 194113
rect 282547 194085 282575 194113
rect 282609 194085 282637 194113
rect 282671 194085 282699 194113
rect 282485 194023 282513 194051
rect 282547 194023 282575 194051
rect 282609 194023 282637 194051
rect 282671 194023 282699 194051
rect 282485 193961 282513 193989
rect 282547 193961 282575 193989
rect 282609 193961 282637 193989
rect 282671 193961 282699 193989
rect 282485 185147 282513 185175
rect 282547 185147 282575 185175
rect 282609 185147 282637 185175
rect 282671 185147 282699 185175
rect 282485 185085 282513 185113
rect 282547 185085 282575 185113
rect 282609 185085 282637 185113
rect 282671 185085 282699 185113
rect 282485 185023 282513 185051
rect 282547 185023 282575 185051
rect 282609 185023 282637 185051
rect 282671 185023 282699 185051
rect 282485 184961 282513 184989
rect 282547 184961 282575 184989
rect 282609 184961 282637 184989
rect 282671 184961 282699 184989
rect 282485 176147 282513 176175
rect 282547 176147 282575 176175
rect 282609 176147 282637 176175
rect 282671 176147 282699 176175
rect 282485 176085 282513 176113
rect 282547 176085 282575 176113
rect 282609 176085 282637 176113
rect 282671 176085 282699 176113
rect 282485 176023 282513 176051
rect 282547 176023 282575 176051
rect 282609 176023 282637 176051
rect 282671 176023 282699 176051
rect 282485 175961 282513 175989
rect 282547 175961 282575 175989
rect 282609 175961 282637 175989
rect 282671 175961 282699 175989
rect 282485 167147 282513 167175
rect 282547 167147 282575 167175
rect 282609 167147 282637 167175
rect 282671 167147 282699 167175
rect 282485 167085 282513 167113
rect 282547 167085 282575 167113
rect 282609 167085 282637 167113
rect 282671 167085 282699 167113
rect 282485 167023 282513 167051
rect 282547 167023 282575 167051
rect 282609 167023 282637 167051
rect 282671 167023 282699 167051
rect 282485 166961 282513 166989
rect 282547 166961 282575 166989
rect 282609 166961 282637 166989
rect 282671 166961 282699 166989
rect 282485 158147 282513 158175
rect 282547 158147 282575 158175
rect 282609 158147 282637 158175
rect 282671 158147 282699 158175
rect 282485 158085 282513 158113
rect 282547 158085 282575 158113
rect 282609 158085 282637 158113
rect 282671 158085 282699 158113
rect 282485 158023 282513 158051
rect 282547 158023 282575 158051
rect 282609 158023 282637 158051
rect 282671 158023 282699 158051
rect 282485 157961 282513 157989
rect 282547 157961 282575 157989
rect 282609 157961 282637 157989
rect 282671 157961 282699 157989
rect 282485 149147 282513 149175
rect 282547 149147 282575 149175
rect 282609 149147 282637 149175
rect 282671 149147 282699 149175
rect 282485 149085 282513 149113
rect 282547 149085 282575 149113
rect 282609 149085 282637 149113
rect 282671 149085 282699 149113
rect 282485 149023 282513 149051
rect 282547 149023 282575 149051
rect 282609 149023 282637 149051
rect 282671 149023 282699 149051
rect 282485 148961 282513 148989
rect 282547 148961 282575 148989
rect 282609 148961 282637 148989
rect 282671 148961 282699 148989
rect 282485 140147 282513 140175
rect 282547 140147 282575 140175
rect 282609 140147 282637 140175
rect 282671 140147 282699 140175
rect 282485 140085 282513 140113
rect 282547 140085 282575 140113
rect 282609 140085 282637 140113
rect 282671 140085 282699 140113
rect 282485 140023 282513 140051
rect 282547 140023 282575 140051
rect 282609 140023 282637 140051
rect 282671 140023 282699 140051
rect 282485 139961 282513 139989
rect 282547 139961 282575 139989
rect 282609 139961 282637 139989
rect 282671 139961 282699 139989
rect 282485 131147 282513 131175
rect 282547 131147 282575 131175
rect 282609 131147 282637 131175
rect 282671 131147 282699 131175
rect 282485 131085 282513 131113
rect 282547 131085 282575 131113
rect 282609 131085 282637 131113
rect 282671 131085 282699 131113
rect 282485 131023 282513 131051
rect 282547 131023 282575 131051
rect 282609 131023 282637 131051
rect 282671 131023 282699 131051
rect 282485 130961 282513 130989
rect 282547 130961 282575 130989
rect 282609 130961 282637 130989
rect 282671 130961 282699 130989
rect 282485 122147 282513 122175
rect 282547 122147 282575 122175
rect 282609 122147 282637 122175
rect 282671 122147 282699 122175
rect 282485 122085 282513 122113
rect 282547 122085 282575 122113
rect 282609 122085 282637 122113
rect 282671 122085 282699 122113
rect 282485 122023 282513 122051
rect 282547 122023 282575 122051
rect 282609 122023 282637 122051
rect 282671 122023 282699 122051
rect 282485 121961 282513 121989
rect 282547 121961 282575 121989
rect 282609 121961 282637 121989
rect 282671 121961 282699 121989
rect 282485 113147 282513 113175
rect 282547 113147 282575 113175
rect 282609 113147 282637 113175
rect 282671 113147 282699 113175
rect 282485 113085 282513 113113
rect 282547 113085 282575 113113
rect 282609 113085 282637 113113
rect 282671 113085 282699 113113
rect 282485 113023 282513 113051
rect 282547 113023 282575 113051
rect 282609 113023 282637 113051
rect 282671 113023 282699 113051
rect 282485 112961 282513 112989
rect 282547 112961 282575 112989
rect 282609 112961 282637 112989
rect 282671 112961 282699 112989
rect 282485 104147 282513 104175
rect 282547 104147 282575 104175
rect 282609 104147 282637 104175
rect 282671 104147 282699 104175
rect 282485 104085 282513 104113
rect 282547 104085 282575 104113
rect 282609 104085 282637 104113
rect 282671 104085 282699 104113
rect 282485 104023 282513 104051
rect 282547 104023 282575 104051
rect 282609 104023 282637 104051
rect 282671 104023 282699 104051
rect 282485 103961 282513 103989
rect 282547 103961 282575 103989
rect 282609 103961 282637 103989
rect 282671 103961 282699 103989
rect 282485 95147 282513 95175
rect 282547 95147 282575 95175
rect 282609 95147 282637 95175
rect 282671 95147 282699 95175
rect 282485 95085 282513 95113
rect 282547 95085 282575 95113
rect 282609 95085 282637 95113
rect 282671 95085 282699 95113
rect 282485 95023 282513 95051
rect 282547 95023 282575 95051
rect 282609 95023 282637 95051
rect 282671 95023 282699 95051
rect 282485 94961 282513 94989
rect 282547 94961 282575 94989
rect 282609 94961 282637 94989
rect 282671 94961 282699 94989
rect 282485 86147 282513 86175
rect 282547 86147 282575 86175
rect 282609 86147 282637 86175
rect 282671 86147 282699 86175
rect 282485 86085 282513 86113
rect 282547 86085 282575 86113
rect 282609 86085 282637 86113
rect 282671 86085 282699 86113
rect 282485 86023 282513 86051
rect 282547 86023 282575 86051
rect 282609 86023 282637 86051
rect 282671 86023 282699 86051
rect 282485 85961 282513 85989
rect 282547 85961 282575 85989
rect 282609 85961 282637 85989
rect 282671 85961 282699 85989
rect 282485 77147 282513 77175
rect 282547 77147 282575 77175
rect 282609 77147 282637 77175
rect 282671 77147 282699 77175
rect 282485 77085 282513 77113
rect 282547 77085 282575 77113
rect 282609 77085 282637 77113
rect 282671 77085 282699 77113
rect 282485 77023 282513 77051
rect 282547 77023 282575 77051
rect 282609 77023 282637 77051
rect 282671 77023 282699 77051
rect 282485 76961 282513 76989
rect 282547 76961 282575 76989
rect 282609 76961 282637 76989
rect 282671 76961 282699 76989
rect 282485 68147 282513 68175
rect 282547 68147 282575 68175
rect 282609 68147 282637 68175
rect 282671 68147 282699 68175
rect 282485 68085 282513 68113
rect 282547 68085 282575 68113
rect 282609 68085 282637 68113
rect 282671 68085 282699 68113
rect 282485 68023 282513 68051
rect 282547 68023 282575 68051
rect 282609 68023 282637 68051
rect 282671 68023 282699 68051
rect 282485 67961 282513 67989
rect 282547 67961 282575 67989
rect 282609 67961 282637 67989
rect 282671 67961 282699 67989
rect 282485 59147 282513 59175
rect 282547 59147 282575 59175
rect 282609 59147 282637 59175
rect 282671 59147 282699 59175
rect 282485 59085 282513 59113
rect 282547 59085 282575 59113
rect 282609 59085 282637 59113
rect 282671 59085 282699 59113
rect 282485 59023 282513 59051
rect 282547 59023 282575 59051
rect 282609 59023 282637 59051
rect 282671 59023 282699 59051
rect 282485 58961 282513 58989
rect 282547 58961 282575 58989
rect 282609 58961 282637 58989
rect 282671 58961 282699 58989
rect 282485 50147 282513 50175
rect 282547 50147 282575 50175
rect 282609 50147 282637 50175
rect 282671 50147 282699 50175
rect 282485 50085 282513 50113
rect 282547 50085 282575 50113
rect 282609 50085 282637 50113
rect 282671 50085 282699 50113
rect 282485 50023 282513 50051
rect 282547 50023 282575 50051
rect 282609 50023 282637 50051
rect 282671 50023 282699 50051
rect 282485 49961 282513 49989
rect 282547 49961 282575 49989
rect 282609 49961 282637 49989
rect 282671 49961 282699 49989
rect 282485 41147 282513 41175
rect 282547 41147 282575 41175
rect 282609 41147 282637 41175
rect 282671 41147 282699 41175
rect 282485 41085 282513 41113
rect 282547 41085 282575 41113
rect 282609 41085 282637 41113
rect 282671 41085 282699 41113
rect 282485 41023 282513 41051
rect 282547 41023 282575 41051
rect 282609 41023 282637 41051
rect 282671 41023 282699 41051
rect 282485 40961 282513 40989
rect 282547 40961 282575 40989
rect 282609 40961 282637 40989
rect 282671 40961 282699 40989
rect 282485 32147 282513 32175
rect 282547 32147 282575 32175
rect 282609 32147 282637 32175
rect 282671 32147 282699 32175
rect 282485 32085 282513 32113
rect 282547 32085 282575 32113
rect 282609 32085 282637 32113
rect 282671 32085 282699 32113
rect 282485 32023 282513 32051
rect 282547 32023 282575 32051
rect 282609 32023 282637 32051
rect 282671 32023 282699 32051
rect 282485 31961 282513 31989
rect 282547 31961 282575 31989
rect 282609 31961 282637 31989
rect 282671 31961 282699 31989
rect 282485 23147 282513 23175
rect 282547 23147 282575 23175
rect 282609 23147 282637 23175
rect 282671 23147 282699 23175
rect 282485 23085 282513 23113
rect 282547 23085 282575 23113
rect 282609 23085 282637 23113
rect 282671 23085 282699 23113
rect 282485 23023 282513 23051
rect 282547 23023 282575 23051
rect 282609 23023 282637 23051
rect 282671 23023 282699 23051
rect 282485 22961 282513 22989
rect 282547 22961 282575 22989
rect 282609 22961 282637 22989
rect 282671 22961 282699 22989
rect 282485 14147 282513 14175
rect 282547 14147 282575 14175
rect 282609 14147 282637 14175
rect 282671 14147 282699 14175
rect 282485 14085 282513 14113
rect 282547 14085 282575 14113
rect 282609 14085 282637 14113
rect 282671 14085 282699 14113
rect 282485 14023 282513 14051
rect 282547 14023 282575 14051
rect 282609 14023 282637 14051
rect 282671 14023 282699 14051
rect 282485 13961 282513 13989
rect 282547 13961 282575 13989
rect 282609 13961 282637 13989
rect 282671 13961 282699 13989
rect 282485 5147 282513 5175
rect 282547 5147 282575 5175
rect 282609 5147 282637 5175
rect 282671 5147 282699 5175
rect 282485 5085 282513 5113
rect 282547 5085 282575 5113
rect 282609 5085 282637 5113
rect 282671 5085 282699 5113
rect 282485 5023 282513 5051
rect 282547 5023 282575 5051
rect 282609 5023 282637 5051
rect 282671 5023 282699 5051
rect 282485 4961 282513 4989
rect 282547 4961 282575 4989
rect 282609 4961 282637 4989
rect 282671 4961 282699 4989
rect 282485 -588 282513 -560
rect 282547 -588 282575 -560
rect 282609 -588 282637 -560
rect 282671 -588 282699 -560
rect 282485 -650 282513 -622
rect 282547 -650 282575 -622
rect 282609 -650 282637 -622
rect 282671 -650 282699 -622
rect 282485 -712 282513 -684
rect 282547 -712 282575 -684
rect 282609 -712 282637 -684
rect 282671 -712 282699 -684
rect 282485 -774 282513 -746
rect 282547 -774 282575 -746
rect 282609 -774 282637 -746
rect 282671 -774 282699 -746
rect 289625 298578 289653 298606
rect 289687 298578 289715 298606
rect 289749 298578 289777 298606
rect 289811 298578 289839 298606
rect 289625 298516 289653 298544
rect 289687 298516 289715 298544
rect 289749 298516 289777 298544
rect 289811 298516 289839 298544
rect 289625 298454 289653 298482
rect 289687 298454 289715 298482
rect 289749 298454 289777 298482
rect 289811 298454 289839 298482
rect 289625 298392 289653 298420
rect 289687 298392 289715 298420
rect 289749 298392 289777 298420
rect 289811 298392 289839 298420
rect 289625 290147 289653 290175
rect 289687 290147 289715 290175
rect 289749 290147 289777 290175
rect 289811 290147 289839 290175
rect 289625 290085 289653 290113
rect 289687 290085 289715 290113
rect 289749 290085 289777 290113
rect 289811 290085 289839 290113
rect 289625 290023 289653 290051
rect 289687 290023 289715 290051
rect 289749 290023 289777 290051
rect 289811 290023 289839 290051
rect 289625 289961 289653 289989
rect 289687 289961 289715 289989
rect 289749 289961 289777 289989
rect 289811 289961 289839 289989
rect 289625 281147 289653 281175
rect 289687 281147 289715 281175
rect 289749 281147 289777 281175
rect 289811 281147 289839 281175
rect 289625 281085 289653 281113
rect 289687 281085 289715 281113
rect 289749 281085 289777 281113
rect 289811 281085 289839 281113
rect 289625 281023 289653 281051
rect 289687 281023 289715 281051
rect 289749 281023 289777 281051
rect 289811 281023 289839 281051
rect 289625 280961 289653 280989
rect 289687 280961 289715 280989
rect 289749 280961 289777 280989
rect 289811 280961 289839 280989
rect 289625 272147 289653 272175
rect 289687 272147 289715 272175
rect 289749 272147 289777 272175
rect 289811 272147 289839 272175
rect 289625 272085 289653 272113
rect 289687 272085 289715 272113
rect 289749 272085 289777 272113
rect 289811 272085 289839 272113
rect 289625 272023 289653 272051
rect 289687 272023 289715 272051
rect 289749 272023 289777 272051
rect 289811 272023 289839 272051
rect 289625 271961 289653 271989
rect 289687 271961 289715 271989
rect 289749 271961 289777 271989
rect 289811 271961 289839 271989
rect 289625 263147 289653 263175
rect 289687 263147 289715 263175
rect 289749 263147 289777 263175
rect 289811 263147 289839 263175
rect 289625 263085 289653 263113
rect 289687 263085 289715 263113
rect 289749 263085 289777 263113
rect 289811 263085 289839 263113
rect 289625 263023 289653 263051
rect 289687 263023 289715 263051
rect 289749 263023 289777 263051
rect 289811 263023 289839 263051
rect 289625 262961 289653 262989
rect 289687 262961 289715 262989
rect 289749 262961 289777 262989
rect 289811 262961 289839 262989
rect 289625 254147 289653 254175
rect 289687 254147 289715 254175
rect 289749 254147 289777 254175
rect 289811 254147 289839 254175
rect 289625 254085 289653 254113
rect 289687 254085 289715 254113
rect 289749 254085 289777 254113
rect 289811 254085 289839 254113
rect 289625 254023 289653 254051
rect 289687 254023 289715 254051
rect 289749 254023 289777 254051
rect 289811 254023 289839 254051
rect 289625 253961 289653 253989
rect 289687 253961 289715 253989
rect 289749 253961 289777 253989
rect 289811 253961 289839 253989
rect 289625 245147 289653 245175
rect 289687 245147 289715 245175
rect 289749 245147 289777 245175
rect 289811 245147 289839 245175
rect 289625 245085 289653 245113
rect 289687 245085 289715 245113
rect 289749 245085 289777 245113
rect 289811 245085 289839 245113
rect 289625 245023 289653 245051
rect 289687 245023 289715 245051
rect 289749 245023 289777 245051
rect 289811 245023 289839 245051
rect 289625 244961 289653 244989
rect 289687 244961 289715 244989
rect 289749 244961 289777 244989
rect 289811 244961 289839 244989
rect 289625 236147 289653 236175
rect 289687 236147 289715 236175
rect 289749 236147 289777 236175
rect 289811 236147 289839 236175
rect 289625 236085 289653 236113
rect 289687 236085 289715 236113
rect 289749 236085 289777 236113
rect 289811 236085 289839 236113
rect 289625 236023 289653 236051
rect 289687 236023 289715 236051
rect 289749 236023 289777 236051
rect 289811 236023 289839 236051
rect 289625 235961 289653 235989
rect 289687 235961 289715 235989
rect 289749 235961 289777 235989
rect 289811 235961 289839 235989
rect 289625 227147 289653 227175
rect 289687 227147 289715 227175
rect 289749 227147 289777 227175
rect 289811 227147 289839 227175
rect 289625 227085 289653 227113
rect 289687 227085 289715 227113
rect 289749 227085 289777 227113
rect 289811 227085 289839 227113
rect 289625 227023 289653 227051
rect 289687 227023 289715 227051
rect 289749 227023 289777 227051
rect 289811 227023 289839 227051
rect 289625 226961 289653 226989
rect 289687 226961 289715 226989
rect 289749 226961 289777 226989
rect 289811 226961 289839 226989
rect 289625 218147 289653 218175
rect 289687 218147 289715 218175
rect 289749 218147 289777 218175
rect 289811 218147 289839 218175
rect 289625 218085 289653 218113
rect 289687 218085 289715 218113
rect 289749 218085 289777 218113
rect 289811 218085 289839 218113
rect 289625 218023 289653 218051
rect 289687 218023 289715 218051
rect 289749 218023 289777 218051
rect 289811 218023 289839 218051
rect 289625 217961 289653 217989
rect 289687 217961 289715 217989
rect 289749 217961 289777 217989
rect 289811 217961 289839 217989
rect 289625 209147 289653 209175
rect 289687 209147 289715 209175
rect 289749 209147 289777 209175
rect 289811 209147 289839 209175
rect 289625 209085 289653 209113
rect 289687 209085 289715 209113
rect 289749 209085 289777 209113
rect 289811 209085 289839 209113
rect 289625 209023 289653 209051
rect 289687 209023 289715 209051
rect 289749 209023 289777 209051
rect 289811 209023 289839 209051
rect 289625 208961 289653 208989
rect 289687 208961 289715 208989
rect 289749 208961 289777 208989
rect 289811 208961 289839 208989
rect 289625 200147 289653 200175
rect 289687 200147 289715 200175
rect 289749 200147 289777 200175
rect 289811 200147 289839 200175
rect 289625 200085 289653 200113
rect 289687 200085 289715 200113
rect 289749 200085 289777 200113
rect 289811 200085 289839 200113
rect 289625 200023 289653 200051
rect 289687 200023 289715 200051
rect 289749 200023 289777 200051
rect 289811 200023 289839 200051
rect 289625 199961 289653 199989
rect 289687 199961 289715 199989
rect 289749 199961 289777 199989
rect 289811 199961 289839 199989
rect 289625 191147 289653 191175
rect 289687 191147 289715 191175
rect 289749 191147 289777 191175
rect 289811 191147 289839 191175
rect 289625 191085 289653 191113
rect 289687 191085 289715 191113
rect 289749 191085 289777 191113
rect 289811 191085 289839 191113
rect 289625 191023 289653 191051
rect 289687 191023 289715 191051
rect 289749 191023 289777 191051
rect 289811 191023 289839 191051
rect 289625 190961 289653 190989
rect 289687 190961 289715 190989
rect 289749 190961 289777 190989
rect 289811 190961 289839 190989
rect 289625 182147 289653 182175
rect 289687 182147 289715 182175
rect 289749 182147 289777 182175
rect 289811 182147 289839 182175
rect 289625 182085 289653 182113
rect 289687 182085 289715 182113
rect 289749 182085 289777 182113
rect 289811 182085 289839 182113
rect 289625 182023 289653 182051
rect 289687 182023 289715 182051
rect 289749 182023 289777 182051
rect 289811 182023 289839 182051
rect 289625 181961 289653 181989
rect 289687 181961 289715 181989
rect 289749 181961 289777 181989
rect 289811 181961 289839 181989
rect 289625 173147 289653 173175
rect 289687 173147 289715 173175
rect 289749 173147 289777 173175
rect 289811 173147 289839 173175
rect 289625 173085 289653 173113
rect 289687 173085 289715 173113
rect 289749 173085 289777 173113
rect 289811 173085 289839 173113
rect 289625 173023 289653 173051
rect 289687 173023 289715 173051
rect 289749 173023 289777 173051
rect 289811 173023 289839 173051
rect 289625 172961 289653 172989
rect 289687 172961 289715 172989
rect 289749 172961 289777 172989
rect 289811 172961 289839 172989
rect 289625 164147 289653 164175
rect 289687 164147 289715 164175
rect 289749 164147 289777 164175
rect 289811 164147 289839 164175
rect 289625 164085 289653 164113
rect 289687 164085 289715 164113
rect 289749 164085 289777 164113
rect 289811 164085 289839 164113
rect 289625 164023 289653 164051
rect 289687 164023 289715 164051
rect 289749 164023 289777 164051
rect 289811 164023 289839 164051
rect 289625 163961 289653 163989
rect 289687 163961 289715 163989
rect 289749 163961 289777 163989
rect 289811 163961 289839 163989
rect 289625 155147 289653 155175
rect 289687 155147 289715 155175
rect 289749 155147 289777 155175
rect 289811 155147 289839 155175
rect 289625 155085 289653 155113
rect 289687 155085 289715 155113
rect 289749 155085 289777 155113
rect 289811 155085 289839 155113
rect 289625 155023 289653 155051
rect 289687 155023 289715 155051
rect 289749 155023 289777 155051
rect 289811 155023 289839 155051
rect 289625 154961 289653 154989
rect 289687 154961 289715 154989
rect 289749 154961 289777 154989
rect 289811 154961 289839 154989
rect 289625 146147 289653 146175
rect 289687 146147 289715 146175
rect 289749 146147 289777 146175
rect 289811 146147 289839 146175
rect 289625 146085 289653 146113
rect 289687 146085 289715 146113
rect 289749 146085 289777 146113
rect 289811 146085 289839 146113
rect 289625 146023 289653 146051
rect 289687 146023 289715 146051
rect 289749 146023 289777 146051
rect 289811 146023 289839 146051
rect 289625 145961 289653 145989
rect 289687 145961 289715 145989
rect 289749 145961 289777 145989
rect 289811 145961 289839 145989
rect 289625 137147 289653 137175
rect 289687 137147 289715 137175
rect 289749 137147 289777 137175
rect 289811 137147 289839 137175
rect 289625 137085 289653 137113
rect 289687 137085 289715 137113
rect 289749 137085 289777 137113
rect 289811 137085 289839 137113
rect 289625 137023 289653 137051
rect 289687 137023 289715 137051
rect 289749 137023 289777 137051
rect 289811 137023 289839 137051
rect 289625 136961 289653 136989
rect 289687 136961 289715 136989
rect 289749 136961 289777 136989
rect 289811 136961 289839 136989
rect 289625 128147 289653 128175
rect 289687 128147 289715 128175
rect 289749 128147 289777 128175
rect 289811 128147 289839 128175
rect 289625 128085 289653 128113
rect 289687 128085 289715 128113
rect 289749 128085 289777 128113
rect 289811 128085 289839 128113
rect 289625 128023 289653 128051
rect 289687 128023 289715 128051
rect 289749 128023 289777 128051
rect 289811 128023 289839 128051
rect 289625 127961 289653 127989
rect 289687 127961 289715 127989
rect 289749 127961 289777 127989
rect 289811 127961 289839 127989
rect 289625 119147 289653 119175
rect 289687 119147 289715 119175
rect 289749 119147 289777 119175
rect 289811 119147 289839 119175
rect 289625 119085 289653 119113
rect 289687 119085 289715 119113
rect 289749 119085 289777 119113
rect 289811 119085 289839 119113
rect 289625 119023 289653 119051
rect 289687 119023 289715 119051
rect 289749 119023 289777 119051
rect 289811 119023 289839 119051
rect 289625 118961 289653 118989
rect 289687 118961 289715 118989
rect 289749 118961 289777 118989
rect 289811 118961 289839 118989
rect 289625 110147 289653 110175
rect 289687 110147 289715 110175
rect 289749 110147 289777 110175
rect 289811 110147 289839 110175
rect 289625 110085 289653 110113
rect 289687 110085 289715 110113
rect 289749 110085 289777 110113
rect 289811 110085 289839 110113
rect 289625 110023 289653 110051
rect 289687 110023 289715 110051
rect 289749 110023 289777 110051
rect 289811 110023 289839 110051
rect 289625 109961 289653 109989
rect 289687 109961 289715 109989
rect 289749 109961 289777 109989
rect 289811 109961 289839 109989
rect 289625 101147 289653 101175
rect 289687 101147 289715 101175
rect 289749 101147 289777 101175
rect 289811 101147 289839 101175
rect 289625 101085 289653 101113
rect 289687 101085 289715 101113
rect 289749 101085 289777 101113
rect 289811 101085 289839 101113
rect 289625 101023 289653 101051
rect 289687 101023 289715 101051
rect 289749 101023 289777 101051
rect 289811 101023 289839 101051
rect 289625 100961 289653 100989
rect 289687 100961 289715 100989
rect 289749 100961 289777 100989
rect 289811 100961 289839 100989
rect 289625 92147 289653 92175
rect 289687 92147 289715 92175
rect 289749 92147 289777 92175
rect 289811 92147 289839 92175
rect 289625 92085 289653 92113
rect 289687 92085 289715 92113
rect 289749 92085 289777 92113
rect 289811 92085 289839 92113
rect 289625 92023 289653 92051
rect 289687 92023 289715 92051
rect 289749 92023 289777 92051
rect 289811 92023 289839 92051
rect 289625 91961 289653 91989
rect 289687 91961 289715 91989
rect 289749 91961 289777 91989
rect 289811 91961 289839 91989
rect 289625 83147 289653 83175
rect 289687 83147 289715 83175
rect 289749 83147 289777 83175
rect 289811 83147 289839 83175
rect 289625 83085 289653 83113
rect 289687 83085 289715 83113
rect 289749 83085 289777 83113
rect 289811 83085 289839 83113
rect 289625 83023 289653 83051
rect 289687 83023 289715 83051
rect 289749 83023 289777 83051
rect 289811 83023 289839 83051
rect 289625 82961 289653 82989
rect 289687 82961 289715 82989
rect 289749 82961 289777 82989
rect 289811 82961 289839 82989
rect 289625 74147 289653 74175
rect 289687 74147 289715 74175
rect 289749 74147 289777 74175
rect 289811 74147 289839 74175
rect 289625 74085 289653 74113
rect 289687 74085 289715 74113
rect 289749 74085 289777 74113
rect 289811 74085 289839 74113
rect 289625 74023 289653 74051
rect 289687 74023 289715 74051
rect 289749 74023 289777 74051
rect 289811 74023 289839 74051
rect 289625 73961 289653 73989
rect 289687 73961 289715 73989
rect 289749 73961 289777 73989
rect 289811 73961 289839 73989
rect 289625 65147 289653 65175
rect 289687 65147 289715 65175
rect 289749 65147 289777 65175
rect 289811 65147 289839 65175
rect 289625 65085 289653 65113
rect 289687 65085 289715 65113
rect 289749 65085 289777 65113
rect 289811 65085 289839 65113
rect 289625 65023 289653 65051
rect 289687 65023 289715 65051
rect 289749 65023 289777 65051
rect 289811 65023 289839 65051
rect 289625 64961 289653 64989
rect 289687 64961 289715 64989
rect 289749 64961 289777 64989
rect 289811 64961 289839 64989
rect 289625 56147 289653 56175
rect 289687 56147 289715 56175
rect 289749 56147 289777 56175
rect 289811 56147 289839 56175
rect 289625 56085 289653 56113
rect 289687 56085 289715 56113
rect 289749 56085 289777 56113
rect 289811 56085 289839 56113
rect 289625 56023 289653 56051
rect 289687 56023 289715 56051
rect 289749 56023 289777 56051
rect 289811 56023 289839 56051
rect 289625 55961 289653 55989
rect 289687 55961 289715 55989
rect 289749 55961 289777 55989
rect 289811 55961 289839 55989
rect 289625 47147 289653 47175
rect 289687 47147 289715 47175
rect 289749 47147 289777 47175
rect 289811 47147 289839 47175
rect 289625 47085 289653 47113
rect 289687 47085 289715 47113
rect 289749 47085 289777 47113
rect 289811 47085 289839 47113
rect 289625 47023 289653 47051
rect 289687 47023 289715 47051
rect 289749 47023 289777 47051
rect 289811 47023 289839 47051
rect 289625 46961 289653 46989
rect 289687 46961 289715 46989
rect 289749 46961 289777 46989
rect 289811 46961 289839 46989
rect 289625 38147 289653 38175
rect 289687 38147 289715 38175
rect 289749 38147 289777 38175
rect 289811 38147 289839 38175
rect 289625 38085 289653 38113
rect 289687 38085 289715 38113
rect 289749 38085 289777 38113
rect 289811 38085 289839 38113
rect 289625 38023 289653 38051
rect 289687 38023 289715 38051
rect 289749 38023 289777 38051
rect 289811 38023 289839 38051
rect 289625 37961 289653 37989
rect 289687 37961 289715 37989
rect 289749 37961 289777 37989
rect 289811 37961 289839 37989
rect 289625 29147 289653 29175
rect 289687 29147 289715 29175
rect 289749 29147 289777 29175
rect 289811 29147 289839 29175
rect 289625 29085 289653 29113
rect 289687 29085 289715 29113
rect 289749 29085 289777 29113
rect 289811 29085 289839 29113
rect 289625 29023 289653 29051
rect 289687 29023 289715 29051
rect 289749 29023 289777 29051
rect 289811 29023 289839 29051
rect 289625 28961 289653 28989
rect 289687 28961 289715 28989
rect 289749 28961 289777 28989
rect 289811 28961 289839 28989
rect 289625 20147 289653 20175
rect 289687 20147 289715 20175
rect 289749 20147 289777 20175
rect 289811 20147 289839 20175
rect 289625 20085 289653 20113
rect 289687 20085 289715 20113
rect 289749 20085 289777 20113
rect 289811 20085 289839 20113
rect 289625 20023 289653 20051
rect 289687 20023 289715 20051
rect 289749 20023 289777 20051
rect 289811 20023 289839 20051
rect 289625 19961 289653 19989
rect 289687 19961 289715 19989
rect 289749 19961 289777 19989
rect 289811 19961 289839 19989
rect 289625 11147 289653 11175
rect 289687 11147 289715 11175
rect 289749 11147 289777 11175
rect 289811 11147 289839 11175
rect 289625 11085 289653 11113
rect 289687 11085 289715 11113
rect 289749 11085 289777 11113
rect 289811 11085 289839 11113
rect 289625 11023 289653 11051
rect 289687 11023 289715 11051
rect 289749 11023 289777 11051
rect 289811 11023 289839 11051
rect 289625 10961 289653 10989
rect 289687 10961 289715 10989
rect 289749 10961 289777 10989
rect 289811 10961 289839 10989
rect 289625 2147 289653 2175
rect 289687 2147 289715 2175
rect 289749 2147 289777 2175
rect 289811 2147 289839 2175
rect 289625 2085 289653 2113
rect 289687 2085 289715 2113
rect 289749 2085 289777 2113
rect 289811 2085 289839 2113
rect 289625 2023 289653 2051
rect 289687 2023 289715 2051
rect 289749 2023 289777 2051
rect 289811 2023 289839 2051
rect 289625 1961 289653 1989
rect 289687 1961 289715 1989
rect 289749 1961 289777 1989
rect 289811 1961 289839 1989
rect 289625 -108 289653 -80
rect 289687 -108 289715 -80
rect 289749 -108 289777 -80
rect 289811 -108 289839 -80
rect 289625 -170 289653 -142
rect 289687 -170 289715 -142
rect 289749 -170 289777 -142
rect 289811 -170 289839 -142
rect 289625 -232 289653 -204
rect 289687 -232 289715 -204
rect 289749 -232 289777 -204
rect 289811 -232 289839 -204
rect 289625 -294 289653 -266
rect 289687 -294 289715 -266
rect 289749 -294 289777 -266
rect 289811 -294 289839 -266
rect 291485 299058 291513 299086
rect 291547 299058 291575 299086
rect 291609 299058 291637 299086
rect 291671 299058 291699 299086
rect 291485 298996 291513 299024
rect 291547 298996 291575 299024
rect 291609 298996 291637 299024
rect 291671 298996 291699 299024
rect 291485 298934 291513 298962
rect 291547 298934 291575 298962
rect 291609 298934 291637 298962
rect 291671 298934 291699 298962
rect 291485 298872 291513 298900
rect 291547 298872 291575 298900
rect 291609 298872 291637 298900
rect 291671 298872 291699 298900
rect 298728 299058 298756 299086
rect 298790 299058 298818 299086
rect 298852 299058 298880 299086
rect 298914 299058 298942 299086
rect 298728 298996 298756 299024
rect 298790 298996 298818 299024
rect 298852 298996 298880 299024
rect 298914 298996 298942 299024
rect 298728 298934 298756 298962
rect 298790 298934 298818 298962
rect 298852 298934 298880 298962
rect 298914 298934 298942 298962
rect 298728 298872 298756 298900
rect 298790 298872 298818 298900
rect 298852 298872 298880 298900
rect 298914 298872 298942 298900
rect 291485 293147 291513 293175
rect 291547 293147 291575 293175
rect 291609 293147 291637 293175
rect 291671 293147 291699 293175
rect 291485 293085 291513 293113
rect 291547 293085 291575 293113
rect 291609 293085 291637 293113
rect 291671 293085 291699 293113
rect 291485 293023 291513 293051
rect 291547 293023 291575 293051
rect 291609 293023 291637 293051
rect 291671 293023 291699 293051
rect 291485 292961 291513 292989
rect 291547 292961 291575 292989
rect 291609 292961 291637 292989
rect 291671 292961 291699 292989
rect 291485 284147 291513 284175
rect 291547 284147 291575 284175
rect 291609 284147 291637 284175
rect 291671 284147 291699 284175
rect 291485 284085 291513 284113
rect 291547 284085 291575 284113
rect 291609 284085 291637 284113
rect 291671 284085 291699 284113
rect 291485 284023 291513 284051
rect 291547 284023 291575 284051
rect 291609 284023 291637 284051
rect 291671 284023 291699 284051
rect 291485 283961 291513 283989
rect 291547 283961 291575 283989
rect 291609 283961 291637 283989
rect 291671 283961 291699 283989
rect 291485 275147 291513 275175
rect 291547 275147 291575 275175
rect 291609 275147 291637 275175
rect 291671 275147 291699 275175
rect 291485 275085 291513 275113
rect 291547 275085 291575 275113
rect 291609 275085 291637 275113
rect 291671 275085 291699 275113
rect 291485 275023 291513 275051
rect 291547 275023 291575 275051
rect 291609 275023 291637 275051
rect 291671 275023 291699 275051
rect 291485 274961 291513 274989
rect 291547 274961 291575 274989
rect 291609 274961 291637 274989
rect 291671 274961 291699 274989
rect 291485 266147 291513 266175
rect 291547 266147 291575 266175
rect 291609 266147 291637 266175
rect 291671 266147 291699 266175
rect 291485 266085 291513 266113
rect 291547 266085 291575 266113
rect 291609 266085 291637 266113
rect 291671 266085 291699 266113
rect 291485 266023 291513 266051
rect 291547 266023 291575 266051
rect 291609 266023 291637 266051
rect 291671 266023 291699 266051
rect 291485 265961 291513 265989
rect 291547 265961 291575 265989
rect 291609 265961 291637 265989
rect 291671 265961 291699 265989
rect 291485 257147 291513 257175
rect 291547 257147 291575 257175
rect 291609 257147 291637 257175
rect 291671 257147 291699 257175
rect 291485 257085 291513 257113
rect 291547 257085 291575 257113
rect 291609 257085 291637 257113
rect 291671 257085 291699 257113
rect 291485 257023 291513 257051
rect 291547 257023 291575 257051
rect 291609 257023 291637 257051
rect 291671 257023 291699 257051
rect 291485 256961 291513 256989
rect 291547 256961 291575 256989
rect 291609 256961 291637 256989
rect 291671 256961 291699 256989
rect 291485 248147 291513 248175
rect 291547 248147 291575 248175
rect 291609 248147 291637 248175
rect 291671 248147 291699 248175
rect 291485 248085 291513 248113
rect 291547 248085 291575 248113
rect 291609 248085 291637 248113
rect 291671 248085 291699 248113
rect 291485 248023 291513 248051
rect 291547 248023 291575 248051
rect 291609 248023 291637 248051
rect 291671 248023 291699 248051
rect 291485 247961 291513 247989
rect 291547 247961 291575 247989
rect 291609 247961 291637 247989
rect 291671 247961 291699 247989
rect 291485 239147 291513 239175
rect 291547 239147 291575 239175
rect 291609 239147 291637 239175
rect 291671 239147 291699 239175
rect 291485 239085 291513 239113
rect 291547 239085 291575 239113
rect 291609 239085 291637 239113
rect 291671 239085 291699 239113
rect 291485 239023 291513 239051
rect 291547 239023 291575 239051
rect 291609 239023 291637 239051
rect 291671 239023 291699 239051
rect 291485 238961 291513 238989
rect 291547 238961 291575 238989
rect 291609 238961 291637 238989
rect 291671 238961 291699 238989
rect 291485 230147 291513 230175
rect 291547 230147 291575 230175
rect 291609 230147 291637 230175
rect 291671 230147 291699 230175
rect 291485 230085 291513 230113
rect 291547 230085 291575 230113
rect 291609 230085 291637 230113
rect 291671 230085 291699 230113
rect 291485 230023 291513 230051
rect 291547 230023 291575 230051
rect 291609 230023 291637 230051
rect 291671 230023 291699 230051
rect 291485 229961 291513 229989
rect 291547 229961 291575 229989
rect 291609 229961 291637 229989
rect 291671 229961 291699 229989
rect 291485 221147 291513 221175
rect 291547 221147 291575 221175
rect 291609 221147 291637 221175
rect 291671 221147 291699 221175
rect 291485 221085 291513 221113
rect 291547 221085 291575 221113
rect 291609 221085 291637 221113
rect 291671 221085 291699 221113
rect 291485 221023 291513 221051
rect 291547 221023 291575 221051
rect 291609 221023 291637 221051
rect 291671 221023 291699 221051
rect 291485 220961 291513 220989
rect 291547 220961 291575 220989
rect 291609 220961 291637 220989
rect 291671 220961 291699 220989
rect 291485 212147 291513 212175
rect 291547 212147 291575 212175
rect 291609 212147 291637 212175
rect 291671 212147 291699 212175
rect 291485 212085 291513 212113
rect 291547 212085 291575 212113
rect 291609 212085 291637 212113
rect 291671 212085 291699 212113
rect 291485 212023 291513 212051
rect 291547 212023 291575 212051
rect 291609 212023 291637 212051
rect 291671 212023 291699 212051
rect 291485 211961 291513 211989
rect 291547 211961 291575 211989
rect 291609 211961 291637 211989
rect 291671 211961 291699 211989
rect 291485 203147 291513 203175
rect 291547 203147 291575 203175
rect 291609 203147 291637 203175
rect 291671 203147 291699 203175
rect 291485 203085 291513 203113
rect 291547 203085 291575 203113
rect 291609 203085 291637 203113
rect 291671 203085 291699 203113
rect 291485 203023 291513 203051
rect 291547 203023 291575 203051
rect 291609 203023 291637 203051
rect 291671 203023 291699 203051
rect 291485 202961 291513 202989
rect 291547 202961 291575 202989
rect 291609 202961 291637 202989
rect 291671 202961 291699 202989
rect 291485 194147 291513 194175
rect 291547 194147 291575 194175
rect 291609 194147 291637 194175
rect 291671 194147 291699 194175
rect 291485 194085 291513 194113
rect 291547 194085 291575 194113
rect 291609 194085 291637 194113
rect 291671 194085 291699 194113
rect 291485 194023 291513 194051
rect 291547 194023 291575 194051
rect 291609 194023 291637 194051
rect 291671 194023 291699 194051
rect 291485 193961 291513 193989
rect 291547 193961 291575 193989
rect 291609 193961 291637 193989
rect 291671 193961 291699 193989
rect 291485 185147 291513 185175
rect 291547 185147 291575 185175
rect 291609 185147 291637 185175
rect 291671 185147 291699 185175
rect 291485 185085 291513 185113
rect 291547 185085 291575 185113
rect 291609 185085 291637 185113
rect 291671 185085 291699 185113
rect 291485 185023 291513 185051
rect 291547 185023 291575 185051
rect 291609 185023 291637 185051
rect 291671 185023 291699 185051
rect 291485 184961 291513 184989
rect 291547 184961 291575 184989
rect 291609 184961 291637 184989
rect 291671 184961 291699 184989
rect 291485 176147 291513 176175
rect 291547 176147 291575 176175
rect 291609 176147 291637 176175
rect 291671 176147 291699 176175
rect 291485 176085 291513 176113
rect 291547 176085 291575 176113
rect 291609 176085 291637 176113
rect 291671 176085 291699 176113
rect 291485 176023 291513 176051
rect 291547 176023 291575 176051
rect 291609 176023 291637 176051
rect 291671 176023 291699 176051
rect 291485 175961 291513 175989
rect 291547 175961 291575 175989
rect 291609 175961 291637 175989
rect 291671 175961 291699 175989
rect 291485 167147 291513 167175
rect 291547 167147 291575 167175
rect 291609 167147 291637 167175
rect 291671 167147 291699 167175
rect 291485 167085 291513 167113
rect 291547 167085 291575 167113
rect 291609 167085 291637 167113
rect 291671 167085 291699 167113
rect 291485 167023 291513 167051
rect 291547 167023 291575 167051
rect 291609 167023 291637 167051
rect 291671 167023 291699 167051
rect 291485 166961 291513 166989
rect 291547 166961 291575 166989
rect 291609 166961 291637 166989
rect 291671 166961 291699 166989
rect 291485 158147 291513 158175
rect 291547 158147 291575 158175
rect 291609 158147 291637 158175
rect 291671 158147 291699 158175
rect 291485 158085 291513 158113
rect 291547 158085 291575 158113
rect 291609 158085 291637 158113
rect 291671 158085 291699 158113
rect 291485 158023 291513 158051
rect 291547 158023 291575 158051
rect 291609 158023 291637 158051
rect 291671 158023 291699 158051
rect 291485 157961 291513 157989
rect 291547 157961 291575 157989
rect 291609 157961 291637 157989
rect 291671 157961 291699 157989
rect 291485 149147 291513 149175
rect 291547 149147 291575 149175
rect 291609 149147 291637 149175
rect 291671 149147 291699 149175
rect 291485 149085 291513 149113
rect 291547 149085 291575 149113
rect 291609 149085 291637 149113
rect 291671 149085 291699 149113
rect 291485 149023 291513 149051
rect 291547 149023 291575 149051
rect 291609 149023 291637 149051
rect 291671 149023 291699 149051
rect 291485 148961 291513 148989
rect 291547 148961 291575 148989
rect 291609 148961 291637 148989
rect 291671 148961 291699 148989
rect 291485 140147 291513 140175
rect 291547 140147 291575 140175
rect 291609 140147 291637 140175
rect 291671 140147 291699 140175
rect 291485 140085 291513 140113
rect 291547 140085 291575 140113
rect 291609 140085 291637 140113
rect 291671 140085 291699 140113
rect 291485 140023 291513 140051
rect 291547 140023 291575 140051
rect 291609 140023 291637 140051
rect 291671 140023 291699 140051
rect 291485 139961 291513 139989
rect 291547 139961 291575 139989
rect 291609 139961 291637 139989
rect 291671 139961 291699 139989
rect 291485 131147 291513 131175
rect 291547 131147 291575 131175
rect 291609 131147 291637 131175
rect 291671 131147 291699 131175
rect 291485 131085 291513 131113
rect 291547 131085 291575 131113
rect 291609 131085 291637 131113
rect 291671 131085 291699 131113
rect 291485 131023 291513 131051
rect 291547 131023 291575 131051
rect 291609 131023 291637 131051
rect 291671 131023 291699 131051
rect 291485 130961 291513 130989
rect 291547 130961 291575 130989
rect 291609 130961 291637 130989
rect 291671 130961 291699 130989
rect 291485 122147 291513 122175
rect 291547 122147 291575 122175
rect 291609 122147 291637 122175
rect 291671 122147 291699 122175
rect 291485 122085 291513 122113
rect 291547 122085 291575 122113
rect 291609 122085 291637 122113
rect 291671 122085 291699 122113
rect 291485 122023 291513 122051
rect 291547 122023 291575 122051
rect 291609 122023 291637 122051
rect 291671 122023 291699 122051
rect 291485 121961 291513 121989
rect 291547 121961 291575 121989
rect 291609 121961 291637 121989
rect 291671 121961 291699 121989
rect 291485 113147 291513 113175
rect 291547 113147 291575 113175
rect 291609 113147 291637 113175
rect 291671 113147 291699 113175
rect 291485 113085 291513 113113
rect 291547 113085 291575 113113
rect 291609 113085 291637 113113
rect 291671 113085 291699 113113
rect 291485 113023 291513 113051
rect 291547 113023 291575 113051
rect 291609 113023 291637 113051
rect 291671 113023 291699 113051
rect 291485 112961 291513 112989
rect 291547 112961 291575 112989
rect 291609 112961 291637 112989
rect 291671 112961 291699 112989
rect 291485 104147 291513 104175
rect 291547 104147 291575 104175
rect 291609 104147 291637 104175
rect 291671 104147 291699 104175
rect 291485 104085 291513 104113
rect 291547 104085 291575 104113
rect 291609 104085 291637 104113
rect 291671 104085 291699 104113
rect 291485 104023 291513 104051
rect 291547 104023 291575 104051
rect 291609 104023 291637 104051
rect 291671 104023 291699 104051
rect 291485 103961 291513 103989
rect 291547 103961 291575 103989
rect 291609 103961 291637 103989
rect 291671 103961 291699 103989
rect 291485 95147 291513 95175
rect 291547 95147 291575 95175
rect 291609 95147 291637 95175
rect 291671 95147 291699 95175
rect 291485 95085 291513 95113
rect 291547 95085 291575 95113
rect 291609 95085 291637 95113
rect 291671 95085 291699 95113
rect 291485 95023 291513 95051
rect 291547 95023 291575 95051
rect 291609 95023 291637 95051
rect 291671 95023 291699 95051
rect 291485 94961 291513 94989
rect 291547 94961 291575 94989
rect 291609 94961 291637 94989
rect 291671 94961 291699 94989
rect 291485 86147 291513 86175
rect 291547 86147 291575 86175
rect 291609 86147 291637 86175
rect 291671 86147 291699 86175
rect 291485 86085 291513 86113
rect 291547 86085 291575 86113
rect 291609 86085 291637 86113
rect 291671 86085 291699 86113
rect 291485 86023 291513 86051
rect 291547 86023 291575 86051
rect 291609 86023 291637 86051
rect 291671 86023 291699 86051
rect 291485 85961 291513 85989
rect 291547 85961 291575 85989
rect 291609 85961 291637 85989
rect 291671 85961 291699 85989
rect 291485 77147 291513 77175
rect 291547 77147 291575 77175
rect 291609 77147 291637 77175
rect 291671 77147 291699 77175
rect 291485 77085 291513 77113
rect 291547 77085 291575 77113
rect 291609 77085 291637 77113
rect 291671 77085 291699 77113
rect 291485 77023 291513 77051
rect 291547 77023 291575 77051
rect 291609 77023 291637 77051
rect 291671 77023 291699 77051
rect 291485 76961 291513 76989
rect 291547 76961 291575 76989
rect 291609 76961 291637 76989
rect 291671 76961 291699 76989
rect 291485 68147 291513 68175
rect 291547 68147 291575 68175
rect 291609 68147 291637 68175
rect 291671 68147 291699 68175
rect 291485 68085 291513 68113
rect 291547 68085 291575 68113
rect 291609 68085 291637 68113
rect 291671 68085 291699 68113
rect 291485 68023 291513 68051
rect 291547 68023 291575 68051
rect 291609 68023 291637 68051
rect 291671 68023 291699 68051
rect 291485 67961 291513 67989
rect 291547 67961 291575 67989
rect 291609 67961 291637 67989
rect 291671 67961 291699 67989
rect 291485 59147 291513 59175
rect 291547 59147 291575 59175
rect 291609 59147 291637 59175
rect 291671 59147 291699 59175
rect 291485 59085 291513 59113
rect 291547 59085 291575 59113
rect 291609 59085 291637 59113
rect 291671 59085 291699 59113
rect 291485 59023 291513 59051
rect 291547 59023 291575 59051
rect 291609 59023 291637 59051
rect 291671 59023 291699 59051
rect 291485 58961 291513 58989
rect 291547 58961 291575 58989
rect 291609 58961 291637 58989
rect 291671 58961 291699 58989
rect 291485 50147 291513 50175
rect 291547 50147 291575 50175
rect 291609 50147 291637 50175
rect 291671 50147 291699 50175
rect 291485 50085 291513 50113
rect 291547 50085 291575 50113
rect 291609 50085 291637 50113
rect 291671 50085 291699 50113
rect 291485 50023 291513 50051
rect 291547 50023 291575 50051
rect 291609 50023 291637 50051
rect 291671 50023 291699 50051
rect 291485 49961 291513 49989
rect 291547 49961 291575 49989
rect 291609 49961 291637 49989
rect 291671 49961 291699 49989
rect 291485 41147 291513 41175
rect 291547 41147 291575 41175
rect 291609 41147 291637 41175
rect 291671 41147 291699 41175
rect 291485 41085 291513 41113
rect 291547 41085 291575 41113
rect 291609 41085 291637 41113
rect 291671 41085 291699 41113
rect 291485 41023 291513 41051
rect 291547 41023 291575 41051
rect 291609 41023 291637 41051
rect 291671 41023 291699 41051
rect 291485 40961 291513 40989
rect 291547 40961 291575 40989
rect 291609 40961 291637 40989
rect 291671 40961 291699 40989
rect 291485 32147 291513 32175
rect 291547 32147 291575 32175
rect 291609 32147 291637 32175
rect 291671 32147 291699 32175
rect 291485 32085 291513 32113
rect 291547 32085 291575 32113
rect 291609 32085 291637 32113
rect 291671 32085 291699 32113
rect 291485 32023 291513 32051
rect 291547 32023 291575 32051
rect 291609 32023 291637 32051
rect 291671 32023 291699 32051
rect 291485 31961 291513 31989
rect 291547 31961 291575 31989
rect 291609 31961 291637 31989
rect 291671 31961 291699 31989
rect 291485 23147 291513 23175
rect 291547 23147 291575 23175
rect 291609 23147 291637 23175
rect 291671 23147 291699 23175
rect 291485 23085 291513 23113
rect 291547 23085 291575 23113
rect 291609 23085 291637 23113
rect 291671 23085 291699 23113
rect 291485 23023 291513 23051
rect 291547 23023 291575 23051
rect 291609 23023 291637 23051
rect 291671 23023 291699 23051
rect 291485 22961 291513 22989
rect 291547 22961 291575 22989
rect 291609 22961 291637 22989
rect 291671 22961 291699 22989
rect 291485 14147 291513 14175
rect 291547 14147 291575 14175
rect 291609 14147 291637 14175
rect 291671 14147 291699 14175
rect 291485 14085 291513 14113
rect 291547 14085 291575 14113
rect 291609 14085 291637 14113
rect 291671 14085 291699 14113
rect 291485 14023 291513 14051
rect 291547 14023 291575 14051
rect 291609 14023 291637 14051
rect 291671 14023 291699 14051
rect 291485 13961 291513 13989
rect 291547 13961 291575 13989
rect 291609 13961 291637 13989
rect 291671 13961 291699 13989
rect 291485 5147 291513 5175
rect 291547 5147 291575 5175
rect 291609 5147 291637 5175
rect 291671 5147 291699 5175
rect 291485 5085 291513 5113
rect 291547 5085 291575 5113
rect 291609 5085 291637 5113
rect 291671 5085 291699 5113
rect 291485 5023 291513 5051
rect 291547 5023 291575 5051
rect 291609 5023 291637 5051
rect 291671 5023 291699 5051
rect 291485 4961 291513 4989
rect 291547 4961 291575 4989
rect 291609 4961 291637 4989
rect 291671 4961 291699 4989
rect 298248 298578 298276 298606
rect 298310 298578 298338 298606
rect 298372 298578 298400 298606
rect 298434 298578 298462 298606
rect 298248 298516 298276 298544
rect 298310 298516 298338 298544
rect 298372 298516 298400 298544
rect 298434 298516 298462 298544
rect 298248 298454 298276 298482
rect 298310 298454 298338 298482
rect 298372 298454 298400 298482
rect 298434 298454 298462 298482
rect 298248 298392 298276 298420
rect 298310 298392 298338 298420
rect 298372 298392 298400 298420
rect 298434 298392 298462 298420
rect 298248 290147 298276 290175
rect 298310 290147 298338 290175
rect 298372 290147 298400 290175
rect 298434 290147 298462 290175
rect 298248 290085 298276 290113
rect 298310 290085 298338 290113
rect 298372 290085 298400 290113
rect 298434 290085 298462 290113
rect 298248 290023 298276 290051
rect 298310 290023 298338 290051
rect 298372 290023 298400 290051
rect 298434 290023 298462 290051
rect 298248 289961 298276 289989
rect 298310 289961 298338 289989
rect 298372 289961 298400 289989
rect 298434 289961 298462 289989
rect 298248 281147 298276 281175
rect 298310 281147 298338 281175
rect 298372 281147 298400 281175
rect 298434 281147 298462 281175
rect 298248 281085 298276 281113
rect 298310 281085 298338 281113
rect 298372 281085 298400 281113
rect 298434 281085 298462 281113
rect 298248 281023 298276 281051
rect 298310 281023 298338 281051
rect 298372 281023 298400 281051
rect 298434 281023 298462 281051
rect 298248 280961 298276 280989
rect 298310 280961 298338 280989
rect 298372 280961 298400 280989
rect 298434 280961 298462 280989
rect 298248 272147 298276 272175
rect 298310 272147 298338 272175
rect 298372 272147 298400 272175
rect 298434 272147 298462 272175
rect 298248 272085 298276 272113
rect 298310 272085 298338 272113
rect 298372 272085 298400 272113
rect 298434 272085 298462 272113
rect 298248 272023 298276 272051
rect 298310 272023 298338 272051
rect 298372 272023 298400 272051
rect 298434 272023 298462 272051
rect 298248 271961 298276 271989
rect 298310 271961 298338 271989
rect 298372 271961 298400 271989
rect 298434 271961 298462 271989
rect 298248 263147 298276 263175
rect 298310 263147 298338 263175
rect 298372 263147 298400 263175
rect 298434 263147 298462 263175
rect 298248 263085 298276 263113
rect 298310 263085 298338 263113
rect 298372 263085 298400 263113
rect 298434 263085 298462 263113
rect 298248 263023 298276 263051
rect 298310 263023 298338 263051
rect 298372 263023 298400 263051
rect 298434 263023 298462 263051
rect 298248 262961 298276 262989
rect 298310 262961 298338 262989
rect 298372 262961 298400 262989
rect 298434 262961 298462 262989
rect 298248 254147 298276 254175
rect 298310 254147 298338 254175
rect 298372 254147 298400 254175
rect 298434 254147 298462 254175
rect 298248 254085 298276 254113
rect 298310 254085 298338 254113
rect 298372 254085 298400 254113
rect 298434 254085 298462 254113
rect 298248 254023 298276 254051
rect 298310 254023 298338 254051
rect 298372 254023 298400 254051
rect 298434 254023 298462 254051
rect 298248 253961 298276 253989
rect 298310 253961 298338 253989
rect 298372 253961 298400 253989
rect 298434 253961 298462 253989
rect 298248 245147 298276 245175
rect 298310 245147 298338 245175
rect 298372 245147 298400 245175
rect 298434 245147 298462 245175
rect 298248 245085 298276 245113
rect 298310 245085 298338 245113
rect 298372 245085 298400 245113
rect 298434 245085 298462 245113
rect 298248 245023 298276 245051
rect 298310 245023 298338 245051
rect 298372 245023 298400 245051
rect 298434 245023 298462 245051
rect 298248 244961 298276 244989
rect 298310 244961 298338 244989
rect 298372 244961 298400 244989
rect 298434 244961 298462 244989
rect 298248 236147 298276 236175
rect 298310 236147 298338 236175
rect 298372 236147 298400 236175
rect 298434 236147 298462 236175
rect 298248 236085 298276 236113
rect 298310 236085 298338 236113
rect 298372 236085 298400 236113
rect 298434 236085 298462 236113
rect 298248 236023 298276 236051
rect 298310 236023 298338 236051
rect 298372 236023 298400 236051
rect 298434 236023 298462 236051
rect 298248 235961 298276 235989
rect 298310 235961 298338 235989
rect 298372 235961 298400 235989
rect 298434 235961 298462 235989
rect 298248 227147 298276 227175
rect 298310 227147 298338 227175
rect 298372 227147 298400 227175
rect 298434 227147 298462 227175
rect 298248 227085 298276 227113
rect 298310 227085 298338 227113
rect 298372 227085 298400 227113
rect 298434 227085 298462 227113
rect 298248 227023 298276 227051
rect 298310 227023 298338 227051
rect 298372 227023 298400 227051
rect 298434 227023 298462 227051
rect 298248 226961 298276 226989
rect 298310 226961 298338 226989
rect 298372 226961 298400 226989
rect 298434 226961 298462 226989
rect 298248 218147 298276 218175
rect 298310 218147 298338 218175
rect 298372 218147 298400 218175
rect 298434 218147 298462 218175
rect 298248 218085 298276 218113
rect 298310 218085 298338 218113
rect 298372 218085 298400 218113
rect 298434 218085 298462 218113
rect 298248 218023 298276 218051
rect 298310 218023 298338 218051
rect 298372 218023 298400 218051
rect 298434 218023 298462 218051
rect 298248 217961 298276 217989
rect 298310 217961 298338 217989
rect 298372 217961 298400 217989
rect 298434 217961 298462 217989
rect 298248 209147 298276 209175
rect 298310 209147 298338 209175
rect 298372 209147 298400 209175
rect 298434 209147 298462 209175
rect 298248 209085 298276 209113
rect 298310 209085 298338 209113
rect 298372 209085 298400 209113
rect 298434 209085 298462 209113
rect 298248 209023 298276 209051
rect 298310 209023 298338 209051
rect 298372 209023 298400 209051
rect 298434 209023 298462 209051
rect 298248 208961 298276 208989
rect 298310 208961 298338 208989
rect 298372 208961 298400 208989
rect 298434 208961 298462 208989
rect 298248 200147 298276 200175
rect 298310 200147 298338 200175
rect 298372 200147 298400 200175
rect 298434 200147 298462 200175
rect 298248 200085 298276 200113
rect 298310 200085 298338 200113
rect 298372 200085 298400 200113
rect 298434 200085 298462 200113
rect 298248 200023 298276 200051
rect 298310 200023 298338 200051
rect 298372 200023 298400 200051
rect 298434 200023 298462 200051
rect 298248 199961 298276 199989
rect 298310 199961 298338 199989
rect 298372 199961 298400 199989
rect 298434 199961 298462 199989
rect 298248 191147 298276 191175
rect 298310 191147 298338 191175
rect 298372 191147 298400 191175
rect 298434 191147 298462 191175
rect 298248 191085 298276 191113
rect 298310 191085 298338 191113
rect 298372 191085 298400 191113
rect 298434 191085 298462 191113
rect 298248 191023 298276 191051
rect 298310 191023 298338 191051
rect 298372 191023 298400 191051
rect 298434 191023 298462 191051
rect 298248 190961 298276 190989
rect 298310 190961 298338 190989
rect 298372 190961 298400 190989
rect 298434 190961 298462 190989
rect 298248 182147 298276 182175
rect 298310 182147 298338 182175
rect 298372 182147 298400 182175
rect 298434 182147 298462 182175
rect 298248 182085 298276 182113
rect 298310 182085 298338 182113
rect 298372 182085 298400 182113
rect 298434 182085 298462 182113
rect 298248 182023 298276 182051
rect 298310 182023 298338 182051
rect 298372 182023 298400 182051
rect 298434 182023 298462 182051
rect 298248 181961 298276 181989
rect 298310 181961 298338 181989
rect 298372 181961 298400 181989
rect 298434 181961 298462 181989
rect 298248 173147 298276 173175
rect 298310 173147 298338 173175
rect 298372 173147 298400 173175
rect 298434 173147 298462 173175
rect 298248 173085 298276 173113
rect 298310 173085 298338 173113
rect 298372 173085 298400 173113
rect 298434 173085 298462 173113
rect 298248 173023 298276 173051
rect 298310 173023 298338 173051
rect 298372 173023 298400 173051
rect 298434 173023 298462 173051
rect 298248 172961 298276 172989
rect 298310 172961 298338 172989
rect 298372 172961 298400 172989
rect 298434 172961 298462 172989
rect 298248 164147 298276 164175
rect 298310 164147 298338 164175
rect 298372 164147 298400 164175
rect 298434 164147 298462 164175
rect 298248 164085 298276 164113
rect 298310 164085 298338 164113
rect 298372 164085 298400 164113
rect 298434 164085 298462 164113
rect 298248 164023 298276 164051
rect 298310 164023 298338 164051
rect 298372 164023 298400 164051
rect 298434 164023 298462 164051
rect 298248 163961 298276 163989
rect 298310 163961 298338 163989
rect 298372 163961 298400 163989
rect 298434 163961 298462 163989
rect 298248 155147 298276 155175
rect 298310 155147 298338 155175
rect 298372 155147 298400 155175
rect 298434 155147 298462 155175
rect 298248 155085 298276 155113
rect 298310 155085 298338 155113
rect 298372 155085 298400 155113
rect 298434 155085 298462 155113
rect 298248 155023 298276 155051
rect 298310 155023 298338 155051
rect 298372 155023 298400 155051
rect 298434 155023 298462 155051
rect 298248 154961 298276 154989
rect 298310 154961 298338 154989
rect 298372 154961 298400 154989
rect 298434 154961 298462 154989
rect 298248 146147 298276 146175
rect 298310 146147 298338 146175
rect 298372 146147 298400 146175
rect 298434 146147 298462 146175
rect 298248 146085 298276 146113
rect 298310 146085 298338 146113
rect 298372 146085 298400 146113
rect 298434 146085 298462 146113
rect 298248 146023 298276 146051
rect 298310 146023 298338 146051
rect 298372 146023 298400 146051
rect 298434 146023 298462 146051
rect 298248 145961 298276 145989
rect 298310 145961 298338 145989
rect 298372 145961 298400 145989
rect 298434 145961 298462 145989
rect 298248 137147 298276 137175
rect 298310 137147 298338 137175
rect 298372 137147 298400 137175
rect 298434 137147 298462 137175
rect 298248 137085 298276 137113
rect 298310 137085 298338 137113
rect 298372 137085 298400 137113
rect 298434 137085 298462 137113
rect 298248 137023 298276 137051
rect 298310 137023 298338 137051
rect 298372 137023 298400 137051
rect 298434 137023 298462 137051
rect 298248 136961 298276 136989
rect 298310 136961 298338 136989
rect 298372 136961 298400 136989
rect 298434 136961 298462 136989
rect 298248 128147 298276 128175
rect 298310 128147 298338 128175
rect 298372 128147 298400 128175
rect 298434 128147 298462 128175
rect 298248 128085 298276 128113
rect 298310 128085 298338 128113
rect 298372 128085 298400 128113
rect 298434 128085 298462 128113
rect 298248 128023 298276 128051
rect 298310 128023 298338 128051
rect 298372 128023 298400 128051
rect 298434 128023 298462 128051
rect 298248 127961 298276 127989
rect 298310 127961 298338 127989
rect 298372 127961 298400 127989
rect 298434 127961 298462 127989
rect 298248 119147 298276 119175
rect 298310 119147 298338 119175
rect 298372 119147 298400 119175
rect 298434 119147 298462 119175
rect 298248 119085 298276 119113
rect 298310 119085 298338 119113
rect 298372 119085 298400 119113
rect 298434 119085 298462 119113
rect 298248 119023 298276 119051
rect 298310 119023 298338 119051
rect 298372 119023 298400 119051
rect 298434 119023 298462 119051
rect 298248 118961 298276 118989
rect 298310 118961 298338 118989
rect 298372 118961 298400 118989
rect 298434 118961 298462 118989
rect 298248 110147 298276 110175
rect 298310 110147 298338 110175
rect 298372 110147 298400 110175
rect 298434 110147 298462 110175
rect 298248 110085 298276 110113
rect 298310 110085 298338 110113
rect 298372 110085 298400 110113
rect 298434 110085 298462 110113
rect 298248 110023 298276 110051
rect 298310 110023 298338 110051
rect 298372 110023 298400 110051
rect 298434 110023 298462 110051
rect 298248 109961 298276 109989
rect 298310 109961 298338 109989
rect 298372 109961 298400 109989
rect 298434 109961 298462 109989
rect 298248 101147 298276 101175
rect 298310 101147 298338 101175
rect 298372 101147 298400 101175
rect 298434 101147 298462 101175
rect 298248 101085 298276 101113
rect 298310 101085 298338 101113
rect 298372 101085 298400 101113
rect 298434 101085 298462 101113
rect 298248 101023 298276 101051
rect 298310 101023 298338 101051
rect 298372 101023 298400 101051
rect 298434 101023 298462 101051
rect 298248 100961 298276 100989
rect 298310 100961 298338 100989
rect 298372 100961 298400 100989
rect 298434 100961 298462 100989
rect 298248 92147 298276 92175
rect 298310 92147 298338 92175
rect 298372 92147 298400 92175
rect 298434 92147 298462 92175
rect 298248 92085 298276 92113
rect 298310 92085 298338 92113
rect 298372 92085 298400 92113
rect 298434 92085 298462 92113
rect 298248 92023 298276 92051
rect 298310 92023 298338 92051
rect 298372 92023 298400 92051
rect 298434 92023 298462 92051
rect 298248 91961 298276 91989
rect 298310 91961 298338 91989
rect 298372 91961 298400 91989
rect 298434 91961 298462 91989
rect 298248 83147 298276 83175
rect 298310 83147 298338 83175
rect 298372 83147 298400 83175
rect 298434 83147 298462 83175
rect 298248 83085 298276 83113
rect 298310 83085 298338 83113
rect 298372 83085 298400 83113
rect 298434 83085 298462 83113
rect 298248 83023 298276 83051
rect 298310 83023 298338 83051
rect 298372 83023 298400 83051
rect 298434 83023 298462 83051
rect 298248 82961 298276 82989
rect 298310 82961 298338 82989
rect 298372 82961 298400 82989
rect 298434 82961 298462 82989
rect 298248 74147 298276 74175
rect 298310 74147 298338 74175
rect 298372 74147 298400 74175
rect 298434 74147 298462 74175
rect 298248 74085 298276 74113
rect 298310 74085 298338 74113
rect 298372 74085 298400 74113
rect 298434 74085 298462 74113
rect 298248 74023 298276 74051
rect 298310 74023 298338 74051
rect 298372 74023 298400 74051
rect 298434 74023 298462 74051
rect 298248 73961 298276 73989
rect 298310 73961 298338 73989
rect 298372 73961 298400 73989
rect 298434 73961 298462 73989
rect 298248 65147 298276 65175
rect 298310 65147 298338 65175
rect 298372 65147 298400 65175
rect 298434 65147 298462 65175
rect 298248 65085 298276 65113
rect 298310 65085 298338 65113
rect 298372 65085 298400 65113
rect 298434 65085 298462 65113
rect 298248 65023 298276 65051
rect 298310 65023 298338 65051
rect 298372 65023 298400 65051
rect 298434 65023 298462 65051
rect 298248 64961 298276 64989
rect 298310 64961 298338 64989
rect 298372 64961 298400 64989
rect 298434 64961 298462 64989
rect 298248 56147 298276 56175
rect 298310 56147 298338 56175
rect 298372 56147 298400 56175
rect 298434 56147 298462 56175
rect 298248 56085 298276 56113
rect 298310 56085 298338 56113
rect 298372 56085 298400 56113
rect 298434 56085 298462 56113
rect 298248 56023 298276 56051
rect 298310 56023 298338 56051
rect 298372 56023 298400 56051
rect 298434 56023 298462 56051
rect 298248 55961 298276 55989
rect 298310 55961 298338 55989
rect 298372 55961 298400 55989
rect 298434 55961 298462 55989
rect 298248 47147 298276 47175
rect 298310 47147 298338 47175
rect 298372 47147 298400 47175
rect 298434 47147 298462 47175
rect 298248 47085 298276 47113
rect 298310 47085 298338 47113
rect 298372 47085 298400 47113
rect 298434 47085 298462 47113
rect 298248 47023 298276 47051
rect 298310 47023 298338 47051
rect 298372 47023 298400 47051
rect 298434 47023 298462 47051
rect 298248 46961 298276 46989
rect 298310 46961 298338 46989
rect 298372 46961 298400 46989
rect 298434 46961 298462 46989
rect 298248 38147 298276 38175
rect 298310 38147 298338 38175
rect 298372 38147 298400 38175
rect 298434 38147 298462 38175
rect 298248 38085 298276 38113
rect 298310 38085 298338 38113
rect 298372 38085 298400 38113
rect 298434 38085 298462 38113
rect 298248 38023 298276 38051
rect 298310 38023 298338 38051
rect 298372 38023 298400 38051
rect 298434 38023 298462 38051
rect 298248 37961 298276 37989
rect 298310 37961 298338 37989
rect 298372 37961 298400 37989
rect 298434 37961 298462 37989
rect 298248 29147 298276 29175
rect 298310 29147 298338 29175
rect 298372 29147 298400 29175
rect 298434 29147 298462 29175
rect 298248 29085 298276 29113
rect 298310 29085 298338 29113
rect 298372 29085 298400 29113
rect 298434 29085 298462 29113
rect 298248 29023 298276 29051
rect 298310 29023 298338 29051
rect 298372 29023 298400 29051
rect 298434 29023 298462 29051
rect 298248 28961 298276 28989
rect 298310 28961 298338 28989
rect 298372 28961 298400 28989
rect 298434 28961 298462 28989
rect 298248 20147 298276 20175
rect 298310 20147 298338 20175
rect 298372 20147 298400 20175
rect 298434 20147 298462 20175
rect 298248 20085 298276 20113
rect 298310 20085 298338 20113
rect 298372 20085 298400 20113
rect 298434 20085 298462 20113
rect 298248 20023 298276 20051
rect 298310 20023 298338 20051
rect 298372 20023 298400 20051
rect 298434 20023 298462 20051
rect 298248 19961 298276 19989
rect 298310 19961 298338 19989
rect 298372 19961 298400 19989
rect 298434 19961 298462 19989
rect 298248 11147 298276 11175
rect 298310 11147 298338 11175
rect 298372 11147 298400 11175
rect 298434 11147 298462 11175
rect 298248 11085 298276 11113
rect 298310 11085 298338 11113
rect 298372 11085 298400 11113
rect 298434 11085 298462 11113
rect 298248 11023 298276 11051
rect 298310 11023 298338 11051
rect 298372 11023 298400 11051
rect 298434 11023 298462 11051
rect 298248 10961 298276 10989
rect 298310 10961 298338 10989
rect 298372 10961 298400 10989
rect 298434 10961 298462 10989
rect 298248 2147 298276 2175
rect 298310 2147 298338 2175
rect 298372 2147 298400 2175
rect 298434 2147 298462 2175
rect 298248 2085 298276 2113
rect 298310 2085 298338 2113
rect 298372 2085 298400 2113
rect 298434 2085 298462 2113
rect 298248 2023 298276 2051
rect 298310 2023 298338 2051
rect 298372 2023 298400 2051
rect 298434 2023 298462 2051
rect 298248 1961 298276 1989
rect 298310 1961 298338 1989
rect 298372 1961 298400 1989
rect 298434 1961 298462 1989
rect 298248 -108 298276 -80
rect 298310 -108 298338 -80
rect 298372 -108 298400 -80
rect 298434 -108 298462 -80
rect 298248 -170 298276 -142
rect 298310 -170 298338 -142
rect 298372 -170 298400 -142
rect 298434 -170 298462 -142
rect 298248 -232 298276 -204
rect 298310 -232 298338 -204
rect 298372 -232 298400 -204
rect 298434 -232 298462 -204
rect 298248 -294 298276 -266
rect 298310 -294 298338 -266
rect 298372 -294 298400 -266
rect 298434 -294 298462 -266
rect 298728 293147 298756 293175
rect 298790 293147 298818 293175
rect 298852 293147 298880 293175
rect 298914 293147 298942 293175
rect 298728 293085 298756 293113
rect 298790 293085 298818 293113
rect 298852 293085 298880 293113
rect 298914 293085 298942 293113
rect 298728 293023 298756 293051
rect 298790 293023 298818 293051
rect 298852 293023 298880 293051
rect 298914 293023 298942 293051
rect 298728 292961 298756 292989
rect 298790 292961 298818 292989
rect 298852 292961 298880 292989
rect 298914 292961 298942 292989
rect 298728 284147 298756 284175
rect 298790 284147 298818 284175
rect 298852 284147 298880 284175
rect 298914 284147 298942 284175
rect 298728 284085 298756 284113
rect 298790 284085 298818 284113
rect 298852 284085 298880 284113
rect 298914 284085 298942 284113
rect 298728 284023 298756 284051
rect 298790 284023 298818 284051
rect 298852 284023 298880 284051
rect 298914 284023 298942 284051
rect 298728 283961 298756 283989
rect 298790 283961 298818 283989
rect 298852 283961 298880 283989
rect 298914 283961 298942 283989
rect 298728 275147 298756 275175
rect 298790 275147 298818 275175
rect 298852 275147 298880 275175
rect 298914 275147 298942 275175
rect 298728 275085 298756 275113
rect 298790 275085 298818 275113
rect 298852 275085 298880 275113
rect 298914 275085 298942 275113
rect 298728 275023 298756 275051
rect 298790 275023 298818 275051
rect 298852 275023 298880 275051
rect 298914 275023 298942 275051
rect 298728 274961 298756 274989
rect 298790 274961 298818 274989
rect 298852 274961 298880 274989
rect 298914 274961 298942 274989
rect 298728 266147 298756 266175
rect 298790 266147 298818 266175
rect 298852 266147 298880 266175
rect 298914 266147 298942 266175
rect 298728 266085 298756 266113
rect 298790 266085 298818 266113
rect 298852 266085 298880 266113
rect 298914 266085 298942 266113
rect 298728 266023 298756 266051
rect 298790 266023 298818 266051
rect 298852 266023 298880 266051
rect 298914 266023 298942 266051
rect 298728 265961 298756 265989
rect 298790 265961 298818 265989
rect 298852 265961 298880 265989
rect 298914 265961 298942 265989
rect 298728 257147 298756 257175
rect 298790 257147 298818 257175
rect 298852 257147 298880 257175
rect 298914 257147 298942 257175
rect 298728 257085 298756 257113
rect 298790 257085 298818 257113
rect 298852 257085 298880 257113
rect 298914 257085 298942 257113
rect 298728 257023 298756 257051
rect 298790 257023 298818 257051
rect 298852 257023 298880 257051
rect 298914 257023 298942 257051
rect 298728 256961 298756 256989
rect 298790 256961 298818 256989
rect 298852 256961 298880 256989
rect 298914 256961 298942 256989
rect 298728 248147 298756 248175
rect 298790 248147 298818 248175
rect 298852 248147 298880 248175
rect 298914 248147 298942 248175
rect 298728 248085 298756 248113
rect 298790 248085 298818 248113
rect 298852 248085 298880 248113
rect 298914 248085 298942 248113
rect 298728 248023 298756 248051
rect 298790 248023 298818 248051
rect 298852 248023 298880 248051
rect 298914 248023 298942 248051
rect 298728 247961 298756 247989
rect 298790 247961 298818 247989
rect 298852 247961 298880 247989
rect 298914 247961 298942 247989
rect 298728 239147 298756 239175
rect 298790 239147 298818 239175
rect 298852 239147 298880 239175
rect 298914 239147 298942 239175
rect 298728 239085 298756 239113
rect 298790 239085 298818 239113
rect 298852 239085 298880 239113
rect 298914 239085 298942 239113
rect 298728 239023 298756 239051
rect 298790 239023 298818 239051
rect 298852 239023 298880 239051
rect 298914 239023 298942 239051
rect 298728 238961 298756 238989
rect 298790 238961 298818 238989
rect 298852 238961 298880 238989
rect 298914 238961 298942 238989
rect 298728 230147 298756 230175
rect 298790 230147 298818 230175
rect 298852 230147 298880 230175
rect 298914 230147 298942 230175
rect 298728 230085 298756 230113
rect 298790 230085 298818 230113
rect 298852 230085 298880 230113
rect 298914 230085 298942 230113
rect 298728 230023 298756 230051
rect 298790 230023 298818 230051
rect 298852 230023 298880 230051
rect 298914 230023 298942 230051
rect 298728 229961 298756 229989
rect 298790 229961 298818 229989
rect 298852 229961 298880 229989
rect 298914 229961 298942 229989
rect 298728 221147 298756 221175
rect 298790 221147 298818 221175
rect 298852 221147 298880 221175
rect 298914 221147 298942 221175
rect 298728 221085 298756 221113
rect 298790 221085 298818 221113
rect 298852 221085 298880 221113
rect 298914 221085 298942 221113
rect 298728 221023 298756 221051
rect 298790 221023 298818 221051
rect 298852 221023 298880 221051
rect 298914 221023 298942 221051
rect 298728 220961 298756 220989
rect 298790 220961 298818 220989
rect 298852 220961 298880 220989
rect 298914 220961 298942 220989
rect 298728 212147 298756 212175
rect 298790 212147 298818 212175
rect 298852 212147 298880 212175
rect 298914 212147 298942 212175
rect 298728 212085 298756 212113
rect 298790 212085 298818 212113
rect 298852 212085 298880 212113
rect 298914 212085 298942 212113
rect 298728 212023 298756 212051
rect 298790 212023 298818 212051
rect 298852 212023 298880 212051
rect 298914 212023 298942 212051
rect 298728 211961 298756 211989
rect 298790 211961 298818 211989
rect 298852 211961 298880 211989
rect 298914 211961 298942 211989
rect 298728 203147 298756 203175
rect 298790 203147 298818 203175
rect 298852 203147 298880 203175
rect 298914 203147 298942 203175
rect 298728 203085 298756 203113
rect 298790 203085 298818 203113
rect 298852 203085 298880 203113
rect 298914 203085 298942 203113
rect 298728 203023 298756 203051
rect 298790 203023 298818 203051
rect 298852 203023 298880 203051
rect 298914 203023 298942 203051
rect 298728 202961 298756 202989
rect 298790 202961 298818 202989
rect 298852 202961 298880 202989
rect 298914 202961 298942 202989
rect 298728 194147 298756 194175
rect 298790 194147 298818 194175
rect 298852 194147 298880 194175
rect 298914 194147 298942 194175
rect 298728 194085 298756 194113
rect 298790 194085 298818 194113
rect 298852 194085 298880 194113
rect 298914 194085 298942 194113
rect 298728 194023 298756 194051
rect 298790 194023 298818 194051
rect 298852 194023 298880 194051
rect 298914 194023 298942 194051
rect 298728 193961 298756 193989
rect 298790 193961 298818 193989
rect 298852 193961 298880 193989
rect 298914 193961 298942 193989
rect 298728 185147 298756 185175
rect 298790 185147 298818 185175
rect 298852 185147 298880 185175
rect 298914 185147 298942 185175
rect 298728 185085 298756 185113
rect 298790 185085 298818 185113
rect 298852 185085 298880 185113
rect 298914 185085 298942 185113
rect 298728 185023 298756 185051
rect 298790 185023 298818 185051
rect 298852 185023 298880 185051
rect 298914 185023 298942 185051
rect 298728 184961 298756 184989
rect 298790 184961 298818 184989
rect 298852 184961 298880 184989
rect 298914 184961 298942 184989
rect 298728 176147 298756 176175
rect 298790 176147 298818 176175
rect 298852 176147 298880 176175
rect 298914 176147 298942 176175
rect 298728 176085 298756 176113
rect 298790 176085 298818 176113
rect 298852 176085 298880 176113
rect 298914 176085 298942 176113
rect 298728 176023 298756 176051
rect 298790 176023 298818 176051
rect 298852 176023 298880 176051
rect 298914 176023 298942 176051
rect 298728 175961 298756 175989
rect 298790 175961 298818 175989
rect 298852 175961 298880 175989
rect 298914 175961 298942 175989
rect 298728 167147 298756 167175
rect 298790 167147 298818 167175
rect 298852 167147 298880 167175
rect 298914 167147 298942 167175
rect 298728 167085 298756 167113
rect 298790 167085 298818 167113
rect 298852 167085 298880 167113
rect 298914 167085 298942 167113
rect 298728 167023 298756 167051
rect 298790 167023 298818 167051
rect 298852 167023 298880 167051
rect 298914 167023 298942 167051
rect 298728 166961 298756 166989
rect 298790 166961 298818 166989
rect 298852 166961 298880 166989
rect 298914 166961 298942 166989
rect 298728 158147 298756 158175
rect 298790 158147 298818 158175
rect 298852 158147 298880 158175
rect 298914 158147 298942 158175
rect 298728 158085 298756 158113
rect 298790 158085 298818 158113
rect 298852 158085 298880 158113
rect 298914 158085 298942 158113
rect 298728 158023 298756 158051
rect 298790 158023 298818 158051
rect 298852 158023 298880 158051
rect 298914 158023 298942 158051
rect 298728 157961 298756 157989
rect 298790 157961 298818 157989
rect 298852 157961 298880 157989
rect 298914 157961 298942 157989
rect 298728 149147 298756 149175
rect 298790 149147 298818 149175
rect 298852 149147 298880 149175
rect 298914 149147 298942 149175
rect 298728 149085 298756 149113
rect 298790 149085 298818 149113
rect 298852 149085 298880 149113
rect 298914 149085 298942 149113
rect 298728 149023 298756 149051
rect 298790 149023 298818 149051
rect 298852 149023 298880 149051
rect 298914 149023 298942 149051
rect 298728 148961 298756 148989
rect 298790 148961 298818 148989
rect 298852 148961 298880 148989
rect 298914 148961 298942 148989
rect 298728 140147 298756 140175
rect 298790 140147 298818 140175
rect 298852 140147 298880 140175
rect 298914 140147 298942 140175
rect 298728 140085 298756 140113
rect 298790 140085 298818 140113
rect 298852 140085 298880 140113
rect 298914 140085 298942 140113
rect 298728 140023 298756 140051
rect 298790 140023 298818 140051
rect 298852 140023 298880 140051
rect 298914 140023 298942 140051
rect 298728 139961 298756 139989
rect 298790 139961 298818 139989
rect 298852 139961 298880 139989
rect 298914 139961 298942 139989
rect 298728 131147 298756 131175
rect 298790 131147 298818 131175
rect 298852 131147 298880 131175
rect 298914 131147 298942 131175
rect 298728 131085 298756 131113
rect 298790 131085 298818 131113
rect 298852 131085 298880 131113
rect 298914 131085 298942 131113
rect 298728 131023 298756 131051
rect 298790 131023 298818 131051
rect 298852 131023 298880 131051
rect 298914 131023 298942 131051
rect 298728 130961 298756 130989
rect 298790 130961 298818 130989
rect 298852 130961 298880 130989
rect 298914 130961 298942 130989
rect 298728 122147 298756 122175
rect 298790 122147 298818 122175
rect 298852 122147 298880 122175
rect 298914 122147 298942 122175
rect 298728 122085 298756 122113
rect 298790 122085 298818 122113
rect 298852 122085 298880 122113
rect 298914 122085 298942 122113
rect 298728 122023 298756 122051
rect 298790 122023 298818 122051
rect 298852 122023 298880 122051
rect 298914 122023 298942 122051
rect 298728 121961 298756 121989
rect 298790 121961 298818 121989
rect 298852 121961 298880 121989
rect 298914 121961 298942 121989
rect 298728 113147 298756 113175
rect 298790 113147 298818 113175
rect 298852 113147 298880 113175
rect 298914 113147 298942 113175
rect 298728 113085 298756 113113
rect 298790 113085 298818 113113
rect 298852 113085 298880 113113
rect 298914 113085 298942 113113
rect 298728 113023 298756 113051
rect 298790 113023 298818 113051
rect 298852 113023 298880 113051
rect 298914 113023 298942 113051
rect 298728 112961 298756 112989
rect 298790 112961 298818 112989
rect 298852 112961 298880 112989
rect 298914 112961 298942 112989
rect 298728 104147 298756 104175
rect 298790 104147 298818 104175
rect 298852 104147 298880 104175
rect 298914 104147 298942 104175
rect 298728 104085 298756 104113
rect 298790 104085 298818 104113
rect 298852 104085 298880 104113
rect 298914 104085 298942 104113
rect 298728 104023 298756 104051
rect 298790 104023 298818 104051
rect 298852 104023 298880 104051
rect 298914 104023 298942 104051
rect 298728 103961 298756 103989
rect 298790 103961 298818 103989
rect 298852 103961 298880 103989
rect 298914 103961 298942 103989
rect 298728 95147 298756 95175
rect 298790 95147 298818 95175
rect 298852 95147 298880 95175
rect 298914 95147 298942 95175
rect 298728 95085 298756 95113
rect 298790 95085 298818 95113
rect 298852 95085 298880 95113
rect 298914 95085 298942 95113
rect 298728 95023 298756 95051
rect 298790 95023 298818 95051
rect 298852 95023 298880 95051
rect 298914 95023 298942 95051
rect 298728 94961 298756 94989
rect 298790 94961 298818 94989
rect 298852 94961 298880 94989
rect 298914 94961 298942 94989
rect 298728 86147 298756 86175
rect 298790 86147 298818 86175
rect 298852 86147 298880 86175
rect 298914 86147 298942 86175
rect 298728 86085 298756 86113
rect 298790 86085 298818 86113
rect 298852 86085 298880 86113
rect 298914 86085 298942 86113
rect 298728 86023 298756 86051
rect 298790 86023 298818 86051
rect 298852 86023 298880 86051
rect 298914 86023 298942 86051
rect 298728 85961 298756 85989
rect 298790 85961 298818 85989
rect 298852 85961 298880 85989
rect 298914 85961 298942 85989
rect 298728 77147 298756 77175
rect 298790 77147 298818 77175
rect 298852 77147 298880 77175
rect 298914 77147 298942 77175
rect 298728 77085 298756 77113
rect 298790 77085 298818 77113
rect 298852 77085 298880 77113
rect 298914 77085 298942 77113
rect 298728 77023 298756 77051
rect 298790 77023 298818 77051
rect 298852 77023 298880 77051
rect 298914 77023 298942 77051
rect 298728 76961 298756 76989
rect 298790 76961 298818 76989
rect 298852 76961 298880 76989
rect 298914 76961 298942 76989
rect 298728 68147 298756 68175
rect 298790 68147 298818 68175
rect 298852 68147 298880 68175
rect 298914 68147 298942 68175
rect 298728 68085 298756 68113
rect 298790 68085 298818 68113
rect 298852 68085 298880 68113
rect 298914 68085 298942 68113
rect 298728 68023 298756 68051
rect 298790 68023 298818 68051
rect 298852 68023 298880 68051
rect 298914 68023 298942 68051
rect 298728 67961 298756 67989
rect 298790 67961 298818 67989
rect 298852 67961 298880 67989
rect 298914 67961 298942 67989
rect 298728 59147 298756 59175
rect 298790 59147 298818 59175
rect 298852 59147 298880 59175
rect 298914 59147 298942 59175
rect 298728 59085 298756 59113
rect 298790 59085 298818 59113
rect 298852 59085 298880 59113
rect 298914 59085 298942 59113
rect 298728 59023 298756 59051
rect 298790 59023 298818 59051
rect 298852 59023 298880 59051
rect 298914 59023 298942 59051
rect 298728 58961 298756 58989
rect 298790 58961 298818 58989
rect 298852 58961 298880 58989
rect 298914 58961 298942 58989
rect 298728 50147 298756 50175
rect 298790 50147 298818 50175
rect 298852 50147 298880 50175
rect 298914 50147 298942 50175
rect 298728 50085 298756 50113
rect 298790 50085 298818 50113
rect 298852 50085 298880 50113
rect 298914 50085 298942 50113
rect 298728 50023 298756 50051
rect 298790 50023 298818 50051
rect 298852 50023 298880 50051
rect 298914 50023 298942 50051
rect 298728 49961 298756 49989
rect 298790 49961 298818 49989
rect 298852 49961 298880 49989
rect 298914 49961 298942 49989
rect 298728 41147 298756 41175
rect 298790 41147 298818 41175
rect 298852 41147 298880 41175
rect 298914 41147 298942 41175
rect 298728 41085 298756 41113
rect 298790 41085 298818 41113
rect 298852 41085 298880 41113
rect 298914 41085 298942 41113
rect 298728 41023 298756 41051
rect 298790 41023 298818 41051
rect 298852 41023 298880 41051
rect 298914 41023 298942 41051
rect 298728 40961 298756 40989
rect 298790 40961 298818 40989
rect 298852 40961 298880 40989
rect 298914 40961 298942 40989
rect 298728 32147 298756 32175
rect 298790 32147 298818 32175
rect 298852 32147 298880 32175
rect 298914 32147 298942 32175
rect 298728 32085 298756 32113
rect 298790 32085 298818 32113
rect 298852 32085 298880 32113
rect 298914 32085 298942 32113
rect 298728 32023 298756 32051
rect 298790 32023 298818 32051
rect 298852 32023 298880 32051
rect 298914 32023 298942 32051
rect 298728 31961 298756 31989
rect 298790 31961 298818 31989
rect 298852 31961 298880 31989
rect 298914 31961 298942 31989
rect 298728 23147 298756 23175
rect 298790 23147 298818 23175
rect 298852 23147 298880 23175
rect 298914 23147 298942 23175
rect 298728 23085 298756 23113
rect 298790 23085 298818 23113
rect 298852 23085 298880 23113
rect 298914 23085 298942 23113
rect 298728 23023 298756 23051
rect 298790 23023 298818 23051
rect 298852 23023 298880 23051
rect 298914 23023 298942 23051
rect 298728 22961 298756 22989
rect 298790 22961 298818 22989
rect 298852 22961 298880 22989
rect 298914 22961 298942 22989
rect 298728 14147 298756 14175
rect 298790 14147 298818 14175
rect 298852 14147 298880 14175
rect 298914 14147 298942 14175
rect 298728 14085 298756 14113
rect 298790 14085 298818 14113
rect 298852 14085 298880 14113
rect 298914 14085 298942 14113
rect 298728 14023 298756 14051
rect 298790 14023 298818 14051
rect 298852 14023 298880 14051
rect 298914 14023 298942 14051
rect 298728 13961 298756 13989
rect 298790 13961 298818 13989
rect 298852 13961 298880 13989
rect 298914 13961 298942 13989
rect 298728 5147 298756 5175
rect 298790 5147 298818 5175
rect 298852 5147 298880 5175
rect 298914 5147 298942 5175
rect 298728 5085 298756 5113
rect 298790 5085 298818 5113
rect 298852 5085 298880 5113
rect 298914 5085 298942 5113
rect 298728 5023 298756 5051
rect 298790 5023 298818 5051
rect 298852 5023 298880 5051
rect 298914 5023 298942 5051
rect 298728 4961 298756 4989
rect 298790 4961 298818 4989
rect 298852 4961 298880 4989
rect 298914 4961 298942 4989
rect 291485 -588 291513 -560
rect 291547 -588 291575 -560
rect 291609 -588 291637 -560
rect 291671 -588 291699 -560
rect 291485 -650 291513 -622
rect 291547 -650 291575 -622
rect 291609 -650 291637 -622
rect 291671 -650 291699 -622
rect 291485 -712 291513 -684
rect 291547 -712 291575 -684
rect 291609 -712 291637 -684
rect 291671 -712 291699 -684
rect 291485 -774 291513 -746
rect 291547 -774 291575 -746
rect 291609 -774 291637 -746
rect 291671 -774 291699 -746
rect 298728 -588 298756 -560
rect 298790 -588 298818 -560
rect 298852 -588 298880 -560
rect 298914 -588 298942 -560
rect 298728 -650 298756 -622
rect 298790 -650 298818 -622
rect 298852 -650 298880 -622
rect 298914 -650 298942 -622
rect 298728 -712 298756 -684
rect 298790 -712 298818 -684
rect 298852 -712 298880 -684
rect 298914 -712 298942 -684
rect 298728 -774 298756 -746
rect 298790 -774 298818 -746
rect 298852 -774 298880 -746
rect 298914 -774 298942 -746
<< metal5 >>
rect -958 299086 298990 299134
rect -958 299058 -910 299086
rect -882 299058 -848 299086
rect -820 299058 -786 299086
rect -758 299058 -724 299086
rect -696 299058 3485 299086
rect 3513 299058 3547 299086
rect 3575 299058 3609 299086
rect 3637 299058 3671 299086
rect 3699 299058 12485 299086
rect 12513 299058 12547 299086
rect 12575 299058 12609 299086
rect 12637 299058 12671 299086
rect 12699 299058 21485 299086
rect 21513 299058 21547 299086
rect 21575 299058 21609 299086
rect 21637 299058 21671 299086
rect 21699 299058 30485 299086
rect 30513 299058 30547 299086
rect 30575 299058 30609 299086
rect 30637 299058 30671 299086
rect 30699 299058 39485 299086
rect 39513 299058 39547 299086
rect 39575 299058 39609 299086
rect 39637 299058 39671 299086
rect 39699 299058 48485 299086
rect 48513 299058 48547 299086
rect 48575 299058 48609 299086
rect 48637 299058 48671 299086
rect 48699 299058 57485 299086
rect 57513 299058 57547 299086
rect 57575 299058 57609 299086
rect 57637 299058 57671 299086
rect 57699 299058 66485 299086
rect 66513 299058 66547 299086
rect 66575 299058 66609 299086
rect 66637 299058 66671 299086
rect 66699 299058 75485 299086
rect 75513 299058 75547 299086
rect 75575 299058 75609 299086
rect 75637 299058 75671 299086
rect 75699 299058 84485 299086
rect 84513 299058 84547 299086
rect 84575 299058 84609 299086
rect 84637 299058 84671 299086
rect 84699 299058 93485 299086
rect 93513 299058 93547 299086
rect 93575 299058 93609 299086
rect 93637 299058 93671 299086
rect 93699 299058 102485 299086
rect 102513 299058 102547 299086
rect 102575 299058 102609 299086
rect 102637 299058 102671 299086
rect 102699 299058 111485 299086
rect 111513 299058 111547 299086
rect 111575 299058 111609 299086
rect 111637 299058 111671 299086
rect 111699 299058 120485 299086
rect 120513 299058 120547 299086
rect 120575 299058 120609 299086
rect 120637 299058 120671 299086
rect 120699 299058 129485 299086
rect 129513 299058 129547 299086
rect 129575 299058 129609 299086
rect 129637 299058 129671 299086
rect 129699 299058 138485 299086
rect 138513 299058 138547 299086
rect 138575 299058 138609 299086
rect 138637 299058 138671 299086
rect 138699 299058 147485 299086
rect 147513 299058 147547 299086
rect 147575 299058 147609 299086
rect 147637 299058 147671 299086
rect 147699 299058 156485 299086
rect 156513 299058 156547 299086
rect 156575 299058 156609 299086
rect 156637 299058 156671 299086
rect 156699 299058 165485 299086
rect 165513 299058 165547 299086
rect 165575 299058 165609 299086
rect 165637 299058 165671 299086
rect 165699 299058 174485 299086
rect 174513 299058 174547 299086
rect 174575 299058 174609 299086
rect 174637 299058 174671 299086
rect 174699 299058 183485 299086
rect 183513 299058 183547 299086
rect 183575 299058 183609 299086
rect 183637 299058 183671 299086
rect 183699 299058 192485 299086
rect 192513 299058 192547 299086
rect 192575 299058 192609 299086
rect 192637 299058 192671 299086
rect 192699 299058 201485 299086
rect 201513 299058 201547 299086
rect 201575 299058 201609 299086
rect 201637 299058 201671 299086
rect 201699 299058 210485 299086
rect 210513 299058 210547 299086
rect 210575 299058 210609 299086
rect 210637 299058 210671 299086
rect 210699 299058 219485 299086
rect 219513 299058 219547 299086
rect 219575 299058 219609 299086
rect 219637 299058 219671 299086
rect 219699 299058 228485 299086
rect 228513 299058 228547 299086
rect 228575 299058 228609 299086
rect 228637 299058 228671 299086
rect 228699 299058 237485 299086
rect 237513 299058 237547 299086
rect 237575 299058 237609 299086
rect 237637 299058 237671 299086
rect 237699 299058 246485 299086
rect 246513 299058 246547 299086
rect 246575 299058 246609 299086
rect 246637 299058 246671 299086
rect 246699 299058 255485 299086
rect 255513 299058 255547 299086
rect 255575 299058 255609 299086
rect 255637 299058 255671 299086
rect 255699 299058 264485 299086
rect 264513 299058 264547 299086
rect 264575 299058 264609 299086
rect 264637 299058 264671 299086
rect 264699 299058 273485 299086
rect 273513 299058 273547 299086
rect 273575 299058 273609 299086
rect 273637 299058 273671 299086
rect 273699 299058 282485 299086
rect 282513 299058 282547 299086
rect 282575 299058 282609 299086
rect 282637 299058 282671 299086
rect 282699 299058 291485 299086
rect 291513 299058 291547 299086
rect 291575 299058 291609 299086
rect 291637 299058 291671 299086
rect 291699 299058 298728 299086
rect 298756 299058 298790 299086
rect 298818 299058 298852 299086
rect 298880 299058 298914 299086
rect 298942 299058 298990 299086
rect -958 299024 298990 299058
rect -958 298996 -910 299024
rect -882 298996 -848 299024
rect -820 298996 -786 299024
rect -758 298996 -724 299024
rect -696 298996 3485 299024
rect 3513 298996 3547 299024
rect 3575 298996 3609 299024
rect 3637 298996 3671 299024
rect 3699 298996 12485 299024
rect 12513 298996 12547 299024
rect 12575 298996 12609 299024
rect 12637 298996 12671 299024
rect 12699 298996 21485 299024
rect 21513 298996 21547 299024
rect 21575 298996 21609 299024
rect 21637 298996 21671 299024
rect 21699 298996 30485 299024
rect 30513 298996 30547 299024
rect 30575 298996 30609 299024
rect 30637 298996 30671 299024
rect 30699 298996 39485 299024
rect 39513 298996 39547 299024
rect 39575 298996 39609 299024
rect 39637 298996 39671 299024
rect 39699 298996 48485 299024
rect 48513 298996 48547 299024
rect 48575 298996 48609 299024
rect 48637 298996 48671 299024
rect 48699 298996 57485 299024
rect 57513 298996 57547 299024
rect 57575 298996 57609 299024
rect 57637 298996 57671 299024
rect 57699 298996 66485 299024
rect 66513 298996 66547 299024
rect 66575 298996 66609 299024
rect 66637 298996 66671 299024
rect 66699 298996 75485 299024
rect 75513 298996 75547 299024
rect 75575 298996 75609 299024
rect 75637 298996 75671 299024
rect 75699 298996 84485 299024
rect 84513 298996 84547 299024
rect 84575 298996 84609 299024
rect 84637 298996 84671 299024
rect 84699 298996 93485 299024
rect 93513 298996 93547 299024
rect 93575 298996 93609 299024
rect 93637 298996 93671 299024
rect 93699 298996 102485 299024
rect 102513 298996 102547 299024
rect 102575 298996 102609 299024
rect 102637 298996 102671 299024
rect 102699 298996 111485 299024
rect 111513 298996 111547 299024
rect 111575 298996 111609 299024
rect 111637 298996 111671 299024
rect 111699 298996 120485 299024
rect 120513 298996 120547 299024
rect 120575 298996 120609 299024
rect 120637 298996 120671 299024
rect 120699 298996 129485 299024
rect 129513 298996 129547 299024
rect 129575 298996 129609 299024
rect 129637 298996 129671 299024
rect 129699 298996 138485 299024
rect 138513 298996 138547 299024
rect 138575 298996 138609 299024
rect 138637 298996 138671 299024
rect 138699 298996 147485 299024
rect 147513 298996 147547 299024
rect 147575 298996 147609 299024
rect 147637 298996 147671 299024
rect 147699 298996 156485 299024
rect 156513 298996 156547 299024
rect 156575 298996 156609 299024
rect 156637 298996 156671 299024
rect 156699 298996 165485 299024
rect 165513 298996 165547 299024
rect 165575 298996 165609 299024
rect 165637 298996 165671 299024
rect 165699 298996 174485 299024
rect 174513 298996 174547 299024
rect 174575 298996 174609 299024
rect 174637 298996 174671 299024
rect 174699 298996 183485 299024
rect 183513 298996 183547 299024
rect 183575 298996 183609 299024
rect 183637 298996 183671 299024
rect 183699 298996 192485 299024
rect 192513 298996 192547 299024
rect 192575 298996 192609 299024
rect 192637 298996 192671 299024
rect 192699 298996 201485 299024
rect 201513 298996 201547 299024
rect 201575 298996 201609 299024
rect 201637 298996 201671 299024
rect 201699 298996 210485 299024
rect 210513 298996 210547 299024
rect 210575 298996 210609 299024
rect 210637 298996 210671 299024
rect 210699 298996 219485 299024
rect 219513 298996 219547 299024
rect 219575 298996 219609 299024
rect 219637 298996 219671 299024
rect 219699 298996 228485 299024
rect 228513 298996 228547 299024
rect 228575 298996 228609 299024
rect 228637 298996 228671 299024
rect 228699 298996 237485 299024
rect 237513 298996 237547 299024
rect 237575 298996 237609 299024
rect 237637 298996 237671 299024
rect 237699 298996 246485 299024
rect 246513 298996 246547 299024
rect 246575 298996 246609 299024
rect 246637 298996 246671 299024
rect 246699 298996 255485 299024
rect 255513 298996 255547 299024
rect 255575 298996 255609 299024
rect 255637 298996 255671 299024
rect 255699 298996 264485 299024
rect 264513 298996 264547 299024
rect 264575 298996 264609 299024
rect 264637 298996 264671 299024
rect 264699 298996 273485 299024
rect 273513 298996 273547 299024
rect 273575 298996 273609 299024
rect 273637 298996 273671 299024
rect 273699 298996 282485 299024
rect 282513 298996 282547 299024
rect 282575 298996 282609 299024
rect 282637 298996 282671 299024
rect 282699 298996 291485 299024
rect 291513 298996 291547 299024
rect 291575 298996 291609 299024
rect 291637 298996 291671 299024
rect 291699 298996 298728 299024
rect 298756 298996 298790 299024
rect 298818 298996 298852 299024
rect 298880 298996 298914 299024
rect 298942 298996 298990 299024
rect -958 298962 298990 298996
rect -958 298934 -910 298962
rect -882 298934 -848 298962
rect -820 298934 -786 298962
rect -758 298934 -724 298962
rect -696 298934 3485 298962
rect 3513 298934 3547 298962
rect 3575 298934 3609 298962
rect 3637 298934 3671 298962
rect 3699 298934 12485 298962
rect 12513 298934 12547 298962
rect 12575 298934 12609 298962
rect 12637 298934 12671 298962
rect 12699 298934 21485 298962
rect 21513 298934 21547 298962
rect 21575 298934 21609 298962
rect 21637 298934 21671 298962
rect 21699 298934 30485 298962
rect 30513 298934 30547 298962
rect 30575 298934 30609 298962
rect 30637 298934 30671 298962
rect 30699 298934 39485 298962
rect 39513 298934 39547 298962
rect 39575 298934 39609 298962
rect 39637 298934 39671 298962
rect 39699 298934 48485 298962
rect 48513 298934 48547 298962
rect 48575 298934 48609 298962
rect 48637 298934 48671 298962
rect 48699 298934 57485 298962
rect 57513 298934 57547 298962
rect 57575 298934 57609 298962
rect 57637 298934 57671 298962
rect 57699 298934 66485 298962
rect 66513 298934 66547 298962
rect 66575 298934 66609 298962
rect 66637 298934 66671 298962
rect 66699 298934 75485 298962
rect 75513 298934 75547 298962
rect 75575 298934 75609 298962
rect 75637 298934 75671 298962
rect 75699 298934 84485 298962
rect 84513 298934 84547 298962
rect 84575 298934 84609 298962
rect 84637 298934 84671 298962
rect 84699 298934 93485 298962
rect 93513 298934 93547 298962
rect 93575 298934 93609 298962
rect 93637 298934 93671 298962
rect 93699 298934 102485 298962
rect 102513 298934 102547 298962
rect 102575 298934 102609 298962
rect 102637 298934 102671 298962
rect 102699 298934 111485 298962
rect 111513 298934 111547 298962
rect 111575 298934 111609 298962
rect 111637 298934 111671 298962
rect 111699 298934 120485 298962
rect 120513 298934 120547 298962
rect 120575 298934 120609 298962
rect 120637 298934 120671 298962
rect 120699 298934 129485 298962
rect 129513 298934 129547 298962
rect 129575 298934 129609 298962
rect 129637 298934 129671 298962
rect 129699 298934 138485 298962
rect 138513 298934 138547 298962
rect 138575 298934 138609 298962
rect 138637 298934 138671 298962
rect 138699 298934 147485 298962
rect 147513 298934 147547 298962
rect 147575 298934 147609 298962
rect 147637 298934 147671 298962
rect 147699 298934 156485 298962
rect 156513 298934 156547 298962
rect 156575 298934 156609 298962
rect 156637 298934 156671 298962
rect 156699 298934 165485 298962
rect 165513 298934 165547 298962
rect 165575 298934 165609 298962
rect 165637 298934 165671 298962
rect 165699 298934 174485 298962
rect 174513 298934 174547 298962
rect 174575 298934 174609 298962
rect 174637 298934 174671 298962
rect 174699 298934 183485 298962
rect 183513 298934 183547 298962
rect 183575 298934 183609 298962
rect 183637 298934 183671 298962
rect 183699 298934 192485 298962
rect 192513 298934 192547 298962
rect 192575 298934 192609 298962
rect 192637 298934 192671 298962
rect 192699 298934 201485 298962
rect 201513 298934 201547 298962
rect 201575 298934 201609 298962
rect 201637 298934 201671 298962
rect 201699 298934 210485 298962
rect 210513 298934 210547 298962
rect 210575 298934 210609 298962
rect 210637 298934 210671 298962
rect 210699 298934 219485 298962
rect 219513 298934 219547 298962
rect 219575 298934 219609 298962
rect 219637 298934 219671 298962
rect 219699 298934 228485 298962
rect 228513 298934 228547 298962
rect 228575 298934 228609 298962
rect 228637 298934 228671 298962
rect 228699 298934 237485 298962
rect 237513 298934 237547 298962
rect 237575 298934 237609 298962
rect 237637 298934 237671 298962
rect 237699 298934 246485 298962
rect 246513 298934 246547 298962
rect 246575 298934 246609 298962
rect 246637 298934 246671 298962
rect 246699 298934 255485 298962
rect 255513 298934 255547 298962
rect 255575 298934 255609 298962
rect 255637 298934 255671 298962
rect 255699 298934 264485 298962
rect 264513 298934 264547 298962
rect 264575 298934 264609 298962
rect 264637 298934 264671 298962
rect 264699 298934 273485 298962
rect 273513 298934 273547 298962
rect 273575 298934 273609 298962
rect 273637 298934 273671 298962
rect 273699 298934 282485 298962
rect 282513 298934 282547 298962
rect 282575 298934 282609 298962
rect 282637 298934 282671 298962
rect 282699 298934 291485 298962
rect 291513 298934 291547 298962
rect 291575 298934 291609 298962
rect 291637 298934 291671 298962
rect 291699 298934 298728 298962
rect 298756 298934 298790 298962
rect 298818 298934 298852 298962
rect 298880 298934 298914 298962
rect 298942 298934 298990 298962
rect -958 298900 298990 298934
rect -958 298872 -910 298900
rect -882 298872 -848 298900
rect -820 298872 -786 298900
rect -758 298872 -724 298900
rect -696 298872 3485 298900
rect 3513 298872 3547 298900
rect 3575 298872 3609 298900
rect 3637 298872 3671 298900
rect 3699 298872 12485 298900
rect 12513 298872 12547 298900
rect 12575 298872 12609 298900
rect 12637 298872 12671 298900
rect 12699 298872 21485 298900
rect 21513 298872 21547 298900
rect 21575 298872 21609 298900
rect 21637 298872 21671 298900
rect 21699 298872 30485 298900
rect 30513 298872 30547 298900
rect 30575 298872 30609 298900
rect 30637 298872 30671 298900
rect 30699 298872 39485 298900
rect 39513 298872 39547 298900
rect 39575 298872 39609 298900
rect 39637 298872 39671 298900
rect 39699 298872 48485 298900
rect 48513 298872 48547 298900
rect 48575 298872 48609 298900
rect 48637 298872 48671 298900
rect 48699 298872 57485 298900
rect 57513 298872 57547 298900
rect 57575 298872 57609 298900
rect 57637 298872 57671 298900
rect 57699 298872 66485 298900
rect 66513 298872 66547 298900
rect 66575 298872 66609 298900
rect 66637 298872 66671 298900
rect 66699 298872 75485 298900
rect 75513 298872 75547 298900
rect 75575 298872 75609 298900
rect 75637 298872 75671 298900
rect 75699 298872 84485 298900
rect 84513 298872 84547 298900
rect 84575 298872 84609 298900
rect 84637 298872 84671 298900
rect 84699 298872 93485 298900
rect 93513 298872 93547 298900
rect 93575 298872 93609 298900
rect 93637 298872 93671 298900
rect 93699 298872 102485 298900
rect 102513 298872 102547 298900
rect 102575 298872 102609 298900
rect 102637 298872 102671 298900
rect 102699 298872 111485 298900
rect 111513 298872 111547 298900
rect 111575 298872 111609 298900
rect 111637 298872 111671 298900
rect 111699 298872 120485 298900
rect 120513 298872 120547 298900
rect 120575 298872 120609 298900
rect 120637 298872 120671 298900
rect 120699 298872 129485 298900
rect 129513 298872 129547 298900
rect 129575 298872 129609 298900
rect 129637 298872 129671 298900
rect 129699 298872 138485 298900
rect 138513 298872 138547 298900
rect 138575 298872 138609 298900
rect 138637 298872 138671 298900
rect 138699 298872 147485 298900
rect 147513 298872 147547 298900
rect 147575 298872 147609 298900
rect 147637 298872 147671 298900
rect 147699 298872 156485 298900
rect 156513 298872 156547 298900
rect 156575 298872 156609 298900
rect 156637 298872 156671 298900
rect 156699 298872 165485 298900
rect 165513 298872 165547 298900
rect 165575 298872 165609 298900
rect 165637 298872 165671 298900
rect 165699 298872 174485 298900
rect 174513 298872 174547 298900
rect 174575 298872 174609 298900
rect 174637 298872 174671 298900
rect 174699 298872 183485 298900
rect 183513 298872 183547 298900
rect 183575 298872 183609 298900
rect 183637 298872 183671 298900
rect 183699 298872 192485 298900
rect 192513 298872 192547 298900
rect 192575 298872 192609 298900
rect 192637 298872 192671 298900
rect 192699 298872 201485 298900
rect 201513 298872 201547 298900
rect 201575 298872 201609 298900
rect 201637 298872 201671 298900
rect 201699 298872 210485 298900
rect 210513 298872 210547 298900
rect 210575 298872 210609 298900
rect 210637 298872 210671 298900
rect 210699 298872 219485 298900
rect 219513 298872 219547 298900
rect 219575 298872 219609 298900
rect 219637 298872 219671 298900
rect 219699 298872 228485 298900
rect 228513 298872 228547 298900
rect 228575 298872 228609 298900
rect 228637 298872 228671 298900
rect 228699 298872 237485 298900
rect 237513 298872 237547 298900
rect 237575 298872 237609 298900
rect 237637 298872 237671 298900
rect 237699 298872 246485 298900
rect 246513 298872 246547 298900
rect 246575 298872 246609 298900
rect 246637 298872 246671 298900
rect 246699 298872 255485 298900
rect 255513 298872 255547 298900
rect 255575 298872 255609 298900
rect 255637 298872 255671 298900
rect 255699 298872 264485 298900
rect 264513 298872 264547 298900
rect 264575 298872 264609 298900
rect 264637 298872 264671 298900
rect 264699 298872 273485 298900
rect 273513 298872 273547 298900
rect 273575 298872 273609 298900
rect 273637 298872 273671 298900
rect 273699 298872 282485 298900
rect 282513 298872 282547 298900
rect 282575 298872 282609 298900
rect 282637 298872 282671 298900
rect 282699 298872 291485 298900
rect 291513 298872 291547 298900
rect 291575 298872 291609 298900
rect 291637 298872 291671 298900
rect 291699 298872 298728 298900
rect 298756 298872 298790 298900
rect 298818 298872 298852 298900
rect 298880 298872 298914 298900
rect 298942 298872 298990 298900
rect -958 298824 298990 298872
rect -478 298606 298510 298654
rect -478 298578 -430 298606
rect -402 298578 -368 298606
rect -340 298578 -306 298606
rect -278 298578 -244 298606
rect -216 298578 1625 298606
rect 1653 298578 1687 298606
rect 1715 298578 1749 298606
rect 1777 298578 1811 298606
rect 1839 298578 10625 298606
rect 10653 298578 10687 298606
rect 10715 298578 10749 298606
rect 10777 298578 10811 298606
rect 10839 298578 19625 298606
rect 19653 298578 19687 298606
rect 19715 298578 19749 298606
rect 19777 298578 19811 298606
rect 19839 298578 28625 298606
rect 28653 298578 28687 298606
rect 28715 298578 28749 298606
rect 28777 298578 28811 298606
rect 28839 298578 37625 298606
rect 37653 298578 37687 298606
rect 37715 298578 37749 298606
rect 37777 298578 37811 298606
rect 37839 298578 46625 298606
rect 46653 298578 46687 298606
rect 46715 298578 46749 298606
rect 46777 298578 46811 298606
rect 46839 298578 55625 298606
rect 55653 298578 55687 298606
rect 55715 298578 55749 298606
rect 55777 298578 55811 298606
rect 55839 298578 64625 298606
rect 64653 298578 64687 298606
rect 64715 298578 64749 298606
rect 64777 298578 64811 298606
rect 64839 298578 73625 298606
rect 73653 298578 73687 298606
rect 73715 298578 73749 298606
rect 73777 298578 73811 298606
rect 73839 298578 82625 298606
rect 82653 298578 82687 298606
rect 82715 298578 82749 298606
rect 82777 298578 82811 298606
rect 82839 298578 91625 298606
rect 91653 298578 91687 298606
rect 91715 298578 91749 298606
rect 91777 298578 91811 298606
rect 91839 298578 100625 298606
rect 100653 298578 100687 298606
rect 100715 298578 100749 298606
rect 100777 298578 100811 298606
rect 100839 298578 109625 298606
rect 109653 298578 109687 298606
rect 109715 298578 109749 298606
rect 109777 298578 109811 298606
rect 109839 298578 118625 298606
rect 118653 298578 118687 298606
rect 118715 298578 118749 298606
rect 118777 298578 118811 298606
rect 118839 298578 127625 298606
rect 127653 298578 127687 298606
rect 127715 298578 127749 298606
rect 127777 298578 127811 298606
rect 127839 298578 136625 298606
rect 136653 298578 136687 298606
rect 136715 298578 136749 298606
rect 136777 298578 136811 298606
rect 136839 298578 145625 298606
rect 145653 298578 145687 298606
rect 145715 298578 145749 298606
rect 145777 298578 145811 298606
rect 145839 298578 154625 298606
rect 154653 298578 154687 298606
rect 154715 298578 154749 298606
rect 154777 298578 154811 298606
rect 154839 298578 163625 298606
rect 163653 298578 163687 298606
rect 163715 298578 163749 298606
rect 163777 298578 163811 298606
rect 163839 298578 172625 298606
rect 172653 298578 172687 298606
rect 172715 298578 172749 298606
rect 172777 298578 172811 298606
rect 172839 298578 181625 298606
rect 181653 298578 181687 298606
rect 181715 298578 181749 298606
rect 181777 298578 181811 298606
rect 181839 298578 190625 298606
rect 190653 298578 190687 298606
rect 190715 298578 190749 298606
rect 190777 298578 190811 298606
rect 190839 298578 199625 298606
rect 199653 298578 199687 298606
rect 199715 298578 199749 298606
rect 199777 298578 199811 298606
rect 199839 298578 208625 298606
rect 208653 298578 208687 298606
rect 208715 298578 208749 298606
rect 208777 298578 208811 298606
rect 208839 298578 217625 298606
rect 217653 298578 217687 298606
rect 217715 298578 217749 298606
rect 217777 298578 217811 298606
rect 217839 298578 226625 298606
rect 226653 298578 226687 298606
rect 226715 298578 226749 298606
rect 226777 298578 226811 298606
rect 226839 298578 235625 298606
rect 235653 298578 235687 298606
rect 235715 298578 235749 298606
rect 235777 298578 235811 298606
rect 235839 298578 244625 298606
rect 244653 298578 244687 298606
rect 244715 298578 244749 298606
rect 244777 298578 244811 298606
rect 244839 298578 253625 298606
rect 253653 298578 253687 298606
rect 253715 298578 253749 298606
rect 253777 298578 253811 298606
rect 253839 298578 262625 298606
rect 262653 298578 262687 298606
rect 262715 298578 262749 298606
rect 262777 298578 262811 298606
rect 262839 298578 271625 298606
rect 271653 298578 271687 298606
rect 271715 298578 271749 298606
rect 271777 298578 271811 298606
rect 271839 298578 280625 298606
rect 280653 298578 280687 298606
rect 280715 298578 280749 298606
rect 280777 298578 280811 298606
rect 280839 298578 289625 298606
rect 289653 298578 289687 298606
rect 289715 298578 289749 298606
rect 289777 298578 289811 298606
rect 289839 298578 298248 298606
rect 298276 298578 298310 298606
rect 298338 298578 298372 298606
rect 298400 298578 298434 298606
rect 298462 298578 298510 298606
rect -478 298544 298510 298578
rect -478 298516 -430 298544
rect -402 298516 -368 298544
rect -340 298516 -306 298544
rect -278 298516 -244 298544
rect -216 298516 1625 298544
rect 1653 298516 1687 298544
rect 1715 298516 1749 298544
rect 1777 298516 1811 298544
rect 1839 298516 10625 298544
rect 10653 298516 10687 298544
rect 10715 298516 10749 298544
rect 10777 298516 10811 298544
rect 10839 298516 19625 298544
rect 19653 298516 19687 298544
rect 19715 298516 19749 298544
rect 19777 298516 19811 298544
rect 19839 298516 28625 298544
rect 28653 298516 28687 298544
rect 28715 298516 28749 298544
rect 28777 298516 28811 298544
rect 28839 298516 37625 298544
rect 37653 298516 37687 298544
rect 37715 298516 37749 298544
rect 37777 298516 37811 298544
rect 37839 298516 46625 298544
rect 46653 298516 46687 298544
rect 46715 298516 46749 298544
rect 46777 298516 46811 298544
rect 46839 298516 55625 298544
rect 55653 298516 55687 298544
rect 55715 298516 55749 298544
rect 55777 298516 55811 298544
rect 55839 298516 64625 298544
rect 64653 298516 64687 298544
rect 64715 298516 64749 298544
rect 64777 298516 64811 298544
rect 64839 298516 73625 298544
rect 73653 298516 73687 298544
rect 73715 298516 73749 298544
rect 73777 298516 73811 298544
rect 73839 298516 82625 298544
rect 82653 298516 82687 298544
rect 82715 298516 82749 298544
rect 82777 298516 82811 298544
rect 82839 298516 91625 298544
rect 91653 298516 91687 298544
rect 91715 298516 91749 298544
rect 91777 298516 91811 298544
rect 91839 298516 100625 298544
rect 100653 298516 100687 298544
rect 100715 298516 100749 298544
rect 100777 298516 100811 298544
rect 100839 298516 109625 298544
rect 109653 298516 109687 298544
rect 109715 298516 109749 298544
rect 109777 298516 109811 298544
rect 109839 298516 118625 298544
rect 118653 298516 118687 298544
rect 118715 298516 118749 298544
rect 118777 298516 118811 298544
rect 118839 298516 127625 298544
rect 127653 298516 127687 298544
rect 127715 298516 127749 298544
rect 127777 298516 127811 298544
rect 127839 298516 136625 298544
rect 136653 298516 136687 298544
rect 136715 298516 136749 298544
rect 136777 298516 136811 298544
rect 136839 298516 145625 298544
rect 145653 298516 145687 298544
rect 145715 298516 145749 298544
rect 145777 298516 145811 298544
rect 145839 298516 154625 298544
rect 154653 298516 154687 298544
rect 154715 298516 154749 298544
rect 154777 298516 154811 298544
rect 154839 298516 163625 298544
rect 163653 298516 163687 298544
rect 163715 298516 163749 298544
rect 163777 298516 163811 298544
rect 163839 298516 172625 298544
rect 172653 298516 172687 298544
rect 172715 298516 172749 298544
rect 172777 298516 172811 298544
rect 172839 298516 181625 298544
rect 181653 298516 181687 298544
rect 181715 298516 181749 298544
rect 181777 298516 181811 298544
rect 181839 298516 190625 298544
rect 190653 298516 190687 298544
rect 190715 298516 190749 298544
rect 190777 298516 190811 298544
rect 190839 298516 199625 298544
rect 199653 298516 199687 298544
rect 199715 298516 199749 298544
rect 199777 298516 199811 298544
rect 199839 298516 208625 298544
rect 208653 298516 208687 298544
rect 208715 298516 208749 298544
rect 208777 298516 208811 298544
rect 208839 298516 217625 298544
rect 217653 298516 217687 298544
rect 217715 298516 217749 298544
rect 217777 298516 217811 298544
rect 217839 298516 226625 298544
rect 226653 298516 226687 298544
rect 226715 298516 226749 298544
rect 226777 298516 226811 298544
rect 226839 298516 235625 298544
rect 235653 298516 235687 298544
rect 235715 298516 235749 298544
rect 235777 298516 235811 298544
rect 235839 298516 244625 298544
rect 244653 298516 244687 298544
rect 244715 298516 244749 298544
rect 244777 298516 244811 298544
rect 244839 298516 253625 298544
rect 253653 298516 253687 298544
rect 253715 298516 253749 298544
rect 253777 298516 253811 298544
rect 253839 298516 262625 298544
rect 262653 298516 262687 298544
rect 262715 298516 262749 298544
rect 262777 298516 262811 298544
rect 262839 298516 271625 298544
rect 271653 298516 271687 298544
rect 271715 298516 271749 298544
rect 271777 298516 271811 298544
rect 271839 298516 280625 298544
rect 280653 298516 280687 298544
rect 280715 298516 280749 298544
rect 280777 298516 280811 298544
rect 280839 298516 289625 298544
rect 289653 298516 289687 298544
rect 289715 298516 289749 298544
rect 289777 298516 289811 298544
rect 289839 298516 298248 298544
rect 298276 298516 298310 298544
rect 298338 298516 298372 298544
rect 298400 298516 298434 298544
rect 298462 298516 298510 298544
rect -478 298482 298510 298516
rect -478 298454 -430 298482
rect -402 298454 -368 298482
rect -340 298454 -306 298482
rect -278 298454 -244 298482
rect -216 298454 1625 298482
rect 1653 298454 1687 298482
rect 1715 298454 1749 298482
rect 1777 298454 1811 298482
rect 1839 298454 10625 298482
rect 10653 298454 10687 298482
rect 10715 298454 10749 298482
rect 10777 298454 10811 298482
rect 10839 298454 19625 298482
rect 19653 298454 19687 298482
rect 19715 298454 19749 298482
rect 19777 298454 19811 298482
rect 19839 298454 28625 298482
rect 28653 298454 28687 298482
rect 28715 298454 28749 298482
rect 28777 298454 28811 298482
rect 28839 298454 37625 298482
rect 37653 298454 37687 298482
rect 37715 298454 37749 298482
rect 37777 298454 37811 298482
rect 37839 298454 46625 298482
rect 46653 298454 46687 298482
rect 46715 298454 46749 298482
rect 46777 298454 46811 298482
rect 46839 298454 55625 298482
rect 55653 298454 55687 298482
rect 55715 298454 55749 298482
rect 55777 298454 55811 298482
rect 55839 298454 64625 298482
rect 64653 298454 64687 298482
rect 64715 298454 64749 298482
rect 64777 298454 64811 298482
rect 64839 298454 73625 298482
rect 73653 298454 73687 298482
rect 73715 298454 73749 298482
rect 73777 298454 73811 298482
rect 73839 298454 82625 298482
rect 82653 298454 82687 298482
rect 82715 298454 82749 298482
rect 82777 298454 82811 298482
rect 82839 298454 91625 298482
rect 91653 298454 91687 298482
rect 91715 298454 91749 298482
rect 91777 298454 91811 298482
rect 91839 298454 100625 298482
rect 100653 298454 100687 298482
rect 100715 298454 100749 298482
rect 100777 298454 100811 298482
rect 100839 298454 109625 298482
rect 109653 298454 109687 298482
rect 109715 298454 109749 298482
rect 109777 298454 109811 298482
rect 109839 298454 118625 298482
rect 118653 298454 118687 298482
rect 118715 298454 118749 298482
rect 118777 298454 118811 298482
rect 118839 298454 127625 298482
rect 127653 298454 127687 298482
rect 127715 298454 127749 298482
rect 127777 298454 127811 298482
rect 127839 298454 136625 298482
rect 136653 298454 136687 298482
rect 136715 298454 136749 298482
rect 136777 298454 136811 298482
rect 136839 298454 145625 298482
rect 145653 298454 145687 298482
rect 145715 298454 145749 298482
rect 145777 298454 145811 298482
rect 145839 298454 154625 298482
rect 154653 298454 154687 298482
rect 154715 298454 154749 298482
rect 154777 298454 154811 298482
rect 154839 298454 163625 298482
rect 163653 298454 163687 298482
rect 163715 298454 163749 298482
rect 163777 298454 163811 298482
rect 163839 298454 172625 298482
rect 172653 298454 172687 298482
rect 172715 298454 172749 298482
rect 172777 298454 172811 298482
rect 172839 298454 181625 298482
rect 181653 298454 181687 298482
rect 181715 298454 181749 298482
rect 181777 298454 181811 298482
rect 181839 298454 190625 298482
rect 190653 298454 190687 298482
rect 190715 298454 190749 298482
rect 190777 298454 190811 298482
rect 190839 298454 199625 298482
rect 199653 298454 199687 298482
rect 199715 298454 199749 298482
rect 199777 298454 199811 298482
rect 199839 298454 208625 298482
rect 208653 298454 208687 298482
rect 208715 298454 208749 298482
rect 208777 298454 208811 298482
rect 208839 298454 217625 298482
rect 217653 298454 217687 298482
rect 217715 298454 217749 298482
rect 217777 298454 217811 298482
rect 217839 298454 226625 298482
rect 226653 298454 226687 298482
rect 226715 298454 226749 298482
rect 226777 298454 226811 298482
rect 226839 298454 235625 298482
rect 235653 298454 235687 298482
rect 235715 298454 235749 298482
rect 235777 298454 235811 298482
rect 235839 298454 244625 298482
rect 244653 298454 244687 298482
rect 244715 298454 244749 298482
rect 244777 298454 244811 298482
rect 244839 298454 253625 298482
rect 253653 298454 253687 298482
rect 253715 298454 253749 298482
rect 253777 298454 253811 298482
rect 253839 298454 262625 298482
rect 262653 298454 262687 298482
rect 262715 298454 262749 298482
rect 262777 298454 262811 298482
rect 262839 298454 271625 298482
rect 271653 298454 271687 298482
rect 271715 298454 271749 298482
rect 271777 298454 271811 298482
rect 271839 298454 280625 298482
rect 280653 298454 280687 298482
rect 280715 298454 280749 298482
rect 280777 298454 280811 298482
rect 280839 298454 289625 298482
rect 289653 298454 289687 298482
rect 289715 298454 289749 298482
rect 289777 298454 289811 298482
rect 289839 298454 298248 298482
rect 298276 298454 298310 298482
rect 298338 298454 298372 298482
rect 298400 298454 298434 298482
rect 298462 298454 298510 298482
rect -478 298420 298510 298454
rect -478 298392 -430 298420
rect -402 298392 -368 298420
rect -340 298392 -306 298420
rect -278 298392 -244 298420
rect -216 298392 1625 298420
rect 1653 298392 1687 298420
rect 1715 298392 1749 298420
rect 1777 298392 1811 298420
rect 1839 298392 10625 298420
rect 10653 298392 10687 298420
rect 10715 298392 10749 298420
rect 10777 298392 10811 298420
rect 10839 298392 19625 298420
rect 19653 298392 19687 298420
rect 19715 298392 19749 298420
rect 19777 298392 19811 298420
rect 19839 298392 28625 298420
rect 28653 298392 28687 298420
rect 28715 298392 28749 298420
rect 28777 298392 28811 298420
rect 28839 298392 37625 298420
rect 37653 298392 37687 298420
rect 37715 298392 37749 298420
rect 37777 298392 37811 298420
rect 37839 298392 46625 298420
rect 46653 298392 46687 298420
rect 46715 298392 46749 298420
rect 46777 298392 46811 298420
rect 46839 298392 55625 298420
rect 55653 298392 55687 298420
rect 55715 298392 55749 298420
rect 55777 298392 55811 298420
rect 55839 298392 64625 298420
rect 64653 298392 64687 298420
rect 64715 298392 64749 298420
rect 64777 298392 64811 298420
rect 64839 298392 73625 298420
rect 73653 298392 73687 298420
rect 73715 298392 73749 298420
rect 73777 298392 73811 298420
rect 73839 298392 82625 298420
rect 82653 298392 82687 298420
rect 82715 298392 82749 298420
rect 82777 298392 82811 298420
rect 82839 298392 91625 298420
rect 91653 298392 91687 298420
rect 91715 298392 91749 298420
rect 91777 298392 91811 298420
rect 91839 298392 100625 298420
rect 100653 298392 100687 298420
rect 100715 298392 100749 298420
rect 100777 298392 100811 298420
rect 100839 298392 109625 298420
rect 109653 298392 109687 298420
rect 109715 298392 109749 298420
rect 109777 298392 109811 298420
rect 109839 298392 118625 298420
rect 118653 298392 118687 298420
rect 118715 298392 118749 298420
rect 118777 298392 118811 298420
rect 118839 298392 127625 298420
rect 127653 298392 127687 298420
rect 127715 298392 127749 298420
rect 127777 298392 127811 298420
rect 127839 298392 136625 298420
rect 136653 298392 136687 298420
rect 136715 298392 136749 298420
rect 136777 298392 136811 298420
rect 136839 298392 145625 298420
rect 145653 298392 145687 298420
rect 145715 298392 145749 298420
rect 145777 298392 145811 298420
rect 145839 298392 154625 298420
rect 154653 298392 154687 298420
rect 154715 298392 154749 298420
rect 154777 298392 154811 298420
rect 154839 298392 163625 298420
rect 163653 298392 163687 298420
rect 163715 298392 163749 298420
rect 163777 298392 163811 298420
rect 163839 298392 172625 298420
rect 172653 298392 172687 298420
rect 172715 298392 172749 298420
rect 172777 298392 172811 298420
rect 172839 298392 181625 298420
rect 181653 298392 181687 298420
rect 181715 298392 181749 298420
rect 181777 298392 181811 298420
rect 181839 298392 190625 298420
rect 190653 298392 190687 298420
rect 190715 298392 190749 298420
rect 190777 298392 190811 298420
rect 190839 298392 199625 298420
rect 199653 298392 199687 298420
rect 199715 298392 199749 298420
rect 199777 298392 199811 298420
rect 199839 298392 208625 298420
rect 208653 298392 208687 298420
rect 208715 298392 208749 298420
rect 208777 298392 208811 298420
rect 208839 298392 217625 298420
rect 217653 298392 217687 298420
rect 217715 298392 217749 298420
rect 217777 298392 217811 298420
rect 217839 298392 226625 298420
rect 226653 298392 226687 298420
rect 226715 298392 226749 298420
rect 226777 298392 226811 298420
rect 226839 298392 235625 298420
rect 235653 298392 235687 298420
rect 235715 298392 235749 298420
rect 235777 298392 235811 298420
rect 235839 298392 244625 298420
rect 244653 298392 244687 298420
rect 244715 298392 244749 298420
rect 244777 298392 244811 298420
rect 244839 298392 253625 298420
rect 253653 298392 253687 298420
rect 253715 298392 253749 298420
rect 253777 298392 253811 298420
rect 253839 298392 262625 298420
rect 262653 298392 262687 298420
rect 262715 298392 262749 298420
rect 262777 298392 262811 298420
rect 262839 298392 271625 298420
rect 271653 298392 271687 298420
rect 271715 298392 271749 298420
rect 271777 298392 271811 298420
rect 271839 298392 280625 298420
rect 280653 298392 280687 298420
rect 280715 298392 280749 298420
rect 280777 298392 280811 298420
rect 280839 298392 289625 298420
rect 289653 298392 289687 298420
rect 289715 298392 289749 298420
rect 289777 298392 289811 298420
rect 289839 298392 298248 298420
rect 298276 298392 298310 298420
rect 298338 298392 298372 298420
rect 298400 298392 298434 298420
rect 298462 298392 298510 298420
rect -478 298344 298510 298392
rect -958 293175 298990 293223
rect -958 293147 -910 293175
rect -882 293147 -848 293175
rect -820 293147 -786 293175
rect -758 293147 -724 293175
rect -696 293147 3485 293175
rect 3513 293147 3547 293175
rect 3575 293147 3609 293175
rect 3637 293147 3671 293175
rect 3699 293147 12485 293175
rect 12513 293147 12547 293175
rect 12575 293147 12609 293175
rect 12637 293147 12671 293175
rect 12699 293147 21485 293175
rect 21513 293147 21547 293175
rect 21575 293147 21609 293175
rect 21637 293147 21671 293175
rect 21699 293147 30485 293175
rect 30513 293147 30547 293175
rect 30575 293147 30609 293175
rect 30637 293147 30671 293175
rect 30699 293147 39485 293175
rect 39513 293147 39547 293175
rect 39575 293147 39609 293175
rect 39637 293147 39671 293175
rect 39699 293147 48485 293175
rect 48513 293147 48547 293175
rect 48575 293147 48609 293175
rect 48637 293147 48671 293175
rect 48699 293147 57485 293175
rect 57513 293147 57547 293175
rect 57575 293147 57609 293175
rect 57637 293147 57671 293175
rect 57699 293147 66485 293175
rect 66513 293147 66547 293175
rect 66575 293147 66609 293175
rect 66637 293147 66671 293175
rect 66699 293147 75485 293175
rect 75513 293147 75547 293175
rect 75575 293147 75609 293175
rect 75637 293147 75671 293175
rect 75699 293147 84485 293175
rect 84513 293147 84547 293175
rect 84575 293147 84609 293175
rect 84637 293147 84671 293175
rect 84699 293147 93485 293175
rect 93513 293147 93547 293175
rect 93575 293147 93609 293175
rect 93637 293147 93671 293175
rect 93699 293147 102485 293175
rect 102513 293147 102547 293175
rect 102575 293147 102609 293175
rect 102637 293147 102671 293175
rect 102699 293147 111485 293175
rect 111513 293147 111547 293175
rect 111575 293147 111609 293175
rect 111637 293147 111671 293175
rect 111699 293147 120485 293175
rect 120513 293147 120547 293175
rect 120575 293147 120609 293175
rect 120637 293147 120671 293175
rect 120699 293147 129485 293175
rect 129513 293147 129547 293175
rect 129575 293147 129609 293175
rect 129637 293147 129671 293175
rect 129699 293147 138485 293175
rect 138513 293147 138547 293175
rect 138575 293147 138609 293175
rect 138637 293147 138671 293175
rect 138699 293147 147485 293175
rect 147513 293147 147547 293175
rect 147575 293147 147609 293175
rect 147637 293147 147671 293175
rect 147699 293147 156485 293175
rect 156513 293147 156547 293175
rect 156575 293147 156609 293175
rect 156637 293147 156671 293175
rect 156699 293147 165485 293175
rect 165513 293147 165547 293175
rect 165575 293147 165609 293175
rect 165637 293147 165671 293175
rect 165699 293147 174485 293175
rect 174513 293147 174547 293175
rect 174575 293147 174609 293175
rect 174637 293147 174671 293175
rect 174699 293147 183485 293175
rect 183513 293147 183547 293175
rect 183575 293147 183609 293175
rect 183637 293147 183671 293175
rect 183699 293147 192485 293175
rect 192513 293147 192547 293175
rect 192575 293147 192609 293175
rect 192637 293147 192671 293175
rect 192699 293147 201485 293175
rect 201513 293147 201547 293175
rect 201575 293147 201609 293175
rect 201637 293147 201671 293175
rect 201699 293147 210485 293175
rect 210513 293147 210547 293175
rect 210575 293147 210609 293175
rect 210637 293147 210671 293175
rect 210699 293147 219485 293175
rect 219513 293147 219547 293175
rect 219575 293147 219609 293175
rect 219637 293147 219671 293175
rect 219699 293147 228485 293175
rect 228513 293147 228547 293175
rect 228575 293147 228609 293175
rect 228637 293147 228671 293175
rect 228699 293147 237485 293175
rect 237513 293147 237547 293175
rect 237575 293147 237609 293175
rect 237637 293147 237671 293175
rect 237699 293147 246485 293175
rect 246513 293147 246547 293175
rect 246575 293147 246609 293175
rect 246637 293147 246671 293175
rect 246699 293147 255485 293175
rect 255513 293147 255547 293175
rect 255575 293147 255609 293175
rect 255637 293147 255671 293175
rect 255699 293147 264485 293175
rect 264513 293147 264547 293175
rect 264575 293147 264609 293175
rect 264637 293147 264671 293175
rect 264699 293147 273485 293175
rect 273513 293147 273547 293175
rect 273575 293147 273609 293175
rect 273637 293147 273671 293175
rect 273699 293147 282485 293175
rect 282513 293147 282547 293175
rect 282575 293147 282609 293175
rect 282637 293147 282671 293175
rect 282699 293147 291485 293175
rect 291513 293147 291547 293175
rect 291575 293147 291609 293175
rect 291637 293147 291671 293175
rect 291699 293147 298728 293175
rect 298756 293147 298790 293175
rect 298818 293147 298852 293175
rect 298880 293147 298914 293175
rect 298942 293147 298990 293175
rect -958 293113 298990 293147
rect -958 293085 -910 293113
rect -882 293085 -848 293113
rect -820 293085 -786 293113
rect -758 293085 -724 293113
rect -696 293085 3485 293113
rect 3513 293085 3547 293113
rect 3575 293085 3609 293113
rect 3637 293085 3671 293113
rect 3699 293085 12485 293113
rect 12513 293085 12547 293113
rect 12575 293085 12609 293113
rect 12637 293085 12671 293113
rect 12699 293085 21485 293113
rect 21513 293085 21547 293113
rect 21575 293085 21609 293113
rect 21637 293085 21671 293113
rect 21699 293085 30485 293113
rect 30513 293085 30547 293113
rect 30575 293085 30609 293113
rect 30637 293085 30671 293113
rect 30699 293085 39485 293113
rect 39513 293085 39547 293113
rect 39575 293085 39609 293113
rect 39637 293085 39671 293113
rect 39699 293085 48485 293113
rect 48513 293085 48547 293113
rect 48575 293085 48609 293113
rect 48637 293085 48671 293113
rect 48699 293085 57485 293113
rect 57513 293085 57547 293113
rect 57575 293085 57609 293113
rect 57637 293085 57671 293113
rect 57699 293085 66485 293113
rect 66513 293085 66547 293113
rect 66575 293085 66609 293113
rect 66637 293085 66671 293113
rect 66699 293085 75485 293113
rect 75513 293085 75547 293113
rect 75575 293085 75609 293113
rect 75637 293085 75671 293113
rect 75699 293085 84485 293113
rect 84513 293085 84547 293113
rect 84575 293085 84609 293113
rect 84637 293085 84671 293113
rect 84699 293085 93485 293113
rect 93513 293085 93547 293113
rect 93575 293085 93609 293113
rect 93637 293085 93671 293113
rect 93699 293085 102485 293113
rect 102513 293085 102547 293113
rect 102575 293085 102609 293113
rect 102637 293085 102671 293113
rect 102699 293085 111485 293113
rect 111513 293085 111547 293113
rect 111575 293085 111609 293113
rect 111637 293085 111671 293113
rect 111699 293085 120485 293113
rect 120513 293085 120547 293113
rect 120575 293085 120609 293113
rect 120637 293085 120671 293113
rect 120699 293085 129485 293113
rect 129513 293085 129547 293113
rect 129575 293085 129609 293113
rect 129637 293085 129671 293113
rect 129699 293085 138485 293113
rect 138513 293085 138547 293113
rect 138575 293085 138609 293113
rect 138637 293085 138671 293113
rect 138699 293085 147485 293113
rect 147513 293085 147547 293113
rect 147575 293085 147609 293113
rect 147637 293085 147671 293113
rect 147699 293085 156485 293113
rect 156513 293085 156547 293113
rect 156575 293085 156609 293113
rect 156637 293085 156671 293113
rect 156699 293085 165485 293113
rect 165513 293085 165547 293113
rect 165575 293085 165609 293113
rect 165637 293085 165671 293113
rect 165699 293085 174485 293113
rect 174513 293085 174547 293113
rect 174575 293085 174609 293113
rect 174637 293085 174671 293113
rect 174699 293085 183485 293113
rect 183513 293085 183547 293113
rect 183575 293085 183609 293113
rect 183637 293085 183671 293113
rect 183699 293085 192485 293113
rect 192513 293085 192547 293113
rect 192575 293085 192609 293113
rect 192637 293085 192671 293113
rect 192699 293085 201485 293113
rect 201513 293085 201547 293113
rect 201575 293085 201609 293113
rect 201637 293085 201671 293113
rect 201699 293085 210485 293113
rect 210513 293085 210547 293113
rect 210575 293085 210609 293113
rect 210637 293085 210671 293113
rect 210699 293085 219485 293113
rect 219513 293085 219547 293113
rect 219575 293085 219609 293113
rect 219637 293085 219671 293113
rect 219699 293085 228485 293113
rect 228513 293085 228547 293113
rect 228575 293085 228609 293113
rect 228637 293085 228671 293113
rect 228699 293085 237485 293113
rect 237513 293085 237547 293113
rect 237575 293085 237609 293113
rect 237637 293085 237671 293113
rect 237699 293085 246485 293113
rect 246513 293085 246547 293113
rect 246575 293085 246609 293113
rect 246637 293085 246671 293113
rect 246699 293085 255485 293113
rect 255513 293085 255547 293113
rect 255575 293085 255609 293113
rect 255637 293085 255671 293113
rect 255699 293085 264485 293113
rect 264513 293085 264547 293113
rect 264575 293085 264609 293113
rect 264637 293085 264671 293113
rect 264699 293085 273485 293113
rect 273513 293085 273547 293113
rect 273575 293085 273609 293113
rect 273637 293085 273671 293113
rect 273699 293085 282485 293113
rect 282513 293085 282547 293113
rect 282575 293085 282609 293113
rect 282637 293085 282671 293113
rect 282699 293085 291485 293113
rect 291513 293085 291547 293113
rect 291575 293085 291609 293113
rect 291637 293085 291671 293113
rect 291699 293085 298728 293113
rect 298756 293085 298790 293113
rect 298818 293085 298852 293113
rect 298880 293085 298914 293113
rect 298942 293085 298990 293113
rect -958 293051 298990 293085
rect -958 293023 -910 293051
rect -882 293023 -848 293051
rect -820 293023 -786 293051
rect -758 293023 -724 293051
rect -696 293023 3485 293051
rect 3513 293023 3547 293051
rect 3575 293023 3609 293051
rect 3637 293023 3671 293051
rect 3699 293023 12485 293051
rect 12513 293023 12547 293051
rect 12575 293023 12609 293051
rect 12637 293023 12671 293051
rect 12699 293023 21485 293051
rect 21513 293023 21547 293051
rect 21575 293023 21609 293051
rect 21637 293023 21671 293051
rect 21699 293023 30485 293051
rect 30513 293023 30547 293051
rect 30575 293023 30609 293051
rect 30637 293023 30671 293051
rect 30699 293023 39485 293051
rect 39513 293023 39547 293051
rect 39575 293023 39609 293051
rect 39637 293023 39671 293051
rect 39699 293023 48485 293051
rect 48513 293023 48547 293051
rect 48575 293023 48609 293051
rect 48637 293023 48671 293051
rect 48699 293023 57485 293051
rect 57513 293023 57547 293051
rect 57575 293023 57609 293051
rect 57637 293023 57671 293051
rect 57699 293023 66485 293051
rect 66513 293023 66547 293051
rect 66575 293023 66609 293051
rect 66637 293023 66671 293051
rect 66699 293023 75485 293051
rect 75513 293023 75547 293051
rect 75575 293023 75609 293051
rect 75637 293023 75671 293051
rect 75699 293023 84485 293051
rect 84513 293023 84547 293051
rect 84575 293023 84609 293051
rect 84637 293023 84671 293051
rect 84699 293023 93485 293051
rect 93513 293023 93547 293051
rect 93575 293023 93609 293051
rect 93637 293023 93671 293051
rect 93699 293023 102485 293051
rect 102513 293023 102547 293051
rect 102575 293023 102609 293051
rect 102637 293023 102671 293051
rect 102699 293023 111485 293051
rect 111513 293023 111547 293051
rect 111575 293023 111609 293051
rect 111637 293023 111671 293051
rect 111699 293023 120485 293051
rect 120513 293023 120547 293051
rect 120575 293023 120609 293051
rect 120637 293023 120671 293051
rect 120699 293023 129485 293051
rect 129513 293023 129547 293051
rect 129575 293023 129609 293051
rect 129637 293023 129671 293051
rect 129699 293023 138485 293051
rect 138513 293023 138547 293051
rect 138575 293023 138609 293051
rect 138637 293023 138671 293051
rect 138699 293023 147485 293051
rect 147513 293023 147547 293051
rect 147575 293023 147609 293051
rect 147637 293023 147671 293051
rect 147699 293023 156485 293051
rect 156513 293023 156547 293051
rect 156575 293023 156609 293051
rect 156637 293023 156671 293051
rect 156699 293023 165485 293051
rect 165513 293023 165547 293051
rect 165575 293023 165609 293051
rect 165637 293023 165671 293051
rect 165699 293023 174485 293051
rect 174513 293023 174547 293051
rect 174575 293023 174609 293051
rect 174637 293023 174671 293051
rect 174699 293023 183485 293051
rect 183513 293023 183547 293051
rect 183575 293023 183609 293051
rect 183637 293023 183671 293051
rect 183699 293023 192485 293051
rect 192513 293023 192547 293051
rect 192575 293023 192609 293051
rect 192637 293023 192671 293051
rect 192699 293023 201485 293051
rect 201513 293023 201547 293051
rect 201575 293023 201609 293051
rect 201637 293023 201671 293051
rect 201699 293023 210485 293051
rect 210513 293023 210547 293051
rect 210575 293023 210609 293051
rect 210637 293023 210671 293051
rect 210699 293023 219485 293051
rect 219513 293023 219547 293051
rect 219575 293023 219609 293051
rect 219637 293023 219671 293051
rect 219699 293023 228485 293051
rect 228513 293023 228547 293051
rect 228575 293023 228609 293051
rect 228637 293023 228671 293051
rect 228699 293023 237485 293051
rect 237513 293023 237547 293051
rect 237575 293023 237609 293051
rect 237637 293023 237671 293051
rect 237699 293023 246485 293051
rect 246513 293023 246547 293051
rect 246575 293023 246609 293051
rect 246637 293023 246671 293051
rect 246699 293023 255485 293051
rect 255513 293023 255547 293051
rect 255575 293023 255609 293051
rect 255637 293023 255671 293051
rect 255699 293023 264485 293051
rect 264513 293023 264547 293051
rect 264575 293023 264609 293051
rect 264637 293023 264671 293051
rect 264699 293023 273485 293051
rect 273513 293023 273547 293051
rect 273575 293023 273609 293051
rect 273637 293023 273671 293051
rect 273699 293023 282485 293051
rect 282513 293023 282547 293051
rect 282575 293023 282609 293051
rect 282637 293023 282671 293051
rect 282699 293023 291485 293051
rect 291513 293023 291547 293051
rect 291575 293023 291609 293051
rect 291637 293023 291671 293051
rect 291699 293023 298728 293051
rect 298756 293023 298790 293051
rect 298818 293023 298852 293051
rect 298880 293023 298914 293051
rect 298942 293023 298990 293051
rect -958 292989 298990 293023
rect -958 292961 -910 292989
rect -882 292961 -848 292989
rect -820 292961 -786 292989
rect -758 292961 -724 292989
rect -696 292961 3485 292989
rect 3513 292961 3547 292989
rect 3575 292961 3609 292989
rect 3637 292961 3671 292989
rect 3699 292961 12485 292989
rect 12513 292961 12547 292989
rect 12575 292961 12609 292989
rect 12637 292961 12671 292989
rect 12699 292961 21485 292989
rect 21513 292961 21547 292989
rect 21575 292961 21609 292989
rect 21637 292961 21671 292989
rect 21699 292961 30485 292989
rect 30513 292961 30547 292989
rect 30575 292961 30609 292989
rect 30637 292961 30671 292989
rect 30699 292961 39485 292989
rect 39513 292961 39547 292989
rect 39575 292961 39609 292989
rect 39637 292961 39671 292989
rect 39699 292961 48485 292989
rect 48513 292961 48547 292989
rect 48575 292961 48609 292989
rect 48637 292961 48671 292989
rect 48699 292961 57485 292989
rect 57513 292961 57547 292989
rect 57575 292961 57609 292989
rect 57637 292961 57671 292989
rect 57699 292961 66485 292989
rect 66513 292961 66547 292989
rect 66575 292961 66609 292989
rect 66637 292961 66671 292989
rect 66699 292961 75485 292989
rect 75513 292961 75547 292989
rect 75575 292961 75609 292989
rect 75637 292961 75671 292989
rect 75699 292961 84485 292989
rect 84513 292961 84547 292989
rect 84575 292961 84609 292989
rect 84637 292961 84671 292989
rect 84699 292961 93485 292989
rect 93513 292961 93547 292989
rect 93575 292961 93609 292989
rect 93637 292961 93671 292989
rect 93699 292961 102485 292989
rect 102513 292961 102547 292989
rect 102575 292961 102609 292989
rect 102637 292961 102671 292989
rect 102699 292961 111485 292989
rect 111513 292961 111547 292989
rect 111575 292961 111609 292989
rect 111637 292961 111671 292989
rect 111699 292961 120485 292989
rect 120513 292961 120547 292989
rect 120575 292961 120609 292989
rect 120637 292961 120671 292989
rect 120699 292961 129485 292989
rect 129513 292961 129547 292989
rect 129575 292961 129609 292989
rect 129637 292961 129671 292989
rect 129699 292961 138485 292989
rect 138513 292961 138547 292989
rect 138575 292961 138609 292989
rect 138637 292961 138671 292989
rect 138699 292961 147485 292989
rect 147513 292961 147547 292989
rect 147575 292961 147609 292989
rect 147637 292961 147671 292989
rect 147699 292961 156485 292989
rect 156513 292961 156547 292989
rect 156575 292961 156609 292989
rect 156637 292961 156671 292989
rect 156699 292961 165485 292989
rect 165513 292961 165547 292989
rect 165575 292961 165609 292989
rect 165637 292961 165671 292989
rect 165699 292961 174485 292989
rect 174513 292961 174547 292989
rect 174575 292961 174609 292989
rect 174637 292961 174671 292989
rect 174699 292961 183485 292989
rect 183513 292961 183547 292989
rect 183575 292961 183609 292989
rect 183637 292961 183671 292989
rect 183699 292961 192485 292989
rect 192513 292961 192547 292989
rect 192575 292961 192609 292989
rect 192637 292961 192671 292989
rect 192699 292961 201485 292989
rect 201513 292961 201547 292989
rect 201575 292961 201609 292989
rect 201637 292961 201671 292989
rect 201699 292961 210485 292989
rect 210513 292961 210547 292989
rect 210575 292961 210609 292989
rect 210637 292961 210671 292989
rect 210699 292961 219485 292989
rect 219513 292961 219547 292989
rect 219575 292961 219609 292989
rect 219637 292961 219671 292989
rect 219699 292961 228485 292989
rect 228513 292961 228547 292989
rect 228575 292961 228609 292989
rect 228637 292961 228671 292989
rect 228699 292961 237485 292989
rect 237513 292961 237547 292989
rect 237575 292961 237609 292989
rect 237637 292961 237671 292989
rect 237699 292961 246485 292989
rect 246513 292961 246547 292989
rect 246575 292961 246609 292989
rect 246637 292961 246671 292989
rect 246699 292961 255485 292989
rect 255513 292961 255547 292989
rect 255575 292961 255609 292989
rect 255637 292961 255671 292989
rect 255699 292961 264485 292989
rect 264513 292961 264547 292989
rect 264575 292961 264609 292989
rect 264637 292961 264671 292989
rect 264699 292961 273485 292989
rect 273513 292961 273547 292989
rect 273575 292961 273609 292989
rect 273637 292961 273671 292989
rect 273699 292961 282485 292989
rect 282513 292961 282547 292989
rect 282575 292961 282609 292989
rect 282637 292961 282671 292989
rect 282699 292961 291485 292989
rect 291513 292961 291547 292989
rect 291575 292961 291609 292989
rect 291637 292961 291671 292989
rect 291699 292961 298728 292989
rect 298756 292961 298790 292989
rect 298818 292961 298852 292989
rect 298880 292961 298914 292989
rect 298942 292961 298990 292989
rect -958 292913 298990 292961
rect -958 290175 298990 290223
rect -958 290147 -430 290175
rect -402 290147 -368 290175
rect -340 290147 -306 290175
rect -278 290147 -244 290175
rect -216 290147 1625 290175
rect 1653 290147 1687 290175
rect 1715 290147 1749 290175
rect 1777 290147 1811 290175
rect 1839 290147 10625 290175
rect 10653 290147 10687 290175
rect 10715 290147 10749 290175
rect 10777 290147 10811 290175
rect 10839 290147 19625 290175
rect 19653 290147 19687 290175
rect 19715 290147 19749 290175
rect 19777 290147 19811 290175
rect 19839 290147 28625 290175
rect 28653 290147 28687 290175
rect 28715 290147 28749 290175
rect 28777 290147 28811 290175
rect 28839 290147 37625 290175
rect 37653 290147 37687 290175
rect 37715 290147 37749 290175
rect 37777 290147 37811 290175
rect 37839 290147 46625 290175
rect 46653 290147 46687 290175
rect 46715 290147 46749 290175
rect 46777 290147 46811 290175
rect 46839 290147 55625 290175
rect 55653 290147 55687 290175
rect 55715 290147 55749 290175
rect 55777 290147 55811 290175
rect 55839 290147 64625 290175
rect 64653 290147 64687 290175
rect 64715 290147 64749 290175
rect 64777 290147 64811 290175
rect 64839 290147 73625 290175
rect 73653 290147 73687 290175
rect 73715 290147 73749 290175
rect 73777 290147 73811 290175
rect 73839 290147 82625 290175
rect 82653 290147 82687 290175
rect 82715 290147 82749 290175
rect 82777 290147 82811 290175
rect 82839 290147 91625 290175
rect 91653 290147 91687 290175
rect 91715 290147 91749 290175
rect 91777 290147 91811 290175
rect 91839 290147 100625 290175
rect 100653 290147 100687 290175
rect 100715 290147 100749 290175
rect 100777 290147 100811 290175
rect 100839 290147 109625 290175
rect 109653 290147 109687 290175
rect 109715 290147 109749 290175
rect 109777 290147 109811 290175
rect 109839 290147 118625 290175
rect 118653 290147 118687 290175
rect 118715 290147 118749 290175
rect 118777 290147 118811 290175
rect 118839 290147 127625 290175
rect 127653 290147 127687 290175
rect 127715 290147 127749 290175
rect 127777 290147 127811 290175
rect 127839 290147 136625 290175
rect 136653 290147 136687 290175
rect 136715 290147 136749 290175
rect 136777 290147 136811 290175
rect 136839 290147 145625 290175
rect 145653 290147 145687 290175
rect 145715 290147 145749 290175
rect 145777 290147 145811 290175
rect 145839 290147 154625 290175
rect 154653 290147 154687 290175
rect 154715 290147 154749 290175
rect 154777 290147 154811 290175
rect 154839 290147 163625 290175
rect 163653 290147 163687 290175
rect 163715 290147 163749 290175
rect 163777 290147 163811 290175
rect 163839 290147 172625 290175
rect 172653 290147 172687 290175
rect 172715 290147 172749 290175
rect 172777 290147 172811 290175
rect 172839 290147 181625 290175
rect 181653 290147 181687 290175
rect 181715 290147 181749 290175
rect 181777 290147 181811 290175
rect 181839 290147 190625 290175
rect 190653 290147 190687 290175
rect 190715 290147 190749 290175
rect 190777 290147 190811 290175
rect 190839 290147 199625 290175
rect 199653 290147 199687 290175
rect 199715 290147 199749 290175
rect 199777 290147 199811 290175
rect 199839 290147 208625 290175
rect 208653 290147 208687 290175
rect 208715 290147 208749 290175
rect 208777 290147 208811 290175
rect 208839 290147 217625 290175
rect 217653 290147 217687 290175
rect 217715 290147 217749 290175
rect 217777 290147 217811 290175
rect 217839 290147 226625 290175
rect 226653 290147 226687 290175
rect 226715 290147 226749 290175
rect 226777 290147 226811 290175
rect 226839 290147 235625 290175
rect 235653 290147 235687 290175
rect 235715 290147 235749 290175
rect 235777 290147 235811 290175
rect 235839 290147 244625 290175
rect 244653 290147 244687 290175
rect 244715 290147 244749 290175
rect 244777 290147 244811 290175
rect 244839 290147 253625 290175
rect 253653 290147 253687 290175
rect 253715 290147 253749 290175
rect 253777 290147 253811 290175
rect 253839 290147 262625 290175
rect 262653 290147 262687 290175
rect 262715 290147 262749 290175
rect 262777 290147 262811 290175
rect 262839 290147 271625 290175
rect 271653 290147 271687 290175
rect 271715 290147 271749 290175
rect 271777 290147 271811 290175
rect 271839 290147 280625 290175
rect 280653 290147 280687 290175
rect 280715 290147 280749 290175
rect 280777 290147 280811 290175
rect 280839 290147 289625 290175
rect 289653 290147 289687 290175
rect 289715 290147 289749 290175
rect 289777 290147 289811 290175
rect 289839 290147 298248 290175
rect 298276 290147 298310 290175
rect 298338 290147 298372 290175
rect 298400 290147 298434 290175
rect 298462 290147 298990 290175
rect -958 290113 298990 290147
rect -958 290085 -430 290113
rect -402 290085 -368 290113
rect -340 290085 -306 290113
rect -278 290085 -244 290113
rect -216 290085 1625 290113
rect 1653 290085 1687 290113
rect 1715 290085 1749 290113
rect 1777 290085 1811 290113
rect 1839 290085 10625 290113
rect 10653 290085 10687 290113
rect 10715 290085 10749 290113
rect 10777 290085 10811 290113
rect 10839 290085 19625 290113
rect 19653 290085 19687 290113
rect 19715 290085 19749 290113
rect 19777 290085 19811 290113
rect 19839 290085 28625 290113
rect 28653 290085 28687 290113
rect 28715 290085 28749 290113
rect 28777 290085 28811 290113
rect 28839 290085 37625 290113
rect 37653 290085 37687 290113
rect 37715 290085 37749 290113
rect 37777 290085 37811 290113
rect 37839 290085 46625 290113
rect 46653 290085 46687 290113
rect 46715 290085 46749 290113
rect 46777 290085 46811 290113
rect 46839 290085 55625 290113
rect 55653 290085 55687 290113
rect 55715 290085 55749 290113
rect 55777 290085 55811 290113
rect 55839 290085 64625 290113
rect 64653 290085 64687 290113
rect 64715 290085 64749 290113
rect 64777 290085 64811 290113
rect 64839 290085 73625 290113
rect 73653 290085 73687 290113
rect 73715 290085 73749 290113
rect 73777 290085 73811 290113
rect 73839 290085 82625 290113
rect 82653 290085 82687 290113
rect 82715 290085 82749 290113
rect 82777 290085 82811 290113
rect 82839 290085 91625 290113
rect 91653 290085 91687 290113
rect 91715 290085 91749 290113
rect 91777 290085 91811 290113
rect 91839 290085 100625 290113
rect 100653 290085 100687 290113
rect 100715 290085 100749 290113
rect 100777 290085 100811 290113
rect 100839 290085 109625 290113
rect 109653 290085 109687 290113
rect 109715 290085 109749 290113
rect 109777 290085 109811 290113
rect 109839 290085 118625 290113
rect 118653 290085 118687 290113
rect 118715 290085 118749 290113
rect 118777 290085 118811 290113
rect 118839 290085 127625 290113
rect 127653 290085 127687 290113
rect 127715 290085 127749 290113
rect 127777 290085 127811 290113
rect 127839 290085 136625 290113
rect 136653 290085 136687 290113
rect 136715 290085 136749 290113
rect 136777 290085 136811 290113
rect 136839 290085 145625 290113
rect 145653 290085 145687 290113
rect 145715 290085 145749 290113
rect 145777 290085 145811 290113
rect 145839 290085 154625 290113
rect 154653 290085 154687 290113
rect 154715 290085 154749 290113
rect 154777 290085 154811 290113
rect 154839 290085 163625 290113
rect 163653 290085 163687 290113
rect 163715 290085 163749 290113
rect 163777 290085 163811 290113
rect 163839 290085 172625 290113
rect 172653 290085 172687 290113
rect 172715 290085 172749 290113
rect 172777 290085 172811 290113
rect 172839 290085 181625 290113
rect 181653 290085 181687 290113
rect 181715 290085 181749 290113
rect 181777 290085 181811 290113
rect 181839 290085 190625 290113
rect 190653 290085 190687 290113
rect 190715 290085 190749 290113
rect 190777 290085 190811 290113
rect 190839 290085 199625 290113
rect 199653 290085 199687 290113
rect 199715 290085 199749 290113
rect 199777 290085 199811 290113
rect 199839 290085 208625 290113
rect 208653 290085 208687 290113
rect 208715 290085 208749 290113
rect 208777 290085 208811 290113
rect 208839 290085 217625 290113
rect 217653 290085 217687 290113
rect 217715 290085 217749 290113
rect 217777 290085 217811 290113
rect 217839 290085 226625 290113
rect 226653 290085 226687 290113
rect 226715 290085 226749 290113
rect 226777 290085 226811 290113
rect 226839 290085 235625 290113
rect 235653 290085 235687 290113
rect 235715 290085 235749 290113
rect 235777 290085 235811 290113
rect 235839 290085 244625 290113
rect 244653 290085 244687 290113
rect 244715 290085 244749 290113
rect 244777 290085 244811 290113
rect 244839 290085 253625 290113
rect 253653 290085 253687 290113
rect 253715 290085 253749 290113
rect 253777 290085 253811 290113
rect 253839 290085 262625 290113
rect 262653 290085 262687 290113
rect 262715 290085 262749 290113
rect 262777 290085 262811 290113
rect 262839 290085 271625 290113
rect 271653 290085 271687 290113
rect 271715 290085 271749 290113
rect 271777 290085 271811 290113
rect 271839 290085 280625 290113
rect 280653 290085 280687 290113
rect 280715 290085 280749 290113
rect 280777 290085 280811 290113
rect 280839 290085 289625 290113
rect 289653 290085 289687 290113
rect 289715 290085 289749 290113
rect 289777 290085 289811 290113
rect 289839 290085 298248 290113
rect 298276 290085 298310 290113
rect 298338 290085 298372 290113
rect 298400 290085 298434 290113
rect 298462 290085 298990 290113
rect -958 290051 298990 290085
rect -958 290023 -430 290051
rect -402 290023 -368 290051
rect -340 290023 -306 290051
rect -278 290023 -244 290051
rect -216 290023 1625 290051
rect 1653 290023 1687 290051
rect 1715 290023 1749 290051
rect 1777 290023 1811 290051
rect 1839 290023 10625 290051
rect 10653 290023 10687 290051
rect 10715 290023 10749 290051
rect 10777 290023 10811 290051
rect 10839 290023 19625 290051
rect 19653 290023 19687 290051
rect 19715 290023 19749 290051
rect 19777 290023 19811 290051
rect 19839 290023 28625 290051
rect 28653 290023 28687 290051
rect 28715 290023 28749 290051
rect 28777 290023 28811 290051
rect 28839 290023 37625 290051
rect 37653 290023 37687 290051
rect 37715 290023 37749 290051
rect 37777 290023 37811 290051
rect 37839 290023 46625 290051
rect 46653 290023 46687 290051
rect 46715 290023 46749 290051
rect 46777 290023 46811 290051
rect 46839 290023 55625 290051
rect 55653 290023 55687 290051
rect 55715 290023 55749 290051
rect 55777 290023 55811 290051
rect 55839 290023 64625 290051
rect 64653 290023 64687 290051
rect 64715 290023 64749 290051
rect 64777 290023 64811 290051
rect 64839 290023 73625 290051
rect 73653 290023 73687 290051
rect 73715 290023 73749 290051
rect 73777 290023 73811 290051
rect 73839 290023 82625 290051
rect 82653 290023 82687 290051
rect 82715 290023 82749 290051
rect 82777 290023 82811 290051
rect 82839 290023 91625 290051
rect 91653 290023 91687 290051
rect 91715 290023 91749 290051
rect 91777 290023 91811 290051
rect 91839 290023 100625 290051
rect 100653 290023 100687 290051
rect 100715 290023 100749 290051
rect 100777 290023 100811 290051
rect 100839 290023 109625 290051
rect 109653 290023 109687 290051
rect 109715 290023 109749 290051
rect 109777 290023 109811 290051
rect 109839 290023 118625 290051
rect 118653 290023 118687 290051
rect 118715 290023 118749 290051
rect 118777 290023 118811 290051
rect 118839 290023 127625 290051
rect 127653 290023 127687 290051
rect 127715 290023 127749 290051
rect 127777 290023 127811 290051
rect 127839 290023 136625 290051
rect 136653 290023 136687 290051
rect 136715 290023 136749 290051
rect 136777 290023 136811 290051
rect 136839 290023 145625 290051
rect 145653 290023 145687 290051
rect 145715 290023 145749 290051
rect 145777 290023 145811 290051
rect 145839 290023 154625 290051
rect 154653 290023 154687 290051
rect 154715 290023 154749 290051
rect 154777 290023 154811 290051
rect 154839 290023 163625 290051
rect 163653 290023 163687 290051
rect 163715 290023 163749 290051
rect 163777 290023 163811 290051
rect 163839 290023 172625 290051
rect 172653 290023 172687 290051
rect 172715 290023 172749 290051
rect 172777 290023 172811 290051
rect 172839 290023 181625 290051
rect 181653 290023 181687 290051
rect 181715 290023 181749 290051
rect 181777 290023 181811 290051
rect 181839 290023 190625 290051
rect 190653 290023 190687 290051
rect 190715 290023 190749 290051
rect 190777 290023 190811 290051
rect 190839 290023 199625 290051
rect 199653 290023 199687 290051
rect 199715 290023 199749 290051
rect 199777 290023 199811 290051
rect 199839 290023 208625 290051
rect 208653 290023 208687 290051
rect 208715 290023 208749 290051
rect 208777 290023 208811 290051
rect 208839 290023 217625 290051
rect 217653 290023 217687 290051
rect 217715 290023 217749 290051
rect 217777 290023 217811 290051
rect 217839 290023 226625 290051
rect 226653 290023 226687 290051
rect 226715 290023 226749 290051
rect 226777 290023 226811 290051
rect 226839 290023 235625 290051
rect 235653 290023 235687 290051
rect 235715 290023 235749 290051
rect 235777 290023 235811 290051
rect 235839 290023 244625 290051
rect 244653 290023 244687 290051
rect 244715 290023 244749 290051
rect 244777 290023 244811 290051
rect 244839 290023 253625 290051
rect 253653 290023 253687 290051
rect 253715 290023 253749 290051
rect 253777 290023 253811 290051
rect 253839 290023 262625 290051
rect 262653 290023 262687 290051
rect 262715 290023 262749 290051
rect 262777 290023 262811 290051
rect 262839 290023 271625 290051
rect 271653 290023 271687 290051
rect 271715 290023 271749 290051
rect 271777 290023 271811 290051
rect 271839 290023 280625 290051
rect 280653 290023 280687 290051
rect 280715 290023 280749 290051
rect 280777 290023 280811 290051
rect 280839 290023 289625 290051
rect 289653 290023 289687 290051
rect 289715 290023 289749 290051
rect 289777 290023 289811 290051
rect 289839 290023 298248 290051
rect 298276 290023 298310 290051
rect 298338 290023 298372 290051
rect 298400 290023 298434 290051
rect 298462 290023 298990 290051
rect -958 289989 298990 290023
rect -958 289961 -430 289989
rect -402 289961 -368 289989
rect -340 289961 -306 289989
rect -278 289961 -244 289989
rect -216 289961 1625 289989
rect 1653 289961 1687 289989
rect 1715 289961 1749 289989
rect 1777 289961 1811 289989
rect 1839 289961 10625 289989
rect 10653 289961 10687 289989
rect 10715 289961 10749 289989
rect 10777 289961 10811 289989
rect 10839 289961 19625 289989
rect 19653 289961 19687 289989
rect 19715 289961 19749 289989
rect 19777 289961 19811 289989
rect 19839 289961 28625 289989
rect 28653 289961 28687 289989
rect 28715 289961 28749 289989
rect 28777 289961 28811 289989
rect 28839 289961 37625 289989
rect 37653 289961 37687 289989
rect 37715 289961 37749 289989
rect 37777 289961 37811 289989
rect 37839 289961 46625 289989
rect 46653 289961 46687 289989
rect 46715 289961 46749 289989
rect 46777 289961 46811 289989
rect 46839 289961 55625 289989
rect 55653 289961 55687 289989
rect 55715 289961 55749 289989
rect 55777 289961 55811 289989
rect 55839 289961 64625 289989
rect 64653 289961 64687 289989
rect 64715 289961 64749 289989
rect 64777 289961 64811 289989
rect 64839 289961 73625 289989
rect 73653 289961 73687 289989
rect 73715 289961 73749 289989
rect 73777 289961 73811 289989
rect 73839 289961 82625 289989
rect 82653 289961 82687 289989
rect 82715 289961 82749 289989
rect 82777 289961 82811 289989
rect 82839 289961 91625 289989
rect 91653 289961 91687 289989
rect 91715 289961 91749 289989
rect 91777 289961 91811 289989
rect 91839 289961 100625 289989
rect 100653 289961 100687 289989
rect 100715 289961 100749 289989
rect 100777 289961 100811 289989
rect 100839 289961 109625 289989
rect 109653 289961 109687 289989
rect 109715 289961 109749 289989
rect 109777 289961 109811 289989
rect 109839 289961 118625 289989
rect 118653 289961 118687 289989
rect 118715 289961 118749 289989
rect 118777 289961 118811 289989
rect 118839 289961 127625 289989
rect 127653 289961 127687 289989
rect 127715 289961 127749 289989
rect 127777 289961 127811 289989
rect 127839 289961 136625 289989
rect 136653 289961 136687 289989
rect 136715 289961 136749 289989
rect 136777 289961 136811 289989
rect 136839 289961 145625 289989
rect 145653 289961 145687 289989
rect 145715 289961 145749 289989
rect 145777 289961 145811 289989
rect 145839 289961 154625 289989
rect 154653 289961 154687 289989
rect 154715 289961 154749 289989
rect 154777 289961 154811 289989
rect 154839 289961 163625 289989
rect 163653 289961 163687 289989
rect 163715 289961 163749 289989
rect 163777 289961 163811 289989
rect 163839 289961 172625 289989
rect 172653 289961 172687 289989
rect 172715 289961 172749 289989
rect 172777 289961 172811 289989
rect 172839 289961 181625 289989
rect 181653 289961 181687 289989
rect 181715 289961 181749 289989
rect 181777 289961 181811 289989
rect 181839 289961 190625 289989
rect 190653 289961 190687 289989
rect 190715 289961 190749 289989
rect 190777 289961 190811 289989
rect 190839 289961 199625 289989
rect 199653 289961 199687 289989
rect 199715 289961 199749 289989
rect 199777 289961 199811 289989
rect 199839 289961 208625 289989
rect 208653 289961 208687 289989
rect 208715 289961 208749 289989
rect 208777 289961 208811 289989
rect 208839 289961 217625 289989
rect 217653 289961 217687 289989
rect 217715 289961 217749 289989
rect 217777 289961 217811 289989
rect 217839 289961 226625 289989
rect 226653 289961 226687 289989
rect 226715 289961 226749 289989
rect 226777 289961 226811 289989
rect 226839 289961 235625 289989
rect 235653 289961 235687 289989
rect 235715 289961 235749 289989
rect 235777 289961 235811 289989
rect 235839 289961 244625 289989
rect 244653 289961 244687 289989
rect 244715 289961 244749 289989
rect 244777 289961 244811 289989
rect 244839 289961 253625 289989
rect 253653 289961 253687 289989
rect 253715 289961 253749 289989
rect 253777 289961 253811 289989
rect 253839 289961 262625 289989
rect 262653 289961 262687 289989
rect 262715 289961 262749 289989
rect 262777 289961 262811 289989
rect 262839 289961 271625 289989
rect 271653 289961 271687 289989
rect 271715 289961 271749 289989
rect 271777 289961 271811 289989
rect 271839 289961 280625 289989
rect 280653 289961 280687 289989
rect 280715 289961 280749 289989
rect 280777 289961 280811 289989
rect 280839 289961 289625 289989
rect 289653 289961 289687 289989
rect 289715 289961 289749 289989
rect 289777 289961 289811 289989
rect 289839 289961 298248 289989
rect 298276 289961 298310 289989
rect 298338 289961 298372 289989
rect 298400 289961 298434 289989
rect 298462 289961 298990 289989
rect -958 289913 298990 289961
rect -958 284175 298990 284223
rect -958 284147 -910 284175
rect -882 284147 -848 284175
rect -820 284147 -786 284175
rect -758 284147 -724 284175
rect -696 284147 3485 284175
rect 3513 284147 3547 284175
rect 3575 284147 3609 284175
rect 3637 284147 3671 284175
rect 3699 284147 12485 284175
rect 12513 284147 12547 284175
rect 12575 284147 12609 284175
rect 12637 284147 12671 284175
rect 12699 284147 21485 284175
rect 21513 284147 21547 284175
rect 21575 284147 21609 284175
rect 21637 284147 21671 284175
rect 21699 284147 30485 284175
rect 30513 284147 30547 284175
rect 30575 284147 30609 284175
rect 30637 284147 30671 284175
rect 30699 284147 39485 284175
rect 39513 284147 39547 284175
rect 39575 284147 39609 284175
rect 39637 284147 39671 284175
rect 39699 284147 48485 284175
rect 48513 284147 48547 284175
rect 48575 284147 48609 284175
rect 48637 284147 48671 284175
rect 48699 284147 57485 284175
rect 57513 284147 57547 284175
rect 57575 284147 57609 284175
rect 57637 284147 57671 284175
rect 57699 284147 66485 284175
rect 66513 284147 66547 284175
rect 66575 284147 66609 284175
rect 66637 284147 66671 284175
rect 66699 284147 75485 284175
rect 75513 284147 75547 284175
rect 75575 284147 75609 284175
rect 75637 284147 75671 284175
rect 75699 284147 84485 284175
rect 84513 284147 84547 284175
rect 84575 284147 84609 284175
rect 84637 284147 84671 284175
rect 84699 284147 93485 284175
rect 93513 284147 93547 284175
rect 93575 284147 93609 284175
rect 93637 284147 93671 284175
rect 93699 284147 102485 284175
rect 102513 284147 102547 284175
rect 102575 284147 102609 284175
rect 102637 284147 102671 284175
rect 102699 284147 111485 284175
rect 111513 284147 111547 284175
rect 111575 284147 111609 284175
rect 111637 284147 111671 284175
rect 111699 284147 120485 284175
rect 120513 284147 120547 284175
rect 120575 284147 120609 284175
rect 120637 284147 120671 284175
rect 120699 284147 129485 284175
rect 129513 284147 129547 284175
rect 129575 284147 129609 284175
rect 129637 284147 129671 284175
rect 129699 284147 138485 284175
rect 138513 284147 138547 284175
rect 138575 284147 138609 284175
rect 138637 284147 138671 284175
rect 138699 284147 147485 284175
rect 147513 284147 147547 284175
rect 147575 284147 147609 284175
rect 147637 284147 147671 284175
rect 147699 284147 156485 284175
rect 156513 284147 156547 284175
rect 156575 284147 156609 284175
rect 156637 284147 156671 284175
rect 156699 284147 165485 284175
rect 165513 284147 165547 284175
rect 165575 284147 165609 284175
rect 165637 284147 165671 284175
rect 165699 284147 174485 284175
rect 174513 284147 174547 284175
rect 174575 284147 174609 284175
rect 174637 284147 174671 284175
rect 174699 284147 183485 284175
rect 183513 284147 183547 284175
rect 183575 284147 183609 284175
rect 183637 284147 183671 284175
rect 183699 284147 192485 284175
rect 192513 284147 192547 284175
rect 192575 284147 192609 284175
rect 192637 284147 192671 284175
rect 192699 284147 201485 284175
rect 201513 284147 201547 284175
rect 201575 284147 201609 284175
rect 201637 284147 201671 284175
rect 201699 284147 210485 284175
rect 210513 284147 210547 284175
rect 210575 284147 210609 284175
rect 210637 284147 210671 284175
rect 210699 284147 219485 284175
rect 219513 284147 219547 284175
rect 219575 284147 219609 284175
rect 219637 284147 219671 284175
rect 219699 284147 228485 284175
rect 228513 284147 228547 284175
rect 228575 284147 228609 284175
rect 228637 284147 228671 284175
rect 228699 284147 237485 284175
rect 237513 284147 237547 284175
rect 237575 284147 237609 284175
rect 237637 284147 237671 284175
rect 237699 284147 246485 284175
rect 246513 284147 246547 284175
rect 246575 284147 246609 284175
rect 246637 284147 246671 284175
rect 246699 284147 255485 284175
rect 255513 284147 255547 284175
rect 255575 284147 255609 284175
rect 255637 284147 255671 284175
rect 255699 284147 264485 284175
rect 264513 284147 264547 284175
rect 264575 284147 264609 284175
rect 264637 284147 264671 284175
rect 264699 284147 273485 284175
rect 273513 284147 273547 284175
rect 273575 284147 273609 284175
rect 273637 284147 273671 284175
rect 273699 284147 282485 284175
rect 282513 284147 282547 284175
rect 282575 284147 282609 284175
rect 282637 284147 282671 284175
rect 282699 284147 291485 284175
rect 291513 284147 291547 284175
rect 291575 284147 291609 284175
rect 291637 284147 291671 284175
rect 291699 284147 298728 284175
rect 298756 284147 298790 284175
rect 298818 284147 298852 284175
rect 298880 284147 298914 284175
rect 298942 284147 298990 284175
rect -958 284113 298990 284147
rect -958 284085 -910 284113
rect -882 284085 -848 284113
rect -820 284085 -786 284113
rect -758 284085 -724 284113
rect -696 284085 3485 284113
rect 3513 284085 3547 284113
rect 3575 284085 3609 284113
rect 3637 284085 3671 284113
rect 3699 284085 12485 284113
rect 12513 284085 12547 284113
rect 12575 284085 12609 284113
rect 12637 284085 12671 284113
rect 12699 284085 21485 284113
rect 21513 284085 21547 284113
rect 21575 284085 21609 284113
rect 21637 284085 21671 284113
rect 21699 284085 30485 284113
rect 30513 284085 30547 284113
rect 30575 284085 30609 284113
rect 30637 284085 30671 284113
rect 30699 284085 39485 284113
rect 39513 284085 39547 284113
rect 39575 284085 39609 284113
rect 39637 284085 39671 284113
rect 39699 284085 48485 284113
rect 48513 284085 48547 284113
rect 48575 284085 48609 284113
rect 48637 284085 48671 284113
rect 48699 284085 57485 284113
rect 57513 284085 57547 284113
rect 57575 284085 57609 284113
rect 57637 284085 57671 284113
rect 57699 284085 66485 284113
rect 66513 284085 66547 284113
rect 66575 284085 66609 284113
rect 66637 284085 66671 284113
rect 66699 284085 75485 284113
rect 75513 284085 75547 284113
rect 75575 284085 75609 284113
rect 75637 284085 75671 284113
rect 75699 284085 84485 284113
rect 84513 284085 84547 284113
rect 84575 284085 84609 284113
rect 84637 284085 84671 284113
rect 84699 284085 93485 284113
rect 93513 284085 93547 284113
rect 93575 284085 93609 284113
rect 93637 284085 93671 284113
rect 93699 284085 102485 284113
rect 102513 284085 102547 284113
rect 102575 284085 102609 284113
rect 102637 284085 102671 284113
rect 102699 284085 111485 284113
rect 111513 284085 111547 284113
rect 111575 284085 111609 284113
rect 111637 284085 111671 284113
rect 111699 284085 120485 284113
rect 120513 284085 120547 284113
rect 120575 284085 120609 284113
rect 120637 284085 120671 284113
rect 120699 284085 129485 284113
rect 129513 284085 129547 284113
rect 129575 284085 129609 284113
rect 129637 284085 129671 284113
rect 129699 284085 138485 284113
rect 138513 284085 138547 284113
rect 138575 284085 138609 284113
rect 138637 284085 138671 284113
rect 138699 284085 147485 284113
rect 147513 284085 147547 284113
rect 147575 284085 147609 284113
rect 147637 284085 147671 284113
rect 147699 284085 156485 284113
rect 156513 284085 156547 284113
rect 156575 284085 156609 284113
rect 156637 284085 156671 284113
rect 156699 284085 165485 284113
rect 165513 284085 165547 284113
rect 165575 284085 165609 284113
rect 165637 284085 165671 284113
rect 165699 284085 174485 284113
rect 174513 284085 174547 284113
rect 174575 284085 174609 284113
rect 174637 284085 174671 284113
rect 174699 284085 183485 284113
rect 183513 284085 183547 284113
rect 183575 284085 183609 284113
rect 183637 284085 183671 284113
rect 183699 284085 192485 284113
rect 192513 284085 192547 284113
rect 192575 284085 192609 284113
rect 192637 284085 192671 284113
rect 192699 284085 201485 284113
rect 201513 284085 201547 284113
rect 201575 284085 201609 284113
rect 201637 284085 201671 284113
rect 201699 284085 210485 284113
rect 210513 284085 210547 284113
rect 210575 284085 210609 284113
rect 210637 284085 210671 284113
rect 210699 284085 219485 284113
rect 219513 284085 219547 284113
rect 219575 284085 219609 284113
rect 219637 284085 219671 284113
rect 219699 284085 228485 284113
rect 228513 284085 228547 284113
rect 228575 284085 228609 284113
rect 228637 284085 228671 284113
rect 228699 284085 237485 284113
rect 237513 284085 237547 284113
rect 237575 284085 237609 284113
rect 237637 284085 237671 284113
rect 237699 284085 246485 284113
rect 246513 284085 246547 284113
rect 246575 284085 246609 284113
rect 246637 284085 246671 284113
rect 246699 284085 255485 284113
rect 255513 284085 255547 284113
rect 255575 284085 255609 284113
rect 255637 284085 255671 284113
rect 255699 284085 264485 284113
rect 264513 284085 264547 284113
rect 264575 284085 264609 284113
rect 264637 284085 264671 284113
rect 264699 284085 273485 284113
rect 273513 284085 273547 284113
rect 273575 284085 273609 284113
rect 273637 284085 273671 284113
rect 273699 284085 282485 284113
rect 282513 284085 282547 284113
rect 282575 284085 282609 284113
rect 282637 284085 282671 284113
rect 282699 284085 291485 284113
rect 291513 284085 291547 284113
rect 291575 284085 291609 284113
rect 291637 284085 291671 284113
rect 291699 284085 298728 284113
rect 298756 284085 298790 284113
rect 298818 284085 298852 284113
rect 298880 284085 298914 284113
rect 298942 284085 298990 284113
rect -958 284051 298990 284085
rect -958 284023 -910 284051
rect -882 284023 -848 284051
rect -820 284023 -786 284051
rect -758 284023 -724 284051
rect -696 284023 3485 284051
rect 3513 284023 3547 284051
rect 3575 284023 3609 284051
rect 3637 284023 3671 284051
rect 3699 284023 12485 284051
rect 12513 284023 12547 284051
rect 12575 284023 12609 284051
rect 12637 284023 12671 284051
rect 12699 284023 21485 284051
rect 21513 284023 21547 284051
rect 21575 284023 21609 284051
rect 21637 284023 21671 284051
rect 21699 284023 30485 284051
rect 30513 284023 30547 284051
rect 30575 284023 30609 284051
rect 30637 284023 30671 284051
rect 30699 284023 39485 284051
rect 39513 284023 39547 284051
rect 39575 284023 39609 284051
rect 39637 284023 39671 284051
rect 39699 284023 48485 284051
rect 48513 284023 48547 284051
rect 48575 284023 48609 284051
rect 48637 284023 48671 284051
rect 48699 284023 57485 284051
rect 57513 284023 57547 284051
rect 57575 284023 57609 284051
rect 57637 284023 57671 284051
rect 57699 284023 66485 284051
rect 66513 284023 66547 284051
rect 66575 284023 66609 284051
rect 66637 284023 66671 284051
rect 66699 284023 75485 284051
rect 75513 284023 75547 284051
rect 75575 284023 75609 284051
rect 75637 284023 75671 284051
rect 75699 284023 84485 284051
rect 84513 284023 84547 284051
rect 84575 284023 84609 284051
rect 84637 284023 84671 284051
rect 84699 284023 93485 284051
rect 93513 284023 93547 284051
rect 93575 284023 93609 284051
rect 93637 284023 93671 284051
rect 93699 284023 102485 284051
rect 102513 284023 102547 284051
rect 102575 284023 102609 284051
rect 102637 284023 102671 284051
rect 102699 284023 111485 284051
rect 111513 284023 111547 284051
rect 111575 284023 111609 284051
rect 111637 284023 111671 284051
rect 111699 284023 120485 284051
rect 120513 284023 120547 284051
rect 120575 284023 120609 284051
rect 120637 284023 120671 284051
rect 120699 284023 129485 284051
rect 129513 284023 129547 284051
rect 129575 284023 129609 284051
rect 129637 284023 129671 284051
rect 129699 284023 138485 284051
rect 138513 284023 138547 284051
rect 138575 284023 138609 284051
rect 138637 284023 138671 284051
rect 138699 284023 147485 284051
rect 147513 284023 147547 284051
rect 147575 284023 147609 284051
rect 147637 284023 147671 284051
rect 147699 284023 156485 284051
rect 156513 284023 156547 284051
rect 156575 284023 156609 284051
rect 156637 284023 156671 284051
rect 156699 284023 165485 284051
rect 165513 284023 165547 284051
rect 165575 284023 165609 284051
rect 165637 284023 165671 284051
rect 165699 284023 174485 284051
rect 174513 284023 174547 284051
rect 174575 284023 174609 284051
rect 174637 284023 174671 284051
rect 174699 284023 183485 284051
rect 183513 284023 183547 284051
rect 183575 284023 183609 284051
rect 183637 284023 183671 284051
rect 183699 284023 192485 284051
rect 192513 284023 192547 284051
rect 192575 284023 192609 284051
rect 192637 284023 192671 284051
rect 192699 284023 201485 284051
rect 201513 284023 201547 284051
rect 201575 284023 201609 284051
rect 201637 284023 201671 284051
rect 201699 284023 210485 284051
rect 210513 284023 210547 284051
rect 210575 284023 210609 284051
rect 210637 284023 210671 284051
rect 210699 284023 219485 284051
rect 219513 284023 219547 284051
rect 219575 284023 219609 284051
rect 219637 284023 219671 284051
rect 219699 284023 228485 284051
rect 228513 284023 228547 284051
rect 228575 284023 228609 284051
rect 228637 284023 228671 284051
rect 228699 284023 237485 284051
rect 237513 284023 237547 284051
rect 237575 284023 237609 284051
rect 237637 284023 237671 284051
rect 237699 284023 246485 284051
rect 246513 284023 246547 284051
rect 246575 284023 246609 284051
rect 246637 284023 246671 284051
rect 246699 284023 255485 284051
rect 255513 284023 255547 284051
rect 255575 284023 255609 284051
rect 255637 284023 255671 284051
rect 255699 284023 264485 284051
rect 264513 284023 264547 284051
rect 264575 284023 264609 284051
rect 264637 284023 264671 284051
rect 264699 284023 273485 284051
rect 273513 284023 273547 284051
rect 273575 284023 273609 284051
rect 273637 284023 273671 284051
rect 273699 284023 282485 284051
rect 282513 284023 282547 284051
rect 282575 284023 282609 284051
rect 282637 284023 282671 284051
rect 282699 284023 291485 284051
rect 291513 284023 291547 284051
rect 291575 284023 291609 284051
rect 291637 284023 291671 284051
rect 291699 284023 298728 284051
rect 298756 284023 298790 284051
rect 298818 284023 298852 284051
rect 298880 284023 298914 284051
rect 298942 284023 298990 284051
rect -958 283989 298990 284023
rect -958 283961 -910 283989
rect -882 283961 -848 283989
rect -820 283961 -786 283989
rect -758 283961 -724 283989
rect -696 283961 3485 283989
rect 3513 283961 3547 283989
rect 3575 283961 3609 283989
rect 3637 283961 3671 283989
rect 3699 283961 12485 283989
rect 12513 283961 12547 283989
rect 12575 283961 12609 283989
rect 12637 283961 12671 283989
rect 12699 283961 21485 283989
rect 21513 283961 21547 283989
rect 21575 283961 21609 283989
rect 21637 283961 21671 283989
rect 21699 283961 30485 283989
rect 30513 283961 30547 283989
rect 30575 283961 30609 283989
rect 30637 283961 30671 283989
rect 30699 283961 39485 283989
rect 39513 283961 39547 283989
rect 39575 283961 39609 283989
rect 39637 283961 39671 283989
rect 39699 283961 48485 283989
rect 48513 283961 48547 283989
rect 48575 283961 48609 283989
rect 48637 283961 48671 283989
rect 48699 283961 57485 283989
rect 57513 283961 57547 283989
rect 57575 283961 57609 283989
rect 57637 283961 57671 283989
rect 57699 283961 66485 283989
rect 66513 283961 66547 283989
rect 66575 283961 66609 283989
rect 66637 283961 66671 283989
rect 66699 283961 75485 283989
rect 75513 283961 75547 283989
rect 75575 283961 75609 283989
rect 75637 283961 75671 283989
rect 75699 283961 84485 283989
rect 84513 283961 84547 283989
rect 84575 283961 84609 283989
rect 84637 283961 84671 283989
rect 84699 283961 93485 283989
rect 93513 283961 93547 283989
rect 93575 283961 93609 283989
rect 93637 283961 93671 283989
rect 93699 283961 102485 283989
rect 102513 283961 102547 283989
rect 102575 283961 102609 283989
rect 102637 283961 102671 283989
rect 102699 283961 111485 283989
rect 111513 283961 111547 283989
rect 111575 283961 111609 283989
rect 111637 283961 111671 283989
rect 111699 283961 120485 283989
rect 120513 283961 120547 283989
rect 120575 283961 120609 283989
rect 120637 283961 120671 283989
rect 120699 283961 129485 283989
rect 129513 283961 129547 283989
rect 129575 283961 129609 283989
rect 129637 283961 129671 283989
rect 129699 283961 138485 283989
rect 138513 283961 138547 283989
rect 138575 283961 138609 283989
rect 138637 283961 138671 283989
rect 138699 283961 147485 283989
rect 147513 283961 147547 283989
rect 147575 283961 147609 283989
rect 147637 283961 147671 283989
rect 147699 283961 156485 283989
rect 156513 283961 156547 283989
rect 156575 283961 156609 283989
rect 156637 283961 156671 283989
rect 156699 283961 165485 283989
rect 165513 283961 165547 283989
rect 165575 283961 165609 283989
rect 165637 283961 165671 283989
rect 165699 283961 174485 283989
rect 174513 283961 174547 283989
rect 174575 283961 174609 283989
rect 174637 283961 174671 283989
rect 174699 283961 183485 283989
rect 183513 283961 183547 283989
rect 183575 283961 183609 283989
rect 183637 283961 183671 283989
rect 183699 283961 192485 283989
rect 192513 283961 192547 283989
rect 192575 283961 192609 283989
rect 192637 283961 192671 283989
rect 192699 283961 201485 283989
rect 201513 283961 201547 283989
rect 201575 283961 201609 283989
rect 201637 283961 201671 283989
rect 201699 283961 210485 283989
rect 210513 283961 210547 283989
rect 210575 283961 210609 283989
rect 210637 283961 210671 283989
rect 210699 283961 219485 283989
rect 219513 283961 219547 283989
rect 219575 283961 219609 283989
rect 219637 283961 219671 283989
rect 219699 283961 228485 283989
rect 228513 283961 228547 283989
rect 228575 283961 228609 283989
rect 228637 283961 228671 283989
rect 228699 283961 237485 283989
rect 237513 283961 237547 283989
rect 237575 283961 237609 283989
rect 237637 283961 237671 283989
rect 237699 283961 246485 283989
rect 246513 283961 246547 283989
rect 246575 283961 246609 283989
rect 246637 283961 246671 283989
rect 246699 283961 255485 283989
rect 255513 283961 255547 283989
rect 255575 283961 255609 283989
rect 255637 283961 255671 283989
rect 255699 283961 264485 283989
rect 264513 283961 264547 283989
rect 264575 283961 264609 283989
rect 264637 283961 264671 283989
rect 264699 283961 273485 283989
rect 273513 283961 273547 283989
rect 273575 283961 273609 283989
rect 273637 283961 273671 283989
rect 273699 283961 282485 283989
rect 282513 283961 282547 283989
rect 282575 283961 282609 283989
rect 282637 283961 282671 283989
rect 282699 283961 291485 283989
rect 291513 283961 291547 283989
rect 291575 283961 291609 283989
rect 291637 283961 291671 283989
rect 291699 283961 298728 283989
rect 298756 283961 298790 283989
rect 298818 283961 298852 283989
rect 298880 283961 298914 283989
rect 298942 283961 298990 283989
rect -958 283913 298990 283961
rect -958 281175 298990 281223
rect -958 281147 -430 281175
rect -402 281147 -368 281175
rect -340 281147 -306 281175
rect -278 281147 -244 281175
rect -216 281147 1625 281175
rect 1653 281147 1687 281175
rect 1715 281147 1749 281175
rect 1777 281147 1811 281175
rect 1839 281147 10625 281175
rect 10653 281147 10687 281175
rect 10715 281147 10749 281175
rect 10777 281147 10811 281175
rect 10839 281147 19625 281175
rect 19653 281147 19687 281175
rect 19715 281147 19749 281175
rect 19777 281147 19811 281175
rect 19839 281147 28625 281175
rect 28653 281147 28687 281175
rect 28715 281147 28749 281175
rect 28777 281147 28811 281175
rect 28839 281147 37625 281175
rect 37653 281147 37687 281175
rect 37715 281147 37749 281175
rect 37777 281147 37811 281175
rect 37839 281147 46625 281175
rect 46653 281147 46687 281175
rect 46715 281147 46749 281175
rect 46777 281147 46811 281175
rect 46839 281147 55625 281175
rect 55653 281147 55687 281175
rect 55715 281147 55749 281175
rect 55777 281147 55811 281175
rect 55839 281147 64625 281175
rect 64653 281147 64687 281175
rect 64715 281147 64749 281175
rect 64777 281147 64811 281175
rect 64839 281147 73625 281175
rect 73653 281147 73687 281175
rect 73715 281147 73749 281175
rect 73777 281147 73811 281175
rect 73839 281147 82625 281175
rect 82653 281147 82687 281175
rect 82715 281147 82749 281175
rect 82777 281147 82811 281175
rect 82839 281147 91625 281175
rect 91653 281147 91687 281175
rect 91715 281147 91749 281175
rect 91777 281147 91811 281175
rect 91839 281147 100625 281175
rect 100653 281147 100687 281175
rect 100715 281147 100749 281175
rect 100777 281147 100811 281175
rect 100839 281147 109625 281175
rect 109653 281147 109687 281175
rect 109715 281147 109749 281175
rect 109777 281147 109811 281175
rect 109839 281147 118625 281175
rect 118653 281147 118687 281175
rect 118715 281147 118749 281175
rect 118777 281147 118811 281175
rect 118839 281147 127625 281175
rect 127653 281147 127687 281175
rect 127715 281147 127749 281175
rect 127777 281147 127811 281175
rect 127839 281147 136625 281175
rect 136653 281147 136687 281175
rect 136715 281147 136749 281175
rect 136777 281147 136811 281175
rect 136839 281147 145625 281175
rect 145653 281147 145687 281175
rect 145715 281147 145749 281175
rect 145777 281147 145811 281175
rect 145839 281147 154625 281175
rect 154653 281147 154687 281175
rect 154715 281147 154749 281175
rect 154777 281147 154811 281175
rect 154839 281147 163625 281175
rect 163653 281147 163687 281175
rect 163715 281147 163749 281175
rect 163777 281147 163811 281175
rect 163839 281147 172625 281175
rect 172653 281147 172687 281175
rect 172715 281147 172749 281175
rect 172777 281147 172811 281175
rect 172839 281147 181625 281175
rect 181653 281147 181687 281175
rect 181715 281147 181749 281175
rect 181777 281147 181811 281175
rect 181839 281147 190625 281175
rect 190653 281147 190687 281175
rect 190715 281147 190749 281175
rect 190777 281147 190811 281175
rect 190839 281147 199625 281175
rect 199653 281147 199687 281175
rect 199715 281147 199749 281175
rect 199777 281147 199811 281175
rect 199839 281147 208625 281175
rect 208653 281147 208687 281175
rect 208715 281147 208749 281175
rect 208777 281147 208811 281175
rect 208839 281147 217625 281175
rect 217653 281147 217687 281175
rect 217715 281147 217749 281175
rect 217777 281147 217811 281175
rect 217839 281147 226625 281175
rect 226653 281147 226687 281175
rect 226715 281147 226749 281175
rect 226777 281147 226811 281175
rect 226839 281147 235625 281175
rect 235653 281147 235687 281175
rect 235715 281147 235749 281175
rect 235777 281147 235811 281175
rect 235839 281147 244625 281175
rect 244653 281147 244687 281175
rect 244715 281147 244749 281175
rect 244777 281147 244811 281175
rect 244839 281147 253625 281175
rect 253653 281147 253687 281175
rect 253715 281147 253749 281175
rect 253777 281147 253811 281175
rect 253839 281147 262625 281175
rect 262653 281147 262687 281175
rect 262715 281147 262749 281175
rect 262777 281147 262811 281175
rect 262839 281147 271625 281175
rect 271653 281147 271687 281175
rect 271715 281147 271749 281175
rect 271777 281147 271811 281175
rect 271839 281147 280625 281175
rect 280653 281147 280687 281175
rect 280715 281147 280749 281175
rect 280777 281147 280811 281175
rect 280839 281147 289625 281175
rect 289653 281147 289687 281175
rect 289715 281147 289749 281175
rect 289777 281147 289811 281175
rect 289839 281147 298248 281175
rect 298276 281147 298310 281175
rect 298338 281147 298372 281175
rect 298400 281147 298434 281175
rect 298462 281147 298990 281175
rect -958 281113 298990 281147
rect -958 281085 -430 281113
rect -402 281085 -368 281113
rect -340 281085 -306 281113
rect -278 281085 -244 281113
rect -216 281085 1625 281113
rect 1653 281085 1687 281113
rect 1715 281085 1749 281113
rect 1777 281085 1811 281113
rect 1839 281085 10625 281113
rect 10653 281085 10687 281113
rect 10715 281085 10749 281113
rect 10777 281085 10811 281113
rect 10839 281085 19625 281113
rect 19653 281085 19687 281113
rect 19715 281085 19749 281113
rect 19777 281085 19811 281113
rect 19839 281085 28625 281113
rect 28653 281085 28687 281113
rect 28715 281085 28749 281113
rect 28777 281085 28811 281113
rect 28839 281085 37625 281113
rect 37653 281085 37687 281113
rect 37715 281085 37749 281113
rect 37777 281085 37811 281113
rect 37839 281085 46625 281113
rect 46653 281085 46687 281113
rect 46715 281085 46749 281113
rect 46777 281085 46811 281113
rect 46839 281085 55625 281113
rect 55653 281085 55687 281113
rect 55715 281085 55749 281113
rect 55777 281085 55811 281113
rect 55839 281085 64625 281113
rect 64653 281085 64687 281113
rect 64715 281085 64749 281113
rect 64777 281085 64811 281113
rect 64839 281085 73625 281113
rect 73653 281085 73687 281113
rect 73715 281085 73749 281113
rect 73777 281085 73811 281113
rect 73839 281085 82625 281113
rect 82653 281085 82687 281113
rect 82715 281085 82749 281113
rect 82777 281085 82811 281113
rect 82839 281085 91625 281113
rect 91653 281085 91687 281113
rect 91715 281085 91749 281113
rect 91777 281085 91811 281113
rect 91839 281085 100625 281113
rect 100653 281085 100687 281113
rect 100715 281085 100749 281113
rect 100777 281085 100811 281113
rect 100839 281085 109625 281113
rect 109653 281085 109687 281113
rect 109715 281085 109749 281113
rect 109777 281085 109811 281113
rect 109839 281085 118625 281113
rect 118653 281085 118687 281113
rect 118715 281085 118749 281113
rect 118777 281085 118811 281113
rect 118839 281085 127625 281113
rect 127653 281085 127687 281113
rect 127715 281085 127749 281113
rect 127777 281085 127811 281113
rect 127839 281085 136625 281113
rect 136653 281085 136687 281113
rect 136715 281085 136749 281113
rect 136777 281085 136811 281113
rect 136839 281085 145625 281113
rect 145653 281085 145687 281113
rect 145715 281085 145749 281113
rect 145777 281085 145811 281113
rect 145839 281085 154625 281113
rect 154653 281085 154687 281113
rect 154715 281085 154749 281113
rect 154777 281085 154811 281113
rect 154839 281085 163625 281113
rect 163653 281085 163687 281113
rect 163715 281085 163749 281113
rect 163777 281085 163811 281113
rect 163839 281085 172625 281113
rect 172653 281085 172687 281113
rect 172715 281085 172749 281113
rect 172777 281085 172811 281113
rect 172839 281085 181625 281113
rect 181653 281085 181687 281113
rect 181715 281085 181749 281113
rect 181777 281085 181811 281113
rect 181839 281085 190625 281113
rect 190653 281085 190687 281113
rect 190715 281085 190749 281113
rect 190777 281085 190811 281113
rect 190839 281085 199625 281113
rect 199653 281085 199687 281113
rect 199715 281085 199749 281113
rect 199777 281085 199811 281113
rect 199839 281085 208625 281113
rect 208653 281085 208687 281113
rect 208715 281085 208749 281113
rect 208777 281085 208811 281113
rect 208839 281085 217625 281113
rect 217653 281085 217687 281113
rect 217715 281085 217749 281113
rect 217777 281085 217811 281113
rect 217839 281085 226625 281113
rect 226653 281085 226687 281113
rect 226715 281085 226749 281113
rect 226777 281085 226811 281113
rect 226839 281085 235625 281113
rect 235653 281085 235687 281113
rect 235715 281085 235749 281113
rect 235777 281085 235811 281113
rect 235839 281085 244625 281113
rect 244653 281085 244687 281113
rect 244715 281085 244749 281113
rect 244777 281085 244811 281113
rect 244839 281085 253625 281113
rect 253653 281085 253687 281113
rect 253715 281085 253749 281113
rect 253777 281085 253811 281113
rect 253839 281085 262625 281113
rect 262653 281085 262687 281113
rect 262715 281085 262749 281113
rect 262777 281085 262811 281113
rect 262839 281085 271625 281113
rect 271653 281085 271687 281113
rect 271715 281085 271749 281113
rect 271777 281085 271811 281113
rect 271839 281085 280625 281113
rect 280653 281085 280687 281113
rect 280715 281085 280749 281113
rect 280777 281085 280811 281113
rect 280839 281085 289625 281113
rect 289653 281085 289687 281113
rect 289715 281085 289749 281113
rect 289777 281085 289811 281113
rect 289839 281085 298248 281113
rect 298276 281085 298310 281113
rect 298338 281085 298372 281113
rect 298400 281085 298434 281113
rect 298462 281085 298990 281113
rect -958 281051 298990 281085
rect -958 281023 -430 281051
rect -402 281023 -368 281051
rect -340 281023 -306 281051
rect -278 281023 -244 281051
rect -216 281023 1625 281051
rect 1653 281023 1687 281051
rect 1715 281023 1749 281051
rect 1777 281023 1811 281051
rect 1839 281023 10625 281051
rect 10653 281023 10687 281051
rect 10715 281023 10749 281051
rect 10777 281023 10811 281051
rect 10839 281023 19625 281051
rect 19653 281023 19687 281051
rect 19715 281023 19749 281051
rect 19777 281023 19811 281051
rect 19839 281023 28625 281051
rect 28653 281023 28687 281051
rect 28715 281023 28749 281051
rect 28777 281023 28811 281051
rect 28839 281023 37625 281051
rect 37653 281023 37687 281051
rect 37715 281023 37749 281051
rect 37777 281023 37811 281051
rect 37839 281023 46625 281051
rect 46653 281023 46687 281051
rect 46715 281023 46749 281051
rect 46777 281023 46811 281051
rect 46839 281023 55625 281051
rect 55653 281023 55687 281051
rect 55715 281023 55749 281051
rect 55777 281023 55811 281051
rect 55839 281023 64625 281051
rect 64653 281023 64687 281051
rect 64715 281023 64749 281051
rect 64777 281023 64811 281051
rect 64839 281023 73625 281051
rect 73653 281023 73687 281051
rect 73715 281023 73749 281051
rect 73777 281023 73811 281051
rect 73839 281023 82625 281051
rect 82653 281023 82687 281051
rect 82715 281023 82749 281051
rect 82777 281023 82811 281051
rect 82839 281023 91625 281051
rect 91653 281023 91687 281051
rect 91715 281023 91749 281051
rect 91777 281023 91811 281051
rect 91839 281023 100625 281051
rect 100653 281023 100687 281051
rect 100715 281023 100749 281051
rect 100777 281023 100811 281051
rect 100839 281023 109625 281051
rect 109653 281023 109687 281051
rect 109715 281023 109749 281051
rect 109777 281023 109811 281051
rect 109839 281023 118625 281051
rect 118653 281023 118687 281051
rect 118715 281023 118749 281051
rect 118777 281023 118811 281051
rect 118839 281023 127625 281051
rect 127653 281023 127687 281051
rect 127715 281023 127749 281051
rect 127777 281023 127811 281051
rect 127839 281023 136625 281051
rect 136653 281023 136687 281051
rect 136715 281023 136749 281051
rect 136777 281023 136811 281051
rect 136839 281023 145625 281051
rect 145653 281023 145687 281051
rect 145715 281023 145749 281051
rect 145777 281023 145811 281051
rect 145839 281023 154625 281051
rect 154653 281023 154687 281051
rect 154715 281023 154749 281051
rect 154777 281023 154811 281051
rect 154839 281023 163625 281051
rect 163653 281023 163687 281051
rect 163715 281023 163749 281051
rect 163777 281023 163811 281051
rect 163839 281023 172625 281051
rect 172653 281023 172687 281051
rect 172715 281023 172749 281051
rect 172777 281023 172811 281051
rect 172839 281023 181625 281051
rect 181653 281023 181687 281051
rect 181715 281023 181749 281051
rect 181777 281023 181811 281051
rect 181839 281023 190625 281051
rect 190653 281023 190687 281051
rect 190715 281023 190749 281051
rect 190777 281023 190811 281051
rect 190839 281023 199625 281051
rect 199653 281023 199687 281051
rect 199715 281023 199749 281051
rect 199777 281023 199811 281051
rect 199839 281023 208625 281051
rect 208653 281023 208687 281051
rect 208715 281023 208749 281051
rect 208777 281023 208811 281051
rect 208839 281023 217625 281051
rect 217653 281023 217687 281051
rect 217715 281023 217749 281051
rect 217777 281023 217811 281051
rect 217839 281023 226625 281051
rect 226653 281023 226687 281051
rect 226715 281023 226749 281051
rect 226777 281023 226811 281051
rect 226839 281023 235625 281051
rect 235653 281023 235687 281051
rect 235715 281023 235749 281051
rect 235777 281023 235811 281051
rect 235839 281023 244625 281051
rect 244653 281023 244687 281051
rect 244715 281023 244749 281051
rect 244777 281023 244811 281051
rect 244839 281023 253625 281051
rect 253653 281023 253687 281051
rect 253715 281023 253749 281051
rect 253777 281023 253811 281051
rect 253839 281023 262625 281051
rect 262653 281023 262687 281051
rect 262715 281023 262749 281051
rect 262777 281023 262811 281051
rect 262839 281023 271625 281051
rect 271653 281023 271687 281051
rect 271715 281023 271749 281051
rect 271777 281023 271811 281051
rect 271839 281023 280625 281051
rect 280653 281023 280687 281051
rect 280715 281023 280749 281051
rect 280777 281023 280811 281051
rect 280839 281023 289625 281051
rect 289653 281023 289687 281051
rect 289715 281023 289749 281051
rect 289777 281023 289811 281051
rect 289839 281023 298248 281051
rect 298276 281023 298310 281051
rect 298338 281023 298372 281051
rect 298400 281023 298434 281051
rect 298462 281023 298990 281051
rect -958 280989 298990 281023
rect -958 280961 -430 280989
rect -402 280961 -368 280989
rect -340 280961 -306 280989
rect -278 280961 -244 280989
rect -216 280961 1625 280989
rect 1653 280961 1687 280989
rect 1715 280961 1749 280989
rect 1777 280961 1811 280989
rect 1839 280961 10625 280989
rect 10653 280961 10687 280989
rect 10715 280961 10749 280989
rect 10777 280961 10811 280989
rect 10839 280961 19625 280989
rect 19653 280961 19687 280989
rect 19715 280961 19749 280989
rect 19777 280961 19811 280989
rect 19839 280961 28625 280989
rect 28653 280961 28687 280989
rect 28715 280961 28749 280989
rect 28777 280961 28811 280989
rect 28839 280961 37625 280989
rect 37653 280961 37687 280989
rect 37715 280961 37749 280989
rect 37777 280961 37811 280989
rect 37839 280961 46625 280989
rect 46653 280961 46687 280989
rect 46715 280961 46749 280989
rect 46777 280961 46811 280989
rect 46839 280961 55625 280989
rect 55653 280961 55687 280989
rect 55715 280961 55749 280989
rect 55777 280961 55811 280989
rect 55839 280961 64625 280989
rect 64653 280961 64687 280989
rect 64715 280961 64749 280989
rect 64777 280961 64811 280989
rect 64839 280961 73625 280989
rect 73653 280961 73687 280989
rect 73715 280961 73749 280989
rect 73777 280961 73811 280989
rect 73839 280961 82625 280989
rect 82653 280961 82687 280989
rect 82715 280961 82749 280989
rect 82777 280961 82811 280989
rect 82839 280961 91625 280989
rect 91653 280961 91687 280989
rect 91715 280961 91749 280989
rect 91777 280961 91811 280989
rect 91839 280961 100625 280989
rect 100653 280961 100687 280989
rect 100715 280961 100749 280989
rect 100777 280961 100811 280989
rect 100839 280961 109625 280989
rect 109653 280961 109687 280989
rect 109715 280961 109749 280989
rect 109777 280961 109811 280989
rect 109839 280961 118625 280989
rect 118653 280961 118687 280989
rect 118715 280961 118749 280989
rect 118777 280961 118811 280989
rect 118839 280961 127625 280989
rect 127653 280961 127687 280989
rect 127715 280961 127749 280989
rect 127777 280961 127811 280989
rect 127839 280961 136625 280989
rect 136653 280961 136687 280989
rect 136715 280961 136749 280989
rect 136777 280961 136811 280989
rect 136839 280961 145625 280989
rect 145653 280961 145687 280989
rect 145715 280961 145749 280989
rect 145777 280961 145811 280989
rect 145839 280961 154625 280989
rect 154653 280961 154687 280989
rect 154715 280961 154749 280989
rect 154777 280961 154811 280989
rect 154839 280961 163625 280989
rect 163653 280961 163687 280989
rect 163715 280961 163749 280989
rect 163777 280961 163811 280989
rect 163839 280961 172625 280989
rect 172653 280961 172687 280989
rect 172715 280961 172749 280989
rect 172777 280961 172811 280989
rect 172839 280961 181625 280989
rect 181653 280961 181687 280989
rect 181715 280961 181749 280989
rect 181777 280961 181811 280989
rect 181839 280961 190625 280989
rect 190653 280961 190687 280989
rect 190715 280961 190749 280989
rect 190777 280961 190811 280989
rect 190839 280961 199625 280989
rect 199653 280961 199687 280989
rect 199715 280961 199749 280989
rect 199777 280961 199811 280989
rect 199839 280961 208625 280989
rect 208653 280961 208687 280989
rect 208715 280961 208749 280989
rect 208777 280961 208811 280989
rect 208839 280961 217625 280989
rect 217653 280961 217687 280989
rect 217715 280961 217749 280989
rect 217777 280961 217811 280989
rect 217839 280961 226625 280989
rect 226653 280961 226687 280989
rect 226715 280961 226749 280989
rect 226777 280961 226811 280989
rect 226839 280961 235625 280989
rect 235653 280961 235687 280989
rect 235715 280961 235749 280989
rect 235777 280961 235811 280989
rect 235839 280961 244625 280989
rect 244653 280961 244687 280989
rect 244715 280961 244749 280989
rect 244777 280961 244811 280989
rect 244839 280961 253625 280989
rect 253653 280961 253687 280989
rect 253715 280961 253749 280989
rect 253777 280961 253811 280989
rect 253839 280961 262625 280989
rect 262653 280961 262687 280989
rect 262715 280961 262749 280989
rect 262777 280961 262811 280989
rect 262839 280961 271625 280989
rect 271653 280961 271687 280989
rect 271715 280961 271749 280989
rect 271777 280961 271811 280989
rect 271839 280961 280625 280989
rect 280653 280961 280687 280989
rect 280715 280961 280749 280989
rect 280777 280961 280811 280989
rect 280839 280961 289625 280989
rect 289653 280961 289687 280989
rect 289715 280961 289749 280989
rect 289777 280961 289811 280989
rect 289839 280961 298248 280989
rect 298276 280961 298310 280989
rect 298338 280961 298372 280989
rect 298400 280961 298434 280989
rect 298462 280961 298990 280989
rect -958 280913 298990 280961
rect -958 275175 298990 275223
rect -958 275147 -910 275175
rect -882 275147 -848 275175
rect -820 275147 -786 275175
rect -758 275147 -724 275175
rect -696 275147 3485 275175
rect 3513 275147 3547 275175
rect 3575 275147 3609 275175
rect 3637 275147 3671 275175
rect 3699 275147 12485 275175
rect 12513 275147 12547 275175
rect 12575 275147 12609 275175
rect 12637 275147 12671 275175
rect 12699 275147 21485 275175
rect 21513 275147 21547 275175
rect 21575 275147 21609 275175
rect 21637 275147 21671 275175
rect 21699 275147 30485 275175
rect 30513 275147 30547 275175
rect 30575 275147 30609 275175
rect 30637 275147 30671 275175
rect 30699 275147 39485 275175
rect 39513 275147 39547 275175
rect 39575 275147 39609 275175
rect 39637 275147 39671 275175
rect 39699 275147 48485 275175
rect 48513 275147 48547 275175
rect 48575 275147 48609 275175
rect 48637 275147 48671 275175
rect 48699 275147 57485 275175
rect 57513 275147 57547 275175
rect 57575 275147 57609 275175
rect 57637 275147 57671 275175
rect 57699 275147 66485 275175
rect 66513 275147 66547 275175
rect 66575 275147 66609 275175
rect 66637 275147 66671 275175
rect 66699 275147 75485 275175
rect 75513 275147 75547 275175
rect 75575 275147 75609 275175
rect 75637 275147 75671 275175
rect 75699 275147 84485 275175
rect 84513 275147 84547 275175
rect 84575 275147 84609 275175
rect 84637 275147 84671 275175
rect 84699 275147 93485 275175
rect 93513 275147 93547 275175
rect 93575 275147 93609 275175
rect 93637 275147 93671 275175
rect 93699 275147 102485 275175
rect 102513 275147 102547 275175
rect 102575 275147 102609 275175
rect 102637 275147 102671 275175
rect 102699 275147 111485 275175
rect 111513 275147 111547 275175
rect 111575 275147 111609 275175
rect 111637 275147 111671 275175
rect 111699 275147 120485 275175
rect 120513 275147 120547 275175
rect 120575 275147 120609 275175
rect 120637 275147 120671 275175
rect 120699 275147 129485 275175
rect 129513 275147 129547 275175
rect 129575 275147 129609 275175
rect 129637 275147 129671 275175
rect 129699 275147 138485 275175
rect 138513 275147 138547 275175
rect 138575 275147 138609 275175
rect 138637 275147 138671 275175
rect 138699 275147 147485 275175
rect 147513 275147 147547 275175
rect 147575 275147 147609 275175
rect 147637 275147 147671 275175
rect 147699 275147 156485 275175
rect 156513 275147 156547 275175
rect 156575 275147 156609 275175
rect 156637 275147 156671 275175
rect 156699 275147 165485 275175
rect 165513 275147 165547 275175
rect 165575 275147 165609 275175
rect 165637 275147 165671 275175
rect 165699 275147 174485 275175
rect 174513 275147 174547 275175
rect 174575 275147 174609 275175
rect 174637 275147 174671 275175
rect 174699 275147 183485 275175
rect 183513 275147 183547 275175
rect 183575 275147 183609 275175
rect 183637 275147 183671 275175
rect 183699 275147 192485 275175
rect 192513 275147 192547 275175
rect 192575 275147 192609 275175
rect 192637 275147 192671 275175
rect 192699 275147 201485 275175
rect 201513 275147 201547 275175
rect 201575 275147 201609 275175
rect 201637 275147 201671 275175
rect 201699 275147 210485 275175
rect 210513 275147 210547 275175
rect 210575 275147 210609 275175
rect 210637 275147 210671 275175
rect 210699 275147 219485 275175
rect 219513 275147 219547 275175
rect 219575 275147 219609 275175
rect 219637 275147 219671 275175
rect 219699 275147 228485 275175
rect 228513 275147 228547 275175
rect 228575 275147 228609 275175
rect 228637 275147 228671 275175
rect 228699 275147 237485 275175
rect 237513 275147 237547 275175
rect 237575 275147 237609 275175
rect 237637 275147 237671 275175
rect 237699 275147 246485 275175
rect 246513 275147 246547 275175
rect 246575 275147 246609 275175
rect 246637 275147 246671 275175
rect 246699 275147 255485 275175
rect 255513 275147 255547 275175
rect 255575 275147 255609 275175
rect 255637 275147 255671 275175
rect 255699 275147 264485 275175
rect 264513 275147 264547 275175
rect 264575 275147 264609 275175
rect 264637 275147 264671 275175
rect 264699 275147 273485 275175
rect 273513 275147 273547 275175
rect 273575 275147 273609 275175
rect 273637 275147 273671 275175
rect 273699 275147 282485 275175
rect 282513 275147 282547 275175
rect 282575 275147 282609 275175
rect 282637 275147 282671 275175
rect 282699 275147 291485 275175
rect 291513 275147 291547 275175
rect 291575 275147 291609 275175
rect 291637 275147 291671 275175
rect 291699 275147 298728 275175
rect 298756 275147 298790 275175
rect 298818 275147 298852 275175
rect 298880 275147 298914 275175
rect 298942 275147 298990 275175
rect -958 275113 298990 275147
rect -958 275085 -910 275113
rect -882 275085 -848 275113
rect -820 275085 -786 275113
rect -758 275085 -724 275113
rect -696 275085 3485 275113
rect 3513 275085 3547 275113
rect 3575 275085 3609 275113
rect 3637 275085 3671 275113
rect 3699 275085 12485 275113
rect 12513 275085 12547 275113
rect 12575 275085 12609 275113
rect 12637 275085 12671 275113
rect 12699 275085 21485 275113
rect 21513 275085 21547 275113
rect 21575 275085 21609 275113
rect 21637 275085 21671 275113
rect 21699 275085 30485 275113
rect 30513 275085 30547 275113
rect 30575 275085 30609 275113
rect 30637 275085 30671 275113
rect 30699 275085 39485 275113
rect 39513 275085 39547 275113
rect 39575 275085 39609 275113
rect 39637 275085 39671 275113
rect 39699 275085 48485 275113
rect 48513 275085 48547 275113
rect 48575 275085 48609 275113
rect 48637 275085 48671 275113
rect 48699 275085 57485 275113
rect 57513 275085 57547 275113
rect 57575 275085 57609 275113
rect 57637 275085 57671 275113
rect 57699 275085 66485 275113
rect 66513 275085 66547 275113
rect 66575 275085 66609 275113
rect 66637 275085 66671 275113
rect 66699 275085 75485 275113
rect 75513 275085 75547 275113
rect 75575 275085 75609 275113
rect 75637 275085 75671 275113
rect 75699 275085 84485 275113
rect 84513 275085 84547 275113
rect 84575 275085 84609 275113
rect 84637 275085 84671 275113
rect 84699 275085 93485 275113
rect 93513 275085 93547 275113
rect 93575 275085 93609 275113
rect 93637 275085 93671 275113
rect 93699 275085 102485 275113
rect 102513 275085 102547 275113
rect 102575 275085 102609 275113
rect 102637 275085 102671 275113
rect 102699 275085 111485 275113
rect 111513 275085 111547 275113
rect 111575 275085 111609 275113
rect 111637 275085 111671 275113
rect 111699 275085 120485 275113
rect 120513 275085 120547 275113
rect 120575 275085 120609 275113
rect 120637 275085 120671 275113
rect 120699 275085 129485 275113
rect 129513 275085 129547 275113
rect 129575 275085 129609 275113
rect 129637 275085 129671 275113
rect 129699 275085 138485 275113
rect 138513 275085 138547 275113
rect 138575 275085 138609 275113
rect 138637 275085 138671 275113
rect 138699 275085 147485 275113
rect 147513 275085 147547 275113
rect 147575 275085 147609 275113
rect 147637 275085 147671 275113
rect 147699 275085 156485 275113
rect 156513 275085 156547 275113
rect 156575 275085 156609 275113
rect 156637 275085 156671 275113
rect 156699 275085 165485 275113
rect 165513 275085 165547 275113
rect 165575 275085 165609 275113
rect 165637 275085 165671 275113
rect 165699 275085 174485 275113
rect 174513 275085 174547 275113
rect 174575 275085 174609 275113
rect 174637 275085 174671 275113
rect 174699 275085 183485 275113
rect 183513 275085 183547 275113
rect 183575 275085 183609 275113
rect 183637 275085 183671 275113
rect 183699 275085 192485 275113
rect 192513 275085 192547 275113
rect 192575 275085 192609 275113
rect 192637 275085 192671 275113
rect 192699 275085 201485 275113
rect 201513 275085 201547 275113
rect 201575 275085 201609 275113
rect 201637 275085 201671 275113
rect 201699 275085 210485 275113
rect 210513 275085 210547 275113
rect 210575 275085 210609 275113
rect 210637 275085 210671 275113
rect 210699 275085 219485 275113
rect 219513 275085 219547 275113
rect 219575 275085 219609 275113
rect 219637 275085 219671 275113
rect 219699 275085 228485 275113
rect 228513 275085 228547 275113
rect 228575 275085 228609 275113
rect 228637 275085 228671 275113
rect 228699 275085 237485 275113
rect 237513 275085 237547 275113
rect 237575 275085 237609 275113
rect 237637 275085 237671 275113
rect 237699 275085 246485 275113
rect 246513 275085 246547 275113
rect 246575 275085 246609 275113
rect 246637 275085 246671 275113
rect 246699 275085 255485 275113
rect 255513 275085 255547 275113
rect 255575 275085 255609 275113
rect 255637 275085 255671 275113
rect 255699 275085 264485 275113
rect 264513 275085 264547 275113
rect 264575 275085 264609 275113
rect 264637 275085 264671 275113
rect 264699 275085 273485 275113
rect 273513 275085 273547 275113
rect 273575 275085 273609 275113
rect 273637 275085 273671 275113
rect 273699 275085 282485 275113
rect 282513 275085 282547 275113
rect 282575 275085 282609 275113
rect 282637 275085 282671 275113
rect 282699 275085 291485 275113
rect 291513 275085 291547 275113
rect 291575 275085 291609 275113
rect 291637 275085 291671 275113
rect 291699 275085 298728 275113
rect 298756 275085 298790 275113
rect 298818 275085 298852 275113
rect 298880 275085 298914 275113
rect 298942 275085 298990 275113
rect -958 275051 298990 275085
rect -958 275023 -910 275051
rect -882 275023 -848 275051
rect -820 275023 -786 275051
rect -758 275023 -724 275051
rect -696 275023 3485 275051
rect 3513 275023 3547 275051
rect 3575 275023 3609 275051
rect 3637 275023 3671 275051
rect 3699 275023 12485 275051
rect 12513 275023 12547 275051
rect 12575 275023 12609 275051
rect 12637 275023 12671 275051
rect 12699 275023 21485 275051
rect 21513 275023 21547 275051
rect 21575 275023 21609 275051
rect 21637 275023 21671 275051
rect 21699 275023 30485 275051
rect 30513 275023 30547 275051
rect 30575 275023 30609 275051
rect 30637 275023 30671 275051
rect 30699 275023 39485 275051
rect 39513 275023 39547 275051
rect 39575 275023 39609 275051
rect 39637 275023 39671 275051
rect 39699 275023 48485 275051
rect 48513 275023 48547 275051
rect 48575 275023 48609 275051
rect 48637 275023 48671 275051
rect 48699 275023 57485 275051
rect 57513 275023 57547 275051
rect 57575 275023 57609 275051
rect 57637 275023 57671 275051
rect 57699 275023 66485 275051
rect 66513 275023 66547 275051
rect 66575 275023 66609 275051
rect 66637 275023 66671 275051
rect 66699 275023 75485 275051
rect 75513 275023 75547 275051
rect 75575 275023 75609 275051
rect 75637 275023 75671 275051
rect 75699 275023 84485 275051
rect 84513 275023 84547 275051
rect 84575 275023 84609 275051
rect 84637 275023 84671 275051
rect 84699 275023 93485 275051
rect 93513 275023 93547 275051
rect 93575 275023 93609 275051
rect 93637 275023 93671 275051
rect 93699 275023 102485 275051
rect 102513 275023 102547 275051
rect 102575 275023 102609 275051
rect 102637 275023 102671 275051
rect 102699 275023 111485 275051
rect 111513 275023 111547 275051
rect 111575 275023 111609 275051
rect 111637 275023 111671 275051
rect 111699 275023 120485 275051
rect 120513 275023 120547 275051
rect 120575 275023 120609 275051
rect 120637 275023 120671 275051
rect 120699 275023 129485 275051
rect 129513 275023 129547 275051
rect 129575 275023 129609 275051
rect 129637 275023 129671 275051
rect 129699 275023 138485 275051
rect 138513 275023 138547 275051
rect 138575 275023 138609 275051
rect 138637 275023 138671 275051
rect 138699 275023 147485 275051
rect 147513 275023 147547 275051
rect 147575 275023 147609 275051
rect 147637 275023 147671 275051
rect 147699 275023 156485 275051
rect 156513 275023 156547 275051
rect 156575 275023 156609 275051
rect 156637 275023 156671 275051
rect 156699 275023 165485 275051
rect 165513 275023 165547 275051
rect 165575 275023 165609 275051
rect 165637 275023 165671 275051
rect 165699 275023 174485 275051
rect 174513 275023 174547 275051
rect 174575 275023 174609 275051
rect 174637 275023 174671 275051
rect 174699 275023 183485 275051
rect 183513 275023 183547 275051
rect 183575 275023 183609 275051
rect 183637 275023 183671 275051
rect 183699 275023 192485 275051
rect 192513 275023 192547 275051
rect 192575 275023 192609 275051
rect 192637 275023 192671 275051
rect 192699 275023 201485 275051
rect 201513 275023 201547 275051
rect 201575 275023 201609 275051
rect 201637 275023 201671 275051
rect 201699 275023 210485 275051
rect 210513 275023 210547 275051
rect 210575 275023 210609 275051
rect 210637 275023 210671 275051
rect 210699 275023 219485 275051
rect 219513 275023 219547 275051
rect 219575 275023 219609 275051
rect 219637 275023 219671 275051
rect 219699 275023 228485 275051
rect 228513 275023 228547 275051
rect 228575 275023 228609 275051
rect 228637 275023 228671 275051
rect 228699 275023 237485 275051
rect 237513 275023 237547 275051
rect 237575 275023 237609 275051
rect 237637 275023 237671 275051
rect 237699 275023 246485 275051
rect 246513 275023 246547 275051
rect 246575 275023 246609 275051
rect 246637 275023 246671 275051
rect 246699 275023 255485 275051
rect 255513 275023 255547 275051
rect 255575 275023 255609 275051
rect 255637 275023 255671 275051
rect 255699 275023 264485 275051
rect 264513 275023 264547 275051
rect 264575 275023 264609 275051
rect 264637 275023 264671 275051
rect 264699 275023 273485 275051
rect 273513 275023 273547 275051
rect 273575 275023 273609 275051
rect 273637 275023 273671 275051
rect 273699 275023 282485 275051
rect 282513 275023 282547 275051
rect 282575 275023 282609 275051
rect 282637 275023 282671 275051
rect 282699 275023 291485 275051
rect 291513 275023 291547 275051
rect 291575 275023 291609 275051
rect 291637 275023 291671 275051
rect 291699 275023 298728 275051
rect 298756 275023 298790 275051
rect 298818 275023 298852 275051
rect 298880 275023 298914 275051
rect 298942 275023 298990 275051
rect -958 274989 298990 275023
rect -958 274961 -910 274989
rect -882 274961 -848 274989
rect -820 274961 -786 274989
rect -758 274961 -724 274989
rect -696 274961 3485 274989
rect 3513 274961 3547 274989
rect 3575 274961 3609 274989
rect 3637 274961 3671 274989
rect 3699 274961 12485 274989
rect 12513 274961 12547 274989
rect 12575 274961 12609 274989
rect 12637 274961 12671 274989
rect 12699 274961 21485 274989
rect 21513 274961 21547 274989
rect 21575 274961 21609 274989
rect 21637 274961 21671 274989
rect 21699 274961 30485 274989
rect 30513 274961 30547 274989
rect 30575 274961 30609 274989
rect 30637 274961 30671 274989
rect 30699 274961 39485 274989
rect 39513 274961 39547 274989
rect 39575 274961 39609 274989
rect 39637 274961 39671 274989
rect 39699 274961 48485 274989
rect 48513 274961 48547 274989
rect 48575 274961 48609 274989
rect 48637 274961 48671 274989
rect 48699 274961 57485 274989
rect 57513 274961 57547 274989
rect 57575 274961 57609 274989
rect 57637 274961 57671 274989
rect 57699 274961 66485 274989
rect 66513 274961 66547 274989
rect 66575 274961 66609 274989
rect 66637 274961 66671 274989
rect 66699 274961 75485 274989
rect 75513 274961 75547 274989
rect 75575 274961 75609 274989
rect 75637 274961 75671 274989
rect 75699 274961 84485 274989
rect 84513 274961 84547 274989
rect 84575 274961 84609 274989
rect 84637 274961 84671 274989
rect 84699 274961 93485 274989
rect 93513 274961 93547 274989
rect 93575 274961 93609 274989
rect 93637 274961 93671 274989
rect 93699 274961 102485 274989
rect 102513 274961 102547 274989
rect 102575 274961 102609 274989
rect 102637 274961 102671 274989
rect 102699 274961 111485 274989
rect 111513 274961 111547 274989
rect 111575 274961 111609 274989
rect 111637 274961 111671 274989
rect 111699 274961 120485 274989
rect 120513 274961 120547 274989
rect 120575 274961 120609 274989
rect 120637 274961 120671 274989
rect 120699 274961 129485 274989
rect 129513 274961 129547 274989
rect 129575 274961 129609 274989
rect 129637 274961 129671 274989
rect 129699 274961 138485 274989
rect 138513 274961 138547 274989
rect 138575 274961 138609 274989
rect 138637 274961 138671 274989
rect 138699 274961 147485 274989
rect 147513 274961 147547 274989
rect 147575 274961 147609 274989
rect 147637 274961 147671 274989
rect 147699 274961 156485 274989
rect 156513 274961 156547 274989
rect 156575 274961 156609 274989
rect 156637 274961 156671 274989
rect 156699 274961 165485 274989
rect 165513 274961 165547 274989
rect 165575 274961 165609 274989
rect 165637 274961 165671 274989
rect 165699 274961 174485 274989
rect 174513 274961 174547 274989
rect 174575 274961 174609 274989
rect 174637 274961 174671 274989
rect 174699 274961 183485 274989
rect 183513 274961 183547 274989
rect 183575 274961 183609 274989
rect 183637 274961 183671 274989
rect 183699 274961 192485 274989
rect 192513 274961 192547 274989
rect 192575 274961 192609 274989
rect 192637 274961 192671 274989
rect 192699 274961 201485 274989
rect 201513 274961 201547 274989
rect 201575 274961 201609 274989
rect 201637 274961 201671 274989
rect 201699 274961 210485 274989
rect 210513 274961 210547 274989
rect 210575 274961 210609 274989
rect 210637 274961 210671 274989
rect 210699 274961 219485 274989
rect 219513 274961 219547 274989
rect 219575 274961 219609 274989
rect 219637 274961 219671 274989
rect 219699 274961 228485 274989
rect 228513 274961 228547 274989
rect 228575 274961 228609 274989
rect 228637 274961 228671 274989
rect 228699 274961 237485 274989
rect 237513 274961 237547 274989
rect 237575 274961 237609 274989
rect 237637 274961 237671 274989
rect 237699 274961 246485 274989
rect 246513 274961 246547 274989
rect 246575 274961 246609 274989
rect 246637 274961 246671 274989
rect 246699 274961 255485 274989
rect 255513 274961 255547 274989
rect 255575 274961 255609 274989
rect 255637 274961 255671 274989
rect 255699 274961 264485 274989
rect 264513 274961 264547 274989
rect 264575 274961 264609 274989
rect 264637 274961 264671 274989
rect 264699 274961 273485 274989
rect 273513 274961 273547 274989
rect 273575 274961 273609 274989
rect 273637 274961 273671 274989
rect 273699 274961 282485 274989
rect 282513 274961 282547 274989
rect 282575 274961 282609 274989
rect 282637 274961 282671 274989
rect 282699 274961 291485 274989
rect 291513 274961 291547 274989
rect 291575 274961 291609 274989
rect 291637 274961 291671 274989
rect 291699 274961 298728 274989
rect 298756 274961 298790 274989
rect 298818 274961 298852 274989
rect 298880 274961 298914 274989
rect 298942 274961 298990 274989
rect -958 274913 298990 274961
rect -958 272175 298990 272223
rect -958 272147 -430 272175
rect -402 272147 -368 272175
rect -340 272147 -306 272175
rect -278 272147 -244 272175
rect -216 272147 1625 272175
rect 1653 272147 1687 272175
rect 1715 272147 1749 272175
rect 1777 272147 1811 272175
rect 1839 272147 10625 272175
rect 10653 272147 10687 272175
rect 10715 272147 10749 272175
rect 10777 272147 10811 272175
rect 10839 272147 19625 272175
rect 19653 272147 19687 272175
rect 19715 272147 19749 272175
rect 19777 272147 19811 272175
rect 19839 272147 28625 272175
rect 28653 272147 28687 272175
rect 28715 272147 28749 272175
rect 28777 272147 28811 272175
rect 28839 272147 37625 272175
rect 37653 272147 37687 272175
rect 37715 272147 37749 272175
rect 37777 272147 37811 272175
rect 37839 272147 46625 272175
rect 46653 272147 46687 272175
rect 46715 272147 46749 272175
rect 46777 272147 46811 272175
rect 46839 272147 55625 272175
rect 55653 272147 55687 272175
rect 55715 272147 55749 272175
rect 55777 272147 55811 272175
rect 55839 272147 64625 272175
rect 64653 272147 64687 272175
rect 64715 272147 64749 272175
rect 64777 272147 64811 272175
rect 64839 272147 73625 272175
rect 73653 272147 73687 272175
rect 73715 272147 73749 272175
rect 73777 272147 73811 272175
rect 73839 272147 82625 272175
rect 82653 272147 82687 272175
rect 82715 272147 82749 272175
rect 82777 272147 82811 272175
rect 82839 272147 91625 272175
rect 91653 272147 91687 272175
rect 91715 272147 91749 272175
rect 91777 272147 91811 272175
rect 91839 272147 100625 272175
rect 100653 272147 100687 272175
rect 100715 272147 100749 272175
rect 100777 272147 100811 272175
rect 100839 272147 109625 272175
rect 109653 272147 109687 272175
rect 109715 272147 109749 272175
rect 109777 272147 109811 272175
rect 109839 272147 118625 272175
rect 118653 272147 118687 272175
rect 118715 272147 118749 272175
rect 118777 272147 118811 272175
rect 118839 272147 127625 272175
rect 127653 272147 127687 272175
rect 127715 272147 127749 272175
rect 127777 272147 127811 272175
rect 127839 272147 136625 272175
rect 136653 272147 136687 272175
rect 136715 272147 136749 272175
rect 136777 272147 136811 272175
rect 136839 272147 145625 272175
rect 145653 272147 145687 272175
rect 145715 272147 145749 272175
rect 145777 272147 145811 272175
rect 145839 272147 154625 272175
rect 154653 272147 154687 272175
rect 154715 272147 154749 272175
rect 154777 272147 154811 272175
rect 154839 272147 163625 272175
rect 163653 272147 163687 272175
rect 163715 272147 163749 272175
rect 163777 272147 163811 272175
rect 163839 272147 172625 272175
rect 172653 272147 172687 272175
rect 172715 272147 172749 272175
rect 172777 272147 172811 272175
rect 172839 272147 181625 272175
rect 181653 272147 181687 272175
rect 181715 272147 181749 272175
rect 181777 272147 181811 272175
rect 181839 272147 190625 272175
rect 190653 272147 190687 272175
rect 190715 272147 190749 272175
rect 190777 272147 190811 272175
rect 190839 272147 199625 272175
rect 199653 272147 199687 272175
rect 199715 272147 199749 272175
rect 199777 272147 199811 272175
rect 199839 272147 208625 272175
rect 208653 272147 208687 272175
rect 208715 272147 208749 272175
rect 208777 272147 208811 272175
rect 208839 272147 217625 272175
rect 217653 272147 217687 272175
rect 217715 272147 217749 272175
rect 217777 272147 217811 272175
rect 217839 272147 226625 272175
rect 226653 272147 226687 272175
rect 226715 272147 226749 272175
rect 226777 272147 226811 272175
rect 226839 272147 235625 272175
rect 235653 272147 235687 272175
rect 235715 272147 235749 272175
rect 235777 272147 235811 272175
rect 235839 272147 244625 272175
rect 244653 272147 244687 272175
rect 244715 272147 244749 272175
rect 244777 272147 244811 272175
rect 244839 272147 253625 272175
rect 253653 272147 253687 272175
rect 253715 272147 253749 272175
rect 253777 272147 253811 272175
rect 253839 272147 262625 272175
rect 262653 272147 262687 272175
rect 262715 272147 262749 272175
rect 262777 272147 262811 272175
rect 262839 272147 271625 272175
rect 271653 272147 271687 272175
rect 271715 272147 271749 272175
rect 271777 272147 271811 272175
rect 271839 272147 280625 272175
rect 280653 272147 280687 272175
rect 280715 272147 280749 272175
rect 280777 272147 280811 272175
rect 280839 272147 289625 272175
rect 289653 272147 289687 272175
rect 289715 272147 289749 272175
rect 289777 272147 289811 272175
rect 289839 272147 298248 272175
rect 298276 272147 298310 272175
rect 298338 272147 298372 272175
rect 298400 272147 298434 272175
rect 298462 272147 298990 272175
rect -958 272113 298990 272147
rect -958 272085 -430 272113
rect -402 272085 -368 272113
rect -340 272085 -306 272113
rect -278 272085 -244 272113
rect -216 272085 1625 272113
rect 1653 272085 1687 272113
rect 1715 272085 1749 272113
rect 1777 272085 1811 272113
rect 1839 272085 10625 272113
rect 10653 272085 10687 272113
rect 10715 272085 10749 272113
rect 10777 272085 10811 272113
rect 10839 272085 19625 272113
rect 19653 272085 19687 272113
rect 19715 272085 19749 272113
rect 19777 272085 19811 272113
rect 19839 272085 28625 272113
rect 28653 272085 28687 272113
rect 28715 272085 28749 272113
rect 28777 272085 28811 272113
rect 28839 272085 37625 272113
rect 37653 272085 37687 272113
rect 37715 272085 37749 272113
rect 37777 272085 37811 272113
rect 37839 272085 46625 272113
rect 46653 272085 46687 272113
rect 46715 272085 46749 272113
rect 46777 272085 46811 272113
rect 46839 272085 55625 272113
rect 55653 272085 55687 272113
rect 55715 272085 55749 272113
rect 55777 272085 55811 272113
rect 55839 272085 64625 272113
rect 64653 272085 64687 272113
rect 64715 272085 64749 272113
rect 64777 272085 64811 272113
rect 64839 272085 73625 272113
rect 73653 272085 73687 272113
rect 73715 272085 73749 272113
rect 73777 272085 73811 272113
rect 73839 272085 82625 272113
rect 82653 272085 82687 272113
rect 82715 272085 82749 272113
rect 82777 272085 82811 272113
rect 82839 272085 91625 272113
rect 91653 272085 91687 272113
rect 91715 272085 91749 272113
rect 91777 272085 91811 272113
rect 91839 272085 100625 272113
rect 100653 272085 100687 272113
rect 100715 272085 100749 272113
rect 100777 272085 100811 272113
rect 100839 272085 109625 272113
rect 109653 272085 109687 272113
rect 109715 272085 109749 272113
rect 109777 272085 109811 272113
rect 109839 272085 118625 272113
rect 118653 272085 118687 272113
rect 118715 272085 118749 272113
rect 118777 272085 118811 272113
rect 118839 272085 127625 272113
rect 127653 272085 127687 272113
rect 127715 272085 127749 272113
rect 127777 272085 127811 272113
rect 127839 272085 136625 272113
rect 136653 272085 136687 272113
rect 136715 272085 136749 272113
rect 136777 272085 136811 272113
rect 136839 272085 145625 272113
rect 145653 272085 145687 272113
rect 145715 272085 145749 272113
rect 145777 272085 145811 272113
rect 145839 272085 154625 272113
rect 154653 272085 154687 272113
rect 154715 272085 154749 272113
rect 154777 272085 154811 272113
rect 154839 272085 163625 272113
rect 163653 272085 163687 272113
rect 163715 272085 163749 272113
rect 163777 272085 163811 272113
rect 163839 272085 172625 272113
rect 172653 272085 172687 272113
rect 172715 272085 172749 272113
rect 172777 272085 172811 272113
rect 172839 272085 181625 272113
rect 181653 272085 181687 272113
rect 181715 272085 181749 272113
rect 181777 272085 181811 272113
rect 181839 272085 190625 272113
rect 190653 272085 190687 272113
rect 190715 272085 190749 272113
rect 190777 272085 190811 272113
rect 190839 272085 199625 272113
rect 199653 272085 199687 272113
rect 199715 272085 199749 272113
rect 199777 272085 199811 272113
rect 199839 272085 208625 272113
rect 208653 272085 208687 272113
rect 208715 272085 208749 272113
rect 208777 272085 208811 272113
rect 208839 272085 217625 272113
rect 217653 272085 217687 272113
rect 217715 272085 217749 272113
rect 217777 272085 217811 272113
rect 217839 272085 226625 272113
rect 226653 272085 226687 272113
rect 226715 272085 226749 272113
rect 226777 272085 226811 272113
rect 226839 272085 235625 272113
rect 235653 272085 235687 272113
rect 235715 272085 235749 272113
rect 235777 272085 235811 272113
rect 235839 272085 244625 272113
rect 244653 272085 244687 272113
rect 244715 272085 244749 272113
rect 244777 272085 244811 272113
rect 244839 272085 253625 272113
rect 253653 272085 253687 272113
rect 253715 272085 253749 272113
rect 253777 272085 253811 272113
rect 253839 272085 262625 272113
rect 262653 272085 262687 272113
rect 262715 272085 262749 272113
rect 262777 272085 262811 272113
rect 262839 272085 271625 272113
rect 271653 272085 271687 272113
rect 271715 272085 271749 272113
rect 271777 272085 271811 272113
rect 271839 272085 280625 272113
rect 280653 272085 280687 272113
rect 280715 272085 280749 272113
rect 280777 272085 280811 272113
rect 280839 272085 289625 272113
rect 289653 272085 289687 272113
rect 289715 272085 289749 272113
rect 289777 272085 289811 272113
rect 289839 272085 298248 272113
rect 298276 272085 298310 272113
rect 298338 272085 298372 272113
rect 298400 272085 298434 272113
rect 298462 272085 298990 272113
rect -958 272051 298990 272085
rect -958 272023 -430 272051
rect -402 272023 -368 272051
rect -340 272023 -306 272051
rect -278 272023 -244 272051
rect -216 272023 1625 272051
rect 1653 272023 1687 272051
rect 1715 272023 1749 272051
rect 1777 272023 1811 272051
rect 1839 272023 10625 272051
rect 10653 272023 10687 272051
rect 10715 272023 10749 272051
rect 10777 272023 10811 272051
rect 10839 272023 19625 272051
rect 19653 272023 19687 272051
rect 19715 272023 19749 272051
rect 19777 272023 19811 272051
rect 19839 272023 28625 272051
rect 28653 272023 28687 272051
rect 28715 272023 28749 272051
rect 28777 272023 28811 272051
rect 28839 272023 37625 272051
rect 37653 272023 37687 272051
rect 37715 272023 37749 272051
rect 37777 272023 37811 272051
rect 37839 272023 46625 272051
rect 46653 272023 46687 272051
rect 46715 272023 46749 272051
rect 46777 272023 46811 272051
rect 46839 272023 55625 272051
rect 55653 272023 55687 272051
rect 55715 272023 55749 272051
rect 55777 272023 55811 272051
rect 55839 272023 64625 272051
rect 64653 272023 64687 272051
rect 64715 272023 64749 272051
rect 64777 272023 64811 272051
rect 64839 272023 73625 272051
rect 73653 272023 73687 272051
rect 73715 272023 73749 272051
rect 73777 272023 73811 272051
rect 73839 272023 82625 272051
rect 82653 272023 82687 272051
rect 82715 272023 82749 272051
rect 82777 272023 82811 272051
rect 82839 272023 91625 272051
rect 91653 272023 91687 272051
rect 91715 272023 91749 272051
rect 91777 272023 91811 272051
rect 91839 272023 100625 272051
rect 100653 272023 100687 272051
rect 100715 272023 100749 272051
rect 100777 272023 100811 272051
rect 100839 272023 109625 272051
rect 109653 272023 109687 272051
rect 109715 272023 109749 272051
rect 109777 272023 109811 272051
rect 109839 272023 118625 272051
rect 118653 272023 118687 272051
rect 118715 272023 118749 272051
rect 118777 272023 118811 272051
rect 118839 272023 127625 272051
rect 127653 272023 127687 272051
rect 127715 272023 127749 272051
rect 127777 272023 127811 272051
rect 127839 272023 136625 272051
rect 136653 272023 136687 272051
rect 136715 272023 136749 272051
rect 136777 272023 136811 272051
rect 136839 272023 145625 272051
rect 145653 272023 145687 272051
rect 145715 272023 145749 272051
rect 145777 272023 145811 272051
rect 145839 272023 154625 272051
rect 154653 272023 154687 272051
rect 154715 272023 154749 272051
rect 154777 272023 154811 272051
rect 154839 272023 163625 272051
rect 163653 272023 163687 272051
rect 163715 272023 163749 272051
rect 163777 272023 163811 272051
rect 163839 272023 172625 272051
rect 172653 272023 172687 272051
rect 172715 272023 172749 272051
rect 172777 272023 172811 272051
rect 172839 272023 181625 272051
rect 181653 272023 181687 272051
rect 181715 272023 181749 272051
rect 181777 272023 181811 272051
rect 181839 272023 190625 272051
rect 190653 272023 190687 272051
rect 190715 272023 190749 272051
rect 190777 272023 190811 272051
rect 190839 272023 199625 272051
rect 199653 272023 199687 272051
rect 199715 272023 199749 272051
rect 199777 272023 199811 272051
rect 199839 272023 208625 272051
rect 208653 272023 208687 272051
rect 208715 272023 208749 272051
rect 208777 272023 208811 272051
rect 208839 272023 217625 272051
rect 217653 272023 217687 272051
rect 217715 272023 217749 272051
rect 217777 272023 217811 272051
rect 217839 272023 226625 272051
rect 226653 272023 226687 272051
rect 226715 272023 226749 272051
rect 226777 272023 226811 272051
rect 226839 272023 235625 272051
rect 235653 272023 235687 272051
rect 235715 272023 235749 272051
rect 235777 272023 235811 272051
rect 235839 272023 244625 272051
rect 244653 272023 244687 272051
rect 244715 272023 244749 272051
rect 244777 272023 244811 272051
rect 244839 272023 253625 272051
rect 253653 272023 253687 272051
rect 253715 272023 253749 272051
rect 253777 272023 253811 272051
rect 253839 272023 262625 272051
rect 262653 272023 262687 272051
rect 262715 272023 262749 272051
rect 262777 272023 262811 272051
rect 262839 272023 271625 272051
rect 271653 272023 271687 272051
rect 271715 272023 271749 272051
rect 271777 272023 271811 272051
rect 271839 272023 280625 272051
rect 280653 272023 280687 272051
rect 280715 272023 280749 272051
rect 280777 272023 280811 272051
rect 280839 272023 289625 272051
rect 289653 272023 289687 272051
rect 289715 272023 289749 272051
rect 289777 272023 289811 272051
rect 289839 272023 298248 272051
rect 298276 272023 298310 272051
rect 298338 272023 298372 272051
rect 298400 272023 298434 272051
rect 298462 272023 298990 272051
rect -958 271989 298990 272023
rect -958 271961 -430 271989
rect -402 271961 -368 271989
rect -340 271961 -306 271989
rect -278 271961 -244 271989
rect -216 271961 1625 271989
rect 1653 271961 1687 271989
rect 1715 271961 1749 271989
rect 1777 271961 1811 271989
rect 1839 271961 10625 271989
rect 10653 271961 10687 271989
rect 10715 271961 10749 271989
rect 10777 271961 10811 271989
rect 10839 271961 19625 271989
rect 19653 271961 19687 271989
rect 19715 271961 19749 271989
rect 19777 271961 19811 271989
rect 19839 271961 28625 271989
rect 28653 271961 28687 271989
rect 28715 271961 28749 271989
rect 28777 271961 28811 271989
rect 28839 271961 37625 271989
rect 37653 271961 37687 271989
rect 37715 271961 37749 271989
rect 37777 271961 37811 271989
rect 37839 271961 46625 271989
rect 46653 271961 46687 271989
rect 46715 271961 46749 271989
rect 46777 271961 46811 271989
rect 46839 271961 55625 271989
rect 55653 271961 55687 271989
rect 55715 271961 55749 271989
rect 55777 271961 55811 271989
rect 55839 271961 64625 271989
rect 64653 271961 64687 271989
rect 64715 271961 64749 271989
rect 64777 271961 64811 271989
rect 64839 271961 73625 271989
rect 73653 271961 73687 271989
rect 73715 271961 73749 271989
rect 73777 271961 73811 271989
rect 73839 271961 82625 271989
rect 82653 271961 82687 271989
rect 82715 271961 82749 271989
rect 82777 271961 82811 271989
rect 82839 271961 91625 271989
rect 91653 271961 91687 271989
rect 91715 271961 91749 271989
rect 91777 271961 91811 271989
rect 91839 271961 100625 271989
rect 100653 271961 100687 271989
rect 100715 271961 100749 271989
rect 100777 271961 100811 271989
rect 100839 271961 109625 271989
rect 109653 271961 109687 271989
rect 109715 271961 109749 271989
rect 109777 271961 109811 271989
rect 109839 271961 118625 271989
rect 118653 271961 118687 271989
rect 118715 271961 118749 271989
rect 118777 271961 118811 271989
rect 118839 271961 127625 271989
rect 127653 271961 127687 271989
rect 127715 271961 127749 271989
rect 127777 271961 127811 271989
rect 127839 271961 136625 271989
rect 136653 271961 136687 271989
rect 136715 271961 136749 271989
rect 136777 271961 136811 271989
rect 136839 271961 145625 271989
rect 145653 271961 145687 271989
rect 145715 271961 145749 271989
rect 145777 271961 145811 271989
rect 145839 271961 154625 271989
rect 154653 271961 154687 271989
rect 154715 271961 154749 271989
rect 154777 271961 154811 271989
rect 154839 271961 163625 271989
rect 163653 271961 163687 271989
rect 163715 271961 163749 271989
rect 163777 271961 163811 271989
rect 163839 271961 172625 271989
rect 172653 271961 172687 271989
rect 172715 271961 172749 271989
rect 172777 271961 172811 271989
rect 172839 271961 181625 271989
rect 181653 271961 181687 271989
rect 181715 271961 181749 271989
rect 181777 271961 181811 271989
rect 181839 271961 190625 271989
rect 190653 271961 190687 271989
rect 190715 271961 190749 271989
rect 190777 271961 190811 271989
rect 190839 271961 199625 271989
rect 199653 271961 199687 271989
rect 199715 271961 199749 271989
rect 199777 271961 199811 271989
rect 199839 271961 208625 271989
rect 208653 271961 208687 271989
rect 208715 271961 208749 271989
rect 208777 271961 208811 271989
rect 208839 271961 217625 271989
rect 217653 271961 217687 271989
rect 217715 271961 217749 271989
rect 217777 271961 217811 271989
rect 217839 271961 226625 271989
rect 226653 271961 226687 271989
rect 226715 271961 226749 271989
rect 226777 271961 226811 271989
rect 226839 271961 235625 271989
rect 235653 271961 235687 271989
rect 235715 271961 235749 271989
rect 235777 271961 235811 271989
rect 235839 271961 244625 271989
rect 244653 271961 244687 271989
rect 244715 271961 244749 271989
rect 244777 271961 244811 271989
rect 244839 271961 253625 271989
rect 253653 271961 253687 271989
rect 253715 271961 253749 271989
rect 253777 271961 253811 271989
rect 253839 271961 262625 271989
rect 262653 271961 262687 271989
rect 262715 271961 262749 271989
rect 262777 271961 262811 271989
rect 262839 271961 271625 271989
rect 271653 271961 271687 271989
rect 271715 271961 271749 271989
rect 271777 271961 271811 271989
rect 271839 271961 280625 271989
rect 280653 271961 280687 271989
rect 280715 271961 280749 271989
rect 280777 271961 280811 271989
rect 280839 271961 289625 271989
rect 289653 271961 289687 271989
rect 289715 271961 289749 271989
rect 289777 271961 289811 271989
rect 289839 271961 298248 271989
rect 298276 271961 298310 271989
rect 298338 271961 298372 271989
rect 298400 271961 298434 271989
rect 298462 271961 298990 271989
rect -958 271913 298990 271961
rect -958 266175 298990 266223
rect -958 266147 -910 266175
rect -882 266147 -848 266175
rect -820 266147 -786 266175
rect -758 266147 -724 266175
rect -696 266147 3485 266175
rect 3513 266147 3547 266175
rect 3575 266147 3609 266175
rect 3637 266147 3671 266175
rect 3699 266147 12485 266175
rect 12513 266147 12547 266175
rect 12575 266147 12609 266175
rect 12637 266147 12671 266175
rect 12699 266147 21485 266175
rect 21513 266147 21547 266175
rect 21575 266147 21609 266175
rect 21637 266147 21671 266175
rect 21699 266147 30485 266175
rect 30513 266147 30547 266175
rect 30575 266147 30609 266175
rect 30637 266147 30671 266175
rect 30699 266147 39485 266175
rect 39513 266147 39547 266175
rect 39575 266147 39609 266175
rect 39637 266147 39671 266175
rect 39699 266147 48485 266175
rect 48513 266147 48547 266175
rect 48575 266147 48609 266175
rect 48637 266147 48671 266175
rect 48699 266147 57485 266175
rect 57513 266147 57547 266175
rect 57575 266147 57609 266175
rect 57637 266147 57671 266175
rect 57699 266147 66485 266175
rect 66513 266147 66547 266175
rect 66575 266147 66609 266175
rect 66637 266147 66671 266175
rect 66699 266147 75485 266175
rect 75513 266147 75547 266175
rect 75575 266147 75609 266175
rect 75637 266147 75671 266175
rect 75699 266147 84485 266175
rect 84513 266147 84547 266175
rect 84575 266147 84609 266175
rect 84637 266147 84671 266175
rect 84699 266147 93485 266175
rect 93513 266147 93547 266175
rect 93575 266147 93609 266175
rect 93637 266147 93671 266175
rect 93699 266147 102485 266175
rect 102513 266147 102547 266175
rect 102575 266147 102609 266175
rect 102637 266147 102671 266175
rect 102699 266147 111485 266175
rect 111513 266147 111547 266175
rect 111575 266147 111609 266175
rect 111637 266147 111671 266175
rect 111699 266147 120485 266175
rect 120513 266147 120547 266175
rect 120575 266147 120609 266175
rect 120637 266147 120671 266175
rect 120699 266147 129485 266175
rect 129513 266147 129547 266175
rect 129575 266147 129609 266175
rect 129637 266147 129671 266175
rect 129699 266147 138485 266175
rect 138513 266147 138547 266175
rect 138575 266147 138609 266175
rect 138637 266147 138671 266175
rect 138699 266147 147485 266175
rect 147513 266147 147547 266175
rect 147575 266147 147609 266175
rect 147637 266147 147671 266175
rect 147699 266147 156485 266175
rect 156513 266147 156547 266175
rect 156575 266147 156609 266175
rect 156637 266147 156671 266175
rect 156699 266147 165485 266175
rect 165513 266147 165547 266175
rect 165575 266147 165609 266175
rect 165637 266147 165671 266175
rect 165699 266147 174485 266175
rect 174513 266147 174547 266175
rect 174575 266147 174609 266175
rect 174637 266147 174671 266175
rect 174699 266147 183485 266175
rect 183513 266147 183547 266175
rect 183575 266147 183609 266175
rect 183637 266147 183671 266175
rect 183699 266147 192485 266175
rect 192513 266147 192547 266175
rect 192575 266147 192609 266175
rect 192637 266147 192671 266175
rect 192699 266147 201485 266175
rect 201513 266147 201547 266175
rect 201575 266147 201609 266175
rect 201637 266147 201671 266175
rect 201699 266147 210485 266175
rect 210513 266147 210547 266175
rect 210575 266147 210609 266175
rect 210637 266147 210671 266175
rect 210699 266147 219485 266175
rect 219513 266147 219547 266175
rect 219575 266147 219609 266175
rect 219637 266147 219671 266175
rect 219699 266147 228485 266175
rect 228513 266147 228547 266175
rect 228575 266147 228609 266175
rect 228637 266147 228671 266175
rect 228699 266147 237485 266175
rect 237513 266147 237547 266175
rect 237575 266147 237609 266175
rect 237637 266147 237671 266175
rect 237699 266147 246485 266175
rect 246513 266147 246547 266175
rect 246575 266147 246609 266175
rect 246637 266147 246671 266175
rect 246699 266147 255485 266175
rect 255513 266147 255547 266175
rect 255575 266147 255609 266175
rect 255637 266147 255671 266175
rect 255699 266147 264485 266175
rect 264513 266147 264547 266175
rect 264575 266147 264609 266175
rect 264637 266147 264671 266175
rect 264699 266147 273485 266175
rect 273513 266147 273547 266175
rect 273575 266147 273609 266175
rect 273637 266147 273671 266175
rect 273699 266147 282485 266175
rect 282513 266147 282547 266175
rect 282575 266147 282609 266175
rect 282637 266147 282671 266175
rect 282699 266147 291485 266175
rect 291513 266147 291547 266175
rect 291575 266147 291609 266175
rect 291637 266147 291671 266175
rect 291699 266147 298728 266175
rect 298756 266147 298790 266175
rect 298818 266147 298852 266175
rect 298880 266147 298914 266175
rect 298942 266147 298990 266175
rect -958 266113 298990 266147
rect -958 266085 -910 266113
rect -882 266085 -848 266113
rect -820 266085 -786 266113
rect -758 266085 -724 266113
rect -696 266085 3485 266113
rect 3513 266085 3547 266113
rect 3575 266085 3609 266113
rect 3637 266085 3671 266113
rect 3699 266085 12485 266113
rect 12513 266085 12547 266113
rect 12575 266085 12609 266113
rect 12637 266085 12671 266113
rect 12699 266085 21485 266113
rect 21513 266085 21547 266113
rect 21575 266085 21609 266113
rect 21637 266085 21671 266113
rect 21699 266085 30485 266113
rect 30513 266085 30547 266113
rect 30575 266085 30609 266113
rect 30637 266085 30671 266113
rect 30699 266085 39485 266113
rect 39513 266085 39547 266113
rect 39575 266085 39609 266113
rect 39637 266085 39671 266113
rect 39699 266085 48485 266113
rect 48513 266085 48547 266113
rect 48575 266085 48609 266113
rect 48637 266085 48671 266113
rect 48699 266085 57485 266113
rect 57513 266085 57547 266113
rect 57575 266085 57609 266113
rect 57637 266085 57671 266113
rect 57699 266085 66485 266113
rect 66513 266085 66547 266113
rect 66575 266085 66609 266113
rect 66637 266085 66671 266113
rect 66699 266085 75485 266113
rect 75513 266085 75547 266113
rect 75575 266085 75609 266113
rect 75637 266085 75671 266113
rect 75699 266085 84485 266113
rect 84513 266085 84547 266113
rect 84575 266085 84609 266113
rect 84637 266085 84671 266113
rect 84699 266085 93485 266113
rect 93513 266085 93547 266113
rect 93575 266085 93609 266113
rect 93637 266085 93671 266113
rect 93699 266085 102485 266113
rect 102513 266085 102547 266113
rect 102575 266085 102609 266113
rect 102637 266085 102671 266113
rect 102699 266085 111485 266113
rect 111513 266085 111547 266113
rect 111575 266085 111609 266113
rect 111637 266085 111671 266113
rect 111699 266085 120485 266113
rect 120513 266085 120547 266113
rect 120575 266085 120609 266113
rect 120637 266085 120671 266113
rect 120699 266085 129485 266113
rect 129513 266085 129547 266113
rect 129575 266085 129609 266113
rect 129637 266085 129671 266113
rect 129699 266085 138485 266113
rect 138513 266085 138547 266113
rect 138575 266085 138609 266113
rect 138637 266085 138671 266113
rect 138699 266085 147485 266113
rect 147513 266085 147547 266113
rect 147575 266085 147609 266113
rect 147637 266085 147671 266113
rect 147699 266085 156485 266113
rect 156513 266085 156547 266113
rect 156575 266085 156609 266113
rect 156637 266085 156671 266113
rect 156699 266085 165485 266113
rect 165513 266085 165547 266113
rect 165575 266085 165609 266113
rect 165637 266085 165671 266113
rect 165699 266085 174485 266113
rect 174513 266085 174547 266113
rect 174575 266085 174609 266113
rect 174637 266085 174671 266113
rect 174699 266085 183485 266113
rect 183513 266085 183547 266113
rect 183575 266085 183609 266113
rect 183637 266085 183671 266113
rect 183699 266085 192485 266113
rect 192513 266085 192547 266113
rect 192575 266085 192609 266113
rect 192637 266085 192671 266113
rect 192699 266085 201485 266113
rect 201513 266085 201547 266113
rect 201575 266085 201609 266113
rect 201637 266085 201671 266113
rect 201699 266085 210485 266113
rect 210513 266085 210547 266113
rect 210575 266085 210609 266113
rect 210637 266085 210671 266113
rect 210699 266085 219485 266113
rect 219513 266085 219547 266113
rect 219575 266085 219609 266113
rect 219637 266085 219671 266113
rect 219699 266085 228485 266113
rect 228513 266085 228547 266113
rect 228575 266085 228609 266113
rect 228637 266085 228671 266113
rect 228699 266085 237485 266113
rect 237513 266085 237547 266113
rect 237575 266085 237609 266113
rect 237637 266085 237671 266113
rect 237699 266085 246485 266113
rect 246513 266085 246547 266113
rect 246575 266085 246609 266113
rect 246637 266085 246671 266113
rect 246699 266085 255485 266113
rect 255513 266085 255547 266113
rect 255575 266085 255609 266113
rect 255637 266085 255671 266113
rect 255699 266085 264485 266113
rect 264513 266085 264547 266113
rect 264575 266085 264609 266113
rect 264637 266085 264671 266113
rect 264699 266085 273485 266113
rect 273513 266085 273547 266113
rect 273575 266085 273609 266113
rect 273637 266085 273671 266113
rect 273699 266085 282485 266113
rect 282513 266085 282547 266113
rect 282575 266085 282609 266113
rect 282637 266085 282671 266113
rect 282699 266085 291485 266113
rect 291513 266085 291547 266113
rect 291575 266085 291609 266113
rect 291637 266085 291671 266113
rect 291699 266085 298728 266113
rect 298756 266085 298790 266113
rect 298818 266085 298852 266113
rect 298880 266085 298914 266113
rect 298942 266085 298990 266113
rect -958 266051 298990 266085
rect -958 266023 -910 266051
rect -882 266023 -848 266051
rect -820 266023 -786 266051
rect -758 266023 -724 266051
rect -696 266023 3485 266051
rect 3513 266023 3547 266051
rect 3575 266023 3609 266051
rect 3637 266023 3671 266051
rect 3699 266023 12485 266051
rect 12513 266023 12547 266051
rect 12575 266023 12609 266051
rect 12637 266023 12671 266051
rect 12699 266023 21485 266051
rect 21513 266023 21547 266051
rect 21575 266023 21609 266051
rect 21637 266023 21671 266051
rect 21699 266023 30485 266051
rect 30513 266023 30547 266051
rect 30575 266023 30609 266051
rect 30637 266023 30671 266051
rect 30699 266023 39485 266051
rect 39513 266023 39547 266051
rect 39575 266023 39609 266051
rect 39637 266023 39671 266051
rect 39699 266023 48485 266051
rect 48513 266023 48547 266051
rect 48575 266023 48609 266051
rect 48637 266023 48671 266051
rect 48699 266023 57485 266051
rect 57513 266023 57547 266051
rect 57575 266023 57609 266051
rect 57637 266023 57671 266051
rect 57699 266023 66485 266051
rect 66513 266023 66547 266051
rect 66575 266023 66609 266051
rect 66637 266023 66671 266051
rect 66699 266023 75485 266051
rect 75513 266023 75547 266051
rect 75575 266023 75609 266051
rect 75637 266023 75671 266051
rect 75699 266023 84485 266051
rect 84513 266023 84547 266051
rect 84575 266023 84609 266051
rect 84637 266023 84671 266051
rect 84699 266023 93485 266051
rect 93513 266023 93547 266051
rect 93575 266023 93609 266051
rect 93637 266023 93671 266051
rect 93699 266023 102485 266051
rect 102513 266023 102547 266051
rect 102575 266023 102609 266051
rect 102637 266023 102671 266051
rect 102699 266023 111485 266051
rect 111513 266023 111547 266051
rect 111575 266023 111609 266051
rect 111637 266023 111671 266051
rect 111699 266023 120485 266051
rect 120513 266023 120547 266051
rect 120575 266023 120609 266051
rect 120637 266023 120671 266051
rect 120699 266023 129485 266051
rect 129513 266023 129547 266051
rect 129575 266023 129609 266051
rect 129637 266023 129671 266051
rect 129699 266023 138485 266051
rect 138513 266023 138547 266051
rect 138575 266023 138609 266051
rect 138637 266023 138671 266051
rect 138699 266023 147485 266051
rect 147513 266023 147547 266051
rect 147575 266023 147609 266051
rect 147637 266023 147671 266051
rect 147699 266023 156485 266051
rect 156513 266023 156547 266051
rect 156575 266023 156609 266051
rect 156637 266023 156671 266051
rect 156699 266023 165485 266051
rect 165513 266023 165547 266051
rect 165575 266023 165609 266051
rect 165637 266023 165671 266051
rect 165699 266023 174485 266051
rect 174513 266023 174547 266051
rect 174575 266023 174609 266051
rect 174637 266023 174671 266051
rect 174699 266023 183485 266051
rect 183513 266023 183547 266051
rect 183575 266023 183609 266051
rect 183637 266023 183671 266051
rect 183699 266023 192485 266051
rect 192513 266023 192547 266051
rect 192575 266023 192609 266051
rect 192637 266023 192671 266051
rect 192699 266023 201485 266051
rect 201513 266023 201547 266051
rect 201575 266023 201609 266051
rect 201637 266023 201671 266051
rect 201699 266023 210485 266051
rect 210513 266023 210547 266051
rect 210575 266023 210609 266051
rect 210637 266023 210671 266051
rect 210699 266023 219485 266051
rect 219513 266023 219547 266051
rect 219575 266023 219609 266051
rect 219637 266023 219671 266051
rect 219699 266023 228485 266051
rect 228513 266023 228547 266051
rect 228575 266023 228609 266051
rect 228637 266023 228671 266051
rect 228699 266023 237485 266051
rect 237513 266023 237547 266051
rect 237575 266023 237609 266051
rect 237637 266023 237671 266051
rect 237699 266023 246485 266051
rect 246513 266023 246547 266051
rect 246575 266023 246609 266051
rect 246637 266023 246671 266051
rect 246699 266023 255485 266051
rect 255513 266023 255547 266051
rect 255575 266023 255609 266051
rect 255637 266023 255671 266051
rect 255699 266023 264485 266051
rect 264513 266023 264547 266051
rect 264575 266023 264609 266051
rect 264637 266023 264671 266051
rect 264699 266023 273485 266051
rect 273513 266023 273547 266051
rect 273575 266023 273609 266051
rect 273637 266023 273671 266051
rect 273699 266023 282485 266051
rect 282513 266023 282547 266051
rect 282575 266023 282609 266051
rect 282637 266023 282671 266051
rect 282699 266023 291485 266051
rect 291513 266023 291547 266051
rect 291575 266023 291609 266051
rect 291637 266023 291671 266051
rect 291699 266023 298728 266051
rect 298756 266023 298790 266051
rect 298818 266023 298852 266051
rect 298880 266023 298914 266051
rect 298942 266023 298990 266051
rect -958 265989 298990 266023
rect -958 265961 -910 265989
rect -882 265961 -848 265989
rect -820 265961 -786 265989
rect -758 265961 -724 265989
rect -696 265961 3485 265989
rect 3513 265961 3547 265989
rect 3575 265961 3609 265989
rect 3637 265961 3671 265989
rect 3699 265961 12485 265989
rect 12513 265961 12547 265989
rect 12575 265961 12609 265989
rect 12637 265961 12671 265989
rect 12699 265961 21485 265989
rect 21513 265961 21547 265989
rect 21575 265961 21609 265989
rect 21637 265961 21671 265989
rect 21699 265961 30485 265989
rect 30513 265961 30547 265989
rect 30575 265961 30609 265989
rect 30637 265961 30671 265989
rect 30699 265961 39485 265989
rect 39513 265961 39547 265989
rect 39575 265961 39609 265989
rect 39637 265961 39671 265989
rect 39699 265961 48485 265989
rect 48513 265961 48547 265989
rect 48575 265961 48609 265989
rect 48637 265961 48671 265989
rect 48699 265961 57485 265989
rect 57513 265961 57547 265989
rect 57575 265961 57609 265989
rect 57637 265961 57671 265989
rect 57699 265961 66485 265989
rect 66513 265961 66547 265989
rect 66575 265961 66609 265989
rect 66637 265961 66671 265989
rect 66699 265961 75485 265989
rect 75513 265961 75547 265989
rect 75575 265961 75609 265989
rect 75637 265961 75671 265989
rect 75699 265961 84485 265989
rect 84513 265961 84547 265989
rect 84575 265961 84609 265989
rect 84637 265961 84671 265989
rect 84699 265961 93485 265989
rect 93513 265961 93547 265989
rect 93575 265961 93609 265989
rect 93637 265961 93671 265989
rect 93699 265961 102485 265989
rect 102513 265961 102547 265989
rect 102575 265961 102609 265989
rect 102637 265961 102671 265989
rect 102699 265961 111485 265989
rect 111513 265961 111547 265989
rect 111575 265961 111609 265989
rect 111637 265961 111671 265989
rect 111699 265961 120485 265989
rect 120513 265961 120547 265989
rect 120575 265961 120609 265989
rect 120637 265961 120671 265989
rect 120699 265961 129485 265989
rect 129513 265961 129547 265989
rect 129575 265961 129609 265989
rect 129637 265961 129671 265989
rect 129699 265961 138485 265989
rect 138513 265961 138547 265989
rect 138575 265961 138609 265989
rect 138637 265961 138671 265989
rect 138699 265961 147485 265989
rect 147513 265961 147547 265989
rect 147575 265961 147609 265989
rect 147637 265961 147671 265989
rect 147699 265961 156485 265989
rect 156513 265961 156547 265989
rect 156575 265961 156609 265989
rect 156637 265961 156671 265989
rect 156699 265961 165485 265989
rect 165513 265961 165547 265989
rect 165575 265961 165609 265989
rect 165637 265961 165671 265989
rect 165699 265961 174485 265989
rect 174513 265961 174547 265989
rect 174575 265961 174609 265989
rect 174637 265961 174671 265989
rect 174699 265961 183485 265989
rect 183513 265961 183547 265989
rect 183575 265961 183609 265989
rect 183637 265961 183671 265989
rect 183699 265961 192485 265989
rect 192513 265961 192547 265989
rect 192575 265961 192609 265989
rect 192637 265961 192671 265989
rect 192699 265961 201485 265989
rect 201513 265961 201547 265989
rect 201575 265961 201609 265989
rect 201637 265961 201671 265989
rect 201699 265961 210485 265989
rect 210513 265961 210547 265989
rect 210575 265961 210609 265989
rect 210637 265961 210671 265989
rect 210699 265961 219485 265989
rect 219513 265961 219547 265989
rect 219575 265961 219609 265989
rect 219637 265961 219671 265989
rect 219699 265961 228485 265989
rect 228513 265961 228547 265989
rect 228575 265961 228609 265989
rect 228637 265961 228671 265989
rect 228699 265961 237485 265989
rect 237513 265961 237547 265989
rect 237575 265961 237609 265989
rect 237637 265961 237671 265989
rect 237699 265961 246485 265989
rect 246513 265961 246547 265989
rect 246575 265961 246609 265989
rect 246637 265961 246671 265989
rect 246699 265961 255485 265989
rect 255513 265961 255547 265989
rect 255575 265961 255609 265989
rect 255637 265961 255671 265989
rect 255699 265961 264485 265989
rect 264513 265961 264547 265989
rect 264575 265961 264609 265989
rect 264637 265961 264671 265989
rect 264699 265961 273485 265989
rect 273513 265961 273547 265989
rect 273575 265961 273609 265989
rect 273637 265961 273671 265989
rect 273699 265961 282485 265989
rect 282513 265961 282547 265989
rect 282575 265961 282609 265989
rect 282637 265961 282671 265989
rect 282699 265961 291485 265989
rect 291513 265961 291547 265989
rect 291575 265961 291609 265989
rect 291637 265961 291671 265989
rect 291699 265961 298728 265989
rect 298756 265961 298790 265989
rect 298818 265961 298852 265989
rect 298880 265961 298914 265989
rect 298942 265961 298990 265989
rect -958 265913 298990 265961
rect -958 263175 298990 263223
rect -958 263147 -430 263175
rect -402 263147 -368 263175
rect -340 263147 -306 263175
rect -278 263147 -244 263175
rect -216 263147 1625 263175
rect 1653 263147 1687 263175
rect 1715 263147 1749 263175
rect 1777 263147 1811 263175
rect 1839 263147 10625 263175
rect 10653 263147 10687 263175
rect 10715 263147 10749 263175
rect 10777 263147 10811 263175
rect 10839 263147 19625 263175
rect 19653 263147 19687 263175
rect 19715 263147 19749 263175
rect 19777 263147 19811 263175
rect 19839 263147 28625 263175
rect 28653 263147 28687 263175
rect 28715 263147 28749 263175
rect 28777 263147 28811 263175
rect 28839 263147 37625 263175
rect 37653 263147 37687 263175
rect 37715 263147 37749 263175
rect 37777 263147 37811 263175
rect 37839 263147 46625 263175
rect 46653 263147 46687 263175
rect 46715 263147 46749 263175
rect 46777 263147 46811 263175
rect 46839 263147 55625 263175
rect 55653 263147 55687 263175
rect 55715 263147 55749 263175
rect 55777 263147 55811 263175
rect 55839 263147 64625 263175
rect 64653 263147 64687 263175
rect 64715 263147 64749 263175
rect 64777 263147 64811 263175
rect 64839 263147 73625 263175
rect 73653 263147 73687 263175
rect 73715 263147 73749 263175
rect 73777 263147 73811 263175
rect 73839 263147 82625 263175
rect 82653 263147 82687 263175
rect 82715 263147 82749 263175
rect 82777 263147 82811 263175
rect 82839 263147 91625 263175
rect 91653 263147 91687 263175
rect 91715 263147 91749 263175
rect 91777 263147 91811 263175
rect 91839 263147 100625 263175
rect 100653 263147 100687 263175
rect 100715 263147 100749 263175
rect 100777 263147 100811 263175
rect 100839 263147 109625 263175
rect 109653 263147 109687 263175
rect 109715 263147 109749 263175
rect 109777 263147 109811 263175
rect 109839 263147 118625 263175
rect 118653 263147 118687 263175
rect 118715 263147 118749 263175
rect 118777 263147 118811 263175
rect 118839 263147 127625 263175
rect 127653 263147 127687 263175
rect 127715 263147 127749 263175
rect 127777 263147 127811 263175
rect 127839 263147 136625 263175
rect 136653 263147 136687 263175
rect 136715 263147 136749 263175
rect 136777 263147 136811 263175
rect 136839 263147 145625 263175
rect 145653 263147 145687 263175
rect 145715 263147 145749 263175
rect 145777 263147 145811 263175
rect 145839 263147 154625 263175
rect 154653 263147 154687 263175
rect 154715 263147 154749 263175
rect 154777 263147 154811 263175
rect 154839 263147 163625 263175
rect 163653 263147 163687 263175
rect 163715 263147 163749 263175
rect 163777 263147 163811 263175
rect 163839 263147 172625 263175
rect 172653 263147 172687 263175
rect 172715 263147 172749 263175
rect 172777 263147 172811 263175
rect 172839 263147 181625 263175
rect 181653 263147 181687 263175
rect 181715 263147 181749 263175
rect 181777 263147 181811 263175
rect 181839 263147 190625 263175
rect 190653 263147 190687 263175
rect 190715 263147 190749 263175
rect 190777 263147 190811 263175
rect 190839 263147 199625 263175
rect 199653 263147 199687 263175
rect 199715 263147 199749 263175
rect 199777 263147 199811 263175
rect 199839 263147 208625 263175
rect 208653 263147 208687 263175
rect 208715 263147 208749 263175
rect 208777 263147 208811 263175
rect 208839 263147 217625 263175
rect 217653 263147 217687 263175
rect 217715 263147 217749 263175
rect 217777 263147 217811 263175
rect 217839 263147 226625 263175
rect 226653 263147 226687 263175
rect 226715 263147 226749 263175
rect 226777 263147 226811 263175
rect 226839 263147 235625 263175
rect 235653 263147 235687 263175
rect 235715 263147 235749 263175
rect 235777 263147 235811 263175
rect 235839 263147 244625 263175
rect 244653 263147 244687 263175
rect 244715 263147 244749 263175
rect 244777 263147 244811 263175
rect 244839 263147 253625 263175
rect 253653 263147 253687 263175
rect 253715 263147 253749 263175
rect 253777 263147 253811 263175
rect 253839 263147 262625 263175
rect 262653 263147 262687 263175
rect 262715 263147 262749 263175
rect 262777 263147 262811 263175
rect 262839 263147 271625 263175
rect 271653 263147 271687 263175
rect 271715 263147 271749 263175
rect 271777 263147 271811 263175
rect 271839 263147 280625 263175
rect 280653 263147 280687 263175
rect 280715 263147 280749 263175
rect 280777 263147 280811 263175
rect 280839 263147 289625 263175
rect 289653 263147 289687 263175
rect 289715 263147 289749 263175
rect 289777 263147 289811 263175
rect 289839 263147 298248 263175
rect 298276 263147 298310 263175
rect 298338 263147 298372 263175
rect 298400 263147 298434 263175
rect 298462 263147 298990 263175
rect -958 263113 298990 263147
rect -958 263085 -430 263113
rect -402 263085 -368 263113
rect -340 263085 -306 263113
rect -278 263085 -244 263113
rect -216 263085 1625 263113
rect 1653 263085 1687 263113
rect 1715 263085 1749 263113
rect 1777 263085 1811 263113
rect 1839 263085 10625 263113
rect 10653 263085 10687 263113
rect 10715 263085 10749 263113
rect 10777 263085 10811 263113
rect 10839 263085 19625 263113
rect 19653 263085 19687 263113
rect 19715 263085 19749 263113
rect 19777 263085 19811 263113
rect 19839 263085 28625 263113
rect 28653 263085 28687 263113
rect 28715 263085 28749 263113
rect 28777 263085 28811 263113
rect 28839 263085 37625 263113
rect 37653 263085 37687 263113
rect 37715 263085 37749 263113
rect 37777 263085 37811 263113
rect 37839 263085 46625 263113
rect 46653 263085 46687 263113
rect 46715 263085 46749 263113
rect 46777 263085 46811 263113
rect 46839 263085 55625 263113
rect 55653 263085 55687 263113
rect 55715 263085 55749 263113
rect 55777 263085 55811 263113
rect 55839 263085 64625 263113
rect 64653 263085 64687 263113
rect 64715 263085 64749 263113
rect 64777 263085 64811 263113
rect 64839 263085 73625 263113
rect 73653 263085 73687 263113
rect 73715 263085 73749 263113
rect 73777 263085 73811 263113
rect 73839 263085 82625 263113
rect 82653 263085 82687 263113
rect 82715 263085 82749 263113
rect 82777 263085 82811 263113
rect 82839 263085 91625 263113
rect 91653 263085 91687 263113
rect 91715 263085 91749 263113
rect 91777 263085 91811 263113
rect 91839 263085 100625 263113
rect 100653 263085 100687 263113
rect 100715 263085 100749 263113
rect 100777 263085 100811 263113
rect 100839 263085 109625 263113
rect 109653 263085 109687 263113
rect 109715 263085 109749 263113
rect 109777 263085 109811 263113
rect 109839 263085 118625 263113
rect 118653 263085 118687 263113
rect 118715 263085 118749 263113
rect 118777 263085 118811 263113
rect 118839 263085 127625 263113
rect 127653 263085 127687 263113
rect 127715 263085 127749 263113
rect 127777 263085 127811 263113
rect 127839 263085 136625 263113
rect 136653 263085 136687 263113
rect 136715 263085 136749 263113
rect 136777 263085 136811 263113
rect 136839 263085 145625 263113
rect 145653 263085 145687 263113
rect 145715 263085 145749 263113
rect 145777 263085 145811 263113
rect 145839 263085 154625 263113
rect 154653 263085 154687 263113
rect 154715 263085 154749 263113
rect 154777 263085 154811 263113
rect 154839 263085 163625 263113
rect 163653 263085 163687 263113
rect 163715 263085 163749 263113
rect 163777 263085 163811 263113
rect 163839 263085 172625 263113
rect 172653 263085 172687 263113
rect 172715 263085 172749 263113
rect 172777 263085 172811 263113
rect 172839 263085 181625 263113
rect 181653 263085 181687 263113
rect 181715 263085 181749 263113
rect 181777 263085 181811 263113
rect 181839 263085 190625 263113
rect 190653 263085 190687 263113
rect 190715 263085 190749 263113
rect 190777 263085 190811 263113
rect 190839 263085 199625 263113
rect 199653 263085 199687 263113
rect 199715 263085 199749 263113
rect 199777 263085 199811 263113
rect 199839 263085 208625 263113
rect 208653 263085 208687 263113
rect 208715 263085 208749 263113
rect 208777 263085 208811 263113
rect 208839 263085 217625 263113
rect 217653 263085 217687 263113
rect 217715 263085 217749 263113
rect 217777 263085 217811 263113
rect 217839 263085 226625 263113
rect 226653 263085 226687 263113
rect 226715 263085 226749 263113
rect 226777 263085 226811 263113
rect 226839 263085 235625 263113
rect 235653 263085 235687 263113
rect 235715 263085 235749 263113
rect 235777 263085 235811 263113
rect 235839 263085 244625 263113
rect 244653 263085 244687 263113
rect 244715 263085 244749 263113
rect 244777 263085 244811 263113
rect 244839 263085 253625 263113
rect 253653 263085 253687 263113
rect 253715 263085 253749 263113
rect 253777 263085 253811 263113
rect 253839 263085 262625 263113
rect 262653 263085 262687 263113
rect 262715 263085 262749 263113
rect 262777 263085 262811 263113
rect 262839 263085 271625 263113
rect 271653 263085 271687 263113
rect 271715 263085 271749 263113
rect 271777 263085 271811 263113
rect 271839 263085 280625 263113
rect 280653 263085 280687 263113
rect 280715 263085 280749 263113
rect 280777 263085 280811 263113
rect 280839 263085 289625 263113
rect 289653 263085 289687 263113
rect 289715 263085 289749 263113
rect 289777 263085 289811 263113
rect 289839 263085 298248 263113
rect 298276 263085 298310 263113
rect 298338 263085 298372 263113
rect 298400 263085 298434 263113
rect 298462 263085 298990 263113
rect -958 263051 298990 263085
rect -958 263023 -430 263051
rect -402 263023 -368 263051
rect -340 263023 -306 263051
rect -278 263023 -244 263051
rect -216 263023 1625 263051
rect 1653 263023 1687 263051
rect 1715 263023 1749 263051
rect 1777 263023 1811 263051
rect 1839 263023 10625 263051
rect 10653 263023 10687 263051
rect 10715 263023 10749 263051
rect 10777 263023 10811 263051
rect 10839 263023 19625 263051
rect 19653 263023 19687 263051
rect 19715 263023 19749 263051
rect 19777 263023 19811 263051
rect 19839 263023 28625 263051
rect 28653 263023 28687 263051
rect 28715 263023 28749 263051
rect 28777 263023 28811 263051
rect 28839 263023 37625 263051
rect 37653 263023 37687 263051
rect 37715 263023 37749 263051
rect 37777 263023 37811 263051
rect 37839 263023 46625 263051
rect 46653 263023 46687 263051
rect 46715 263023 46749 263051
rect 46777 263023 46811 263051
rect 46839 263023 55625 263051
rect 55653 263023 55687 263051
rect 55715 263023 55749 263051
rect 55777 263023 55811 263051
rect 55839 263023 64625 263051
rect 64653 263023 64687 263051
rect 64715 263023 64749 263051
rect 64777 263023 64811 263051
rect 64839 263023 73625 263051
rect 73653 263023 73687 263051
rect 73715 263023 73749 263051
rect 73777 263023 73811 263051
rect 73839 263023 82625 263051
rect 82653 263023 82687 263051
rect 82715 263023 82749 263051
rect 82777 263023 82811 263051
rect 82839 263023 91625 263051
rect 91653 263023 91687 263051
rect 91715 263023 91749 263051
rect 91777 263023 91811 263051
rect 91839 263023 100625 263051
rect 100653 263023 100687 263051
rect 100715 263023 100749 263051
rect 100777 263023 100811 263051
rect 100839 263023 109625 263051
rect 109653 263023 109687 263051
rect 109715 263023 109749 263051
rect 109777 263023 109811 263051
rect 109839 263023 118625 263051
rect 118653 263023 118687 263051
rect 118715 263023 118749 263051
rect 118777 263023 118811 263051
rect 118839 263023 127625 263051
rect 127653 263023 127687 263051
rect 127715 263023 127749 263051
rect 127777 263023 127811 263051
rect 127839 263023 136625 263051
rect 136653 263023 136687 263051
rect 136715 263023 136749 263051
rect 136777 263023 136811 263051
rect 136839 263023 145625 263051
rect 145653 263023 145687 263051
rect 145715 263023 145749 263051
rect 145777 263023 145811 263051
rect 145839 263023 154625 263051
rect 154653 263023 154687 263051
rect 154715 263023 154749 263051
rect 154777 263023 154811 263051
rect 154839 263023 163625 263051
rect 163653 263023 163687 263051
rect 163715 263023 163749 263051
rect 163777 263023 163811 263051
rect 163839 263023 172625 263051
rect 172653 263023 172687 263051
rect 172715 263023 172749 263051
rect 172777 263023 172811 263051
rect 172839 263023 181625 263051
rect 181653 263023 181687 263051
rect 181715 263023 181749 263051
rect 181777 263023 181811 263051
rect 181839 263023 190625 263051
rect 190653 263023 190687 263051
rect 190715 263023 190749 263051
rect 190777 263023 190811 263051
rect 190839 263023 199625 263051
rect 199653 263023 199687 263051
rect 199715 263023 199749 263051
rect 199777 263023 199811 263051
rect 199839 263023 208625 263051
rect 208653 263023 208687 263051
rect 208715 263023 208749 263051
rect 208777 263023 208811 263051
rect 208839 263023 217625 263051
rect 217653 263023 217687 263051
rect 217715 263023 217749 263051
rect 217777 263023 217811 263051
rect 217839 263023 226625 263051
rect 226653 263023 226687 263051
rect 226715 263023 226749 263051
rect 226777 263023 226811 263051
rect 226839 263023 235625 263051
rect 235653 263023 235687 263051
rect 235715 263023 235749 263051
rect 235777 263023 235811 263051
rect 235839 263023 244625 263051
rect 244653 263023 244687 263051
rect 244715 263023 244749 263051
rect 244777 263023 244811 263051
rect 244839 263023 253625 263051
rect 253653 263023 253687 263051
rect 253715 263023 253749 263051
rect 253777 263023 253811 263051
rect 253839 263023 262625 263051
rect 262653 263023 262687 263051
rect 262715 263023 262749 263051
rect 262777 263023 262811 263051
rect 262839 263023 271625 263051
rect 271653 263023 271687 263051
rect 271715 263023 271749 263051
rect 271777 263023 271811 263051
rect 271839 263023 280625 263051
rect 280653 263023 280687 263051
rect 280715 263023 280749 263051
rect 280777 263023 280811 263051
rect 280839 263023 289625 263051
rect 289653 263023 289687 263051
rect 289715 263023 289749 263051
rect 289777 263023 289811 263051
rect 289839 263023 298248 263051
rect 298276 263023 298310 263051
rect 298338 263023 298372 263051
rect 298400 263023 298434 263051
rect 298462 263023 298990 263051
rect -958 262989 298990 263023
rect -958 262961 -430 262989
rect -402 262961 -368 262989
rect -340 262961 -306 262989
rect -278 262961 -244 262989
rect -216 262961 1625 262989
rect 1653 262961 1687 262989
rect 1715 262961 1749 262989
rect 1777 262961 1811 262989
rect 1839 262961 10625 262989
rect 10653 262961 10687 262989
rect 10715 262961 10749 262989
rect 10777 262961 10811 262989
rect 10839 262961 19625 262989
rect 19653 262961 19687 262989
rect 19715 262961 19749 262989
rect 19777 262961 19811 262989
rect 19839 262961 28625 262989
rect 28653 262961 28687 262989
rect 28715 262961 28749 262989
rect 28777 262961 28811 262989
rect 28839 262961 37625 262989
rect 37653 262961 37687 262989
rect 37715 262961 37749 262989
rect 37777 262961 37811 262989
rect 37839 262961 46625 262989
rect 46653 262961 46687 262989
rect 46715 262961 46749 262989
rect 46777 262961 46811 262989
rect 46839 262961 55625 262989
rect 55653 262961 55687 262989
rect 55715 262961 55749 262989
rect 55777 262961 55811 262989
rect 55839 262961 64625 262989
rect 64653 262961 64687 262989
rect 64715 262961 64749 262989
rect 64777 262961 64811 262989
rect 64839 262961 73625 262989
rect 73653 262961 73687 262989
rect 73715 262961 73749 262989
rect 73777 262961 73811 262989
rect 73839 262961 82625 262989
rect 82653 262961 82687 262989
rect 82715 262961 82749 262989
rect 82777 262961 82811 262989
rect 82839 262961 91625 262989
rect 91653 262961 91687 262989
rect 91715 262961 91749 262989
rect 91777 262961 91811 262989
rect 91839 262961 100625 262989
rect 100653 262961 100687 262989
rect 100715 262961 100749 262989
rect 100777 262961 100811 262989
rect 100839 262961 109625 262989
rect 109653 262961 109687 262989
rect 109715 262961 109749 262989
rect 109777 262961 109811 262989
rect 109839 262961 118625 262989
rect 118653 262961 118687 262989
rect 118715 262961 118749 262989
rect 118777 262961 118811 262989
rect 118839 262961 127625 262989
rect 127653 262961 127687 262989
rect 127715 262961 127749 262989
rect 127777 262961 127811 262989
rect 127839 262961 136625 262989
rect 136653 262961 136687 262989
rect 136715 262961 136749 262989
rect 136777 262961 136811 262989
rect 136839 262961 145625 262989
rect 145653 262961 145687 262989
rect 145715 262961 145749 262989
rect 145777 262961 145811 262989
rect 145839 262961 154625 262989
rect 154653 262961 154687 262989
rect 154715 262961 154749 262989
rect 154777 262961 154811 262989
rect 154839 262961 163625 262989
rect 163653 262961 163687 262989
rect 163715 262961 163749 262989
rect 163777 262961 163811 262989
rect 163839 262961 172625 262989
rect 172653 262961 172687 262989
rect 172715 262961 172749 262989
rect 172777 262961 172811 262989
rect 172839 262961 181625 262989
rect 181653 262961 181687 262989
rect 181715 262961 181749 262989
rect 181777 262961 181811 262989
rect 181839 262961 190625 262989
rect 190653 262961 190687 262989
rect 190715 262961 190749 262989
rect 190777 262961 190811 262989
rect 190839 262961 199625 262989
rect 199653 262961 199687 262989
rect 199715 262961 199749 262989
rect 199777 262961 199811 262989
rect 199839 262961 208625 262989
rect 208653 262961 208687 262989
rect 208715 262961 208749 262989
rect 208777 262961 208811 262989
rect 208839 262961 217625 262989
rect 217653 262961 217687 262989
rect 217715 262961 217749 262989
rect 217777 262961 217811 262989
rect 217839 262961 226625 262989
rect 226653 262961 226687 262989
rect 226715 262961 226749 262989
rect 226777 262961 226811 262989
rect 226839 262961 235625 262989
rect 235653 262961 235687 262989
rect 235715 262961 235749 262989
rect 235777 262961 235811 262989
rect 235839 262961 244625 262989
rect 244653 262961 244687 262989
rect 244715 262961 244749 262989
rect 244777 262961 244811 262989
rect 244839 262961 253625 262989
rect 253653 262961 253687 262989
rect 253715 262961 253749 262989
rect 253777 262961 253811 262989
rect 253839 262961 262625 262989
rect 262653 262961 262687 262989
rect 262715 262961 262749 262989
rect 262777 262961 262811 262989
rect 262839 262961 271625 262989
rect 271653 262961 271687 262989
rect 271715 262961 271749 262989
rect 271777 262961 271811 262989
rect 271839 262961 280625 262989
rect 280653 262961 280687 262989
rect 280715 262961 280749 262989
rect 280777 262961 280811 262989
rect 280839 262961 289625 262989
rect 289653 262961 289687 262989
rect 289715 262961 289749 262989
rect 289777 262961 289811 262989
rect 289839 262961 298248 262989
rect 298276 262961 298310 262989
rect 298338 262961 298372 262989
rect 298400 262961 298434 262989
rect 298462 262961 298990 262989
rect -958 262913 298990 262961
rect -958 257175 298990 257223
rect -958 257147 -910 257175
rect -882 257147 -848 257175
rect -820 257147 -786 257175
rect -758 257147 -724 257175
rect -696 257147 3485 257175
rect 3513 257147 3547 257175
rect 3575 257147 3609 257175
rect 3637 257147 3671 257175
rect 3699 257147 12485 257175
rect 12513 257147 12547 257175
rect 12575 257147 12609 257175
rect 12637 257147 12671 257175
rect 12699 257147 21485 257175
rect 21513 257147 21547 257175
rect 21575 257147 21609 257175
rect 21637 257147 21671 257175
rect 21699 257147 30485 257175
rect 30513 257147 30547 257175
rect 30575 257147 30609 257175
rect 30637 257147 30671 257175
rect 30699 257147 39485 257175
rect 39513 257147 39547 257175
rect 39575 257147 39609 257175
rect 39637 257147 39671 257175
rect 39699 257147 48485 257175
rect 48513 257147 48547 257175
rect 48575 257147 48609 257175
rect 48637 257147 48671 257175
rect 48699 257147 59939 257175
rect 59967 257147 60001 257175
rect 60029 257147 75299 257175
rect 75327 257147 75361 257175
rect 75389 257147 90659 257175
rect 90687 257147 90721 257175
rect 90749 257147 106019 257175
rect 106047 257147 106081 257175
rect 106109 257147 121379 257175
rect 121407 257147 121441 257175
rect 121469 257147 136739 257175
rect 136767 257147 136801 257175
rect 136829 257147 156485 257175
rect 156513 257147 156547 257175
rect 156575 257147 156609 257175
rect 156637 257147 156671 257175
rect 156699 257147 165485 257175
rect 165513 257147 165547 257175
rect 165575 257147 165609 257175
rect 165637 257147 165671 257175
rect 165699 257147 174485 257175
rect 174513 257147 174547 257175
rect 174575 257147 174609 257175
rect 174637 257147 174671 257175
rect 174699 257147 183485 257175
rect 183513 257147 183547 257175
rect 183575 257147 183609 257175
rect 183637 257147 183671 257175
rect 183699 257147 192485 257175
rect 192513 257147 192547 257175
rect 192575 257147 192609 257175
rect 192637 257147 192671 257175
rect 192699 257147 201485 257175
rect 201513 257147 201547 257175
rect 201575 257147 201609 257175
rect 201637 257147 201671 257175
rect 201699 257147 210485 257175
rect 210513 257147 210547 257175
rect 210575 257147 210609 257175
rect 210637 257147 210671 257175
rect 210699 257147 219485 257175
rect 219513 257147 219547 257175
rect 219575 257147 219609 257175
rect 219637 257147 219671 257175
rect 219699 257147 228485 257175
rect 228513 257147 228547 257175
rect 228575 257147 228609 257175
rect 228637 257147 228671 257175
rect 228699 257147 237485 257175
rect 237513 257147 237547 257175
rect 237575 257147 237609 257175
rect 237637 257147 237671 257175
rect 237699 257147 246485 257175
rect 246513 257147 246547 257175
rect 246575 257147 246609 257175
rect 246637 257147 246671 257175
rect 246699 257147 255485 257175
rect 255513 257147 255547 257175
rect 255575 257147 255609 257175
rect 255637 257147 255671 257175
rect 255699 257147 264485 257175
rect 264513 257147 264547 257175
rect 264575 257147 264609 257175
rect 264637 257147 264671 257175
rect 264699 257147 273485 257175
rect 273513 257147 273547 257175
rect 273575 257147 273609 257175
rect 273637 257147 273671 257175
rect 273699 257147 282485 257175
rect 282513 257147 282547 257175
rect 282575 257147 282609 257175
rect 282637 257147 282671 257175
rect 282699 257147 291485 257175
rect 291513 257147 291547 257175
rect 291575 257147 291609 257175
rect 291637 257147 291671 257175
rect 291699 257147 298728 257175
rect 298756 257147 298790 257175
rect 298818 257147 298852 257175
rect 298880 257147 298914 257175
rect 298942 257147 298990 257175
rect -958 257113 298990 257147
rect -958 257085 -910 257113
rect -882 257085 -848 257113
rect -820 257085 -786 257113
rect -758 257085 -724 257113
rect -696 257085 3485 257113
rect 3513 257085 3547 257113
rect 3575 257085 3609 257113
rect 3637 257085 3671 257113
rect 3699 257085 12485 257113
rect 12513 257085 12547 257113
rect 12575 257085 12609 257113
rect 12637 257085 12671 257113
rect 12699 257085 21485 257113
rect 21513 257085 21547 257113
rect 21575 257085 21609 257113
rect 21637 257085 21671 257113
rect 21699 257085 30485 257113
rect 30513 257085 30547 257113
rect 30575 257085 30609 257113
rect 30637 257085 30671 257113
rect 30699 257085 39485 257113
rect 39513 257085 39547 257113
rect 39575 257085 39609 257113
rect 39637 257085 39671 257113
rect 39699 257085 48485 257113
rect 48513 257085 48547 257113
rect 48575 257085 48609 257113
rect 48637 257085 48671 257113
rect 48699 257085 59939 257113
rect 59967 257085 60001 257113
rect 60029 257085 75299 257113
rect 75327 257085 75361 257113
rect 75389 257085 90659 257113
rect 90687 257085 90721 257113
rect 90749 257085 106019 257113
rect 106047 257085 106081 257113
rect 106109 257085 121379 257113
rect 121407 257085 121441 257113
rect 121469 257085 136739 257113
rect 136767 257085 136801 257113
rect 136829 257085 156485 257113
rect 156513 257085 156547 257113
rect 156575 257085 156609 257113
rect 156637 257085 156671 257113
rect 156699 257085 165485 257113
rect 165513 257085 165547 257113
rect 165575 257085 165609 257113
rect 165637 257085 165671 257113
rect 165699 257085 174485 257113
rect 174513 257085 174547 257113
rect 174575 257085 174609 257113
rect 174637 257085 174671 257113
rect 174699 257085 183485 257113
rect 183513 257085 183547 257113
rect 183575 257085 183609 257113
rect 183637 257085 183671 257113
rect 183699 257085 192485 257113
rect 192513 257085 192547 257113
rect 192575 257085 192609 257113
rect 192637 257085 192671 257113
rect 192699 257085 201485 257113
rect 201513 257085 201547 257113
rect 201575 257085 201609 257113
rect 201637 257085 201671 257113
rect 201699 257085 210485 257113
rect 210513 257085 210547 257113
rect 210575 257085 210609 257113
rect 210637 257085 210671 257113
rect 210699 257085 219485 257113
rect 219513 257085 219547 257113
rect 219575 257085 219609 257113
rect 219637 257085 219671 257113
rect 219699 257085 228485 257113
rect 228513 257085 228547 257113
rect 228575 257085 228609 257113
rect 228637 257085 228671 257113
rect 228699 257085 237485 257113
rect 237513 257085 237547 257113
rect 237575 257085 237609 257113
rect 237637 257085 237671 257113
rect 237699 257085 246485 257113
rect 246513 257085 246547 257113
rect 246575 257085 246609 257113
rect 246637 257085 246671 257113
rect 246699 257085 255485 257113
rect 255513 257085 255547 257113
rect 255575 257085 255609 257113
rect 255637 257085 255671 257113
rect 255699 257085 264485 257113
rect 264513 257085 264547 257113
rect 264575 257085 264609 257113
rect 264637 257085 264671 257113
rect 264699 257085 273485 257113
rect 273513 257085 273547 257113
rect 273575 257085 273609 257113
rect 273637 257085 273671 257113
rect 273699 257085 282485 257113
rect 282513 257085 282547 257113
rect 282575 257085 282609 257113
rect 282637 257085 282671 257113
rect 282699 257085 291485 257113
rect 291513 257085 291547 257113
rect 291575 257085 291609 257113
rect 291637 257085 291671 257113
rect 291699 257085 298728 257113
rect 298756 257085 298790 257113
rect 298818 257085 298852 257113
rect 298880 257085 298914 257113
rect 298942 257085 298990 257113
rect -958 257051 298990 257085
rect -958 257023 -910 257051
rect -882 257023 -848 257051
rect -820 257023 -786 257051
rect -758 257023 -724 257051
rect -696 257023 3485 257051
rect 3513 257023 3547 257051
rect 3575 257023 3609 257051
rect 3637 257023 3671 257051
rect 3699 257023 12485 257051
rect 12513 257023 12547 257051
rect 12575 257023 12609 257051
rect 12637 257023 12671 257051
rect 12699 257023 21485 257051
rect 21513 257023 21547 257051
rect 21575 257023 21609 257051
rect 21637 257023 21671 257051
rect 21699 257023 30485 257051
rect 30513 257023 30547 257051
rect 30575 257023 30609 257051
rect 30637 257023 30671 257051
rect 30699 257023 39485 257051
rect 39513 257023 39547 257051
rect 39575 257023 39609 257051
rect 39637 257023 39671 257051
rect 39699 257023 48485 257051
rect 48513 257023 48547 257051
rect 48575 257023 48609 257051
rect 48637 257023 48671 257051
rect 48699 257023 59939 257051
rect 59967 257023 60001 257051
rect 60029 257023 75299 257051
rect 75327 257023 75361 257051
rect 75389 257023 90659 257051
rect 90687 257023 90721 257051
rect 90749 257023 106019 257051
rect 106047 257023 106081 257051
rect 106109 257023 121379 257051
rect 121407 257023 121441 257051
rect 121469 257023 136739 257051
rect 136767 257023 136801 257051
rect 136829 257023 156485 257051
rect 156513 257023 156547 257051
rect 156575 257023 156609 257051
rect 156637 257023 156671 257051
rect 156699 257023 165485 257051
rect 165513 257023 165547 257051
rect 165575 257023 165609 257051
rect 165637 257023 165671 257051
rect 165699 257023 174485 257051
rect 174513 257023 174547 257051
rect 174575 257023 174609 257051
rect 174637 257023 174671 257051
rect 174699 257023 183485 257051
rect 183513 257023 183547 257051
rect 183575 257023 183609 257051
rect 183637 257023 183671 257051
rect 183699 257023 192485 257051
rect 192513 257023 192547 257051
rect 192575 257023 192609 257051
rect 192637 257023 192671 257051
rect 192699 257023 201485 257051
rect 201513 257023 201547 257051
rect 201575 257023 201609 257051
rect 201637 257023 201671 257051
rect 201699 257023 210485 257051
rect 210513 257023 210547 257051
rect 210575 257023 210609 257051
rect 210637 257023 210671 257051
rect 210699 257023 219485 257051
rect 219513 257023 219547 257051
rect 219575 257023 219609 257051
rect 219637 257023 219671 257051
rect 219699 257023 228485 257051
rect 228513 257023 228547 257051
rect 228575 257023 228609 257051
rect 228637 257023 228671 257051
rect 228699 257023 237485 257051
rect 237513 257023 237547 257051
rect 237575 257023 237609 257051
rect 237637 257023 237671 257051
rect 237699 257023 246485 257051
rect 246513 257023 246547 257051
rect 246575 257023 246609 257051
rect 246637 257023 246671 257051
rect 246699 257023 255485 257051
rect 255513 257023 255547 257051
rect 255575 257023 255609 257051
rect 255637 257023 255671 257051
rect 255699 257023 264485 257051
rect 264513 257023 264547 257051
rect 264575 257023 264609 257051
rect 264637 257023 264671 257051
rect 264699 257023 273485 257051
rect 273513 257023 273547 257051
rect 273575 257023 273609 257051
rect 273637 257023 273671 257051
rect 273699 257023 282485 257051
rect 282513 257023 282547 257051
rect 282575 257023 282609 257051
rect 282637 257023 282671 257051
rect 282699 257023 291485 257051
rect 291513 257023 291547 257051
rect 291575 257023 291609 257051
rect 291637 257023 291671 257051
rect 291699 257023 298728 257051
rect 298756 257023 298790 257051
rect 298818 257023 298852 257051
rect 298880 257023 298914 257051
rect 298942 257023 298990 257051
rect -958 256989 298990 257023
rect -958 256961 -910 256989
rect -882 256961 -848 256989
rect -820 256961 -786 256989
rect -758 256961 -724 256989
rect -696 256961 3485 256989
rect 3513 256961 3547 256989
rect 3575 256961 3609 256989
rect 3637 256961 3671 256989
rect 3699 256961 12485 256989
rect 12513 256961 12547 256989
rect 12575 256961 12609 256989
rect 12637 256961 12671 256989
rect 12699 256961 21485 256989
rect 21513 256961 21547 256989
rect 21575 256961 21609 256989
rect 21637 256961 21671 256989
rect 21699 256961 30485 256989
rect 30513 256961 30547 256989
rect 30575 256961 30609 256989
rect 30637 256961 30671 256989
rect 30699 256961 39485 256989
rect 39513 256961 39547 256989
rect 39575 256961 39609 256989
rect 39637 256961 39671 256989
rect 39699 256961 48485 256989
rect 48513 256961 48547 256989
rect 48575 256961 48609 256989
rect 48637 256961 48671 256989
rect 48699 256961 59939 256989
rect 59967 256961 60001 256989
rect 60029 256961 75299 256989
rect 75327 256961 75361 256989
rect 75389 256961 90659 256989
rect 90687 256961 90721 256989
rect 90749 256961 106019 256989
rect 106047 256961 106081 256989
rect 106109 256961 121379 256989
rect 121407 256961 121441 256989
rect 121469 256961 136739 256989
rect 136767 256961 136801 256989
rect 136829 256961 156485 256989
rect 156513 256961 156547 256989
rect 156575 256961 156609 256989
rect 156637 256961 156671 256989
rect 156699 256961 165485 256989
rect 165513 256961 165547 256989
rect 165575 256961 165609 256989
rect 165637 256961 165671 256989
rect 165699 256961 174485 256989
rect 174513 256961 174547 256989
rect 174575 256961 174609 256989
rect 174637 256961 174671 256989
rect 174699 256961 183485 256989
rect 183513 256961 183547 256989
rect 183575 256961 183609 256989
rect 183637 256961 183671 256989
rect 183699 256961 192485 256989
rect 192513 256961 192547 256989
rect 192575 256961 192609 256989
rect 192637 256961 192671 256989
rect 192699 256961 201485 256989
rect 201513 256961 201547 256989
rect 201575 256961 201609 256989
rect 201637 256961 201671 256989
rect 201699 256961 210485 256989
rect 210513 256961 210547 256989
rect 210575 256961 210609 256989
rect 210637 256961 210671 256989
rect 210699 256961 219485 256989
rect 219513 256961 219547 256989
rect 219575 256961 219609 256989
rect 219637 256961 219671 256989
rect 219699 256961 228485 256989
rect 228513 256961 228547 256989
rect 228575 256961 228609 256989
rect 228637 256961 228671 256989
rect 228699 256961 237485 256989
rect 237513 256961 237547 256989
rect 237575 256961 237609 256989
rect 237637 256961 237671 256989
rect 237699 256961 246485 256989
rect 246513 256961 246547 256989
rect 246575 256961 246609 256989
rect 246637 256961 246671 256989
rect 246699 256961 255485 256989
rect 255513 256961 255547 256989
rect 255575 256961 255609 256989
rect 255637 256961 255671 256989
rect 255699 256961 264485 256989
rect 264513 256961 264547 256989
rect 264575 256961 264609 256989
rect 264637 256961 264671 256989
rect 264699 256961 273485 256989
rect 273513 256961 273547 256989
rect 273575 256961 273609 256989
rect 273637 256961 273671 256989
rect 273699 256961 282485 256989
rect 282513 256961 282547 256989
rect 282575 256961 282609 256989
rect 282637 256961 282671 256989
rect 282699 256961 291485 256989
rect 291513 256961 291547 256989
rect 291575 256961 291609 256989
rect 291637 256961 291671 256989
rect 291699 256961 298728 256989
rect 298756 256961 298790 256989
rect 298818 256961 298852 256989
rect 298880 256961 298914 256989
rect 298942 256961 298990 256989
rect -958 256913 298990 256961
rect -958 254175 298990 254223
rect -958 254147 -430 254175
rect -402 254147 -368 254175
rect -340 254147 -306 254175
rect -278 254147 -244 254175
rect -216 254147 1625 254175
rect 1653 254147 1687 254175
rect 1715 254147 1749 254175
rect 1777 254147 1811 254175
rect 1839 254147 10625 254175
rect 10653 254147 10687 254175
rect 10715 254147 10749 254175
rect 10777 254147 10811 254175
rect 10839 254147 19625 254175
rect 19653 254147 19687 254175
rect 19715 254147 19749 254175
rect 19777 254147 19811 254175
rect 19839 254147 28625 254175
rect 28653 254147 28687 254175
rect 28715 254147 28749 254175
rect 28777 254147 28811 254175
rect 28839 254147 37625 254175
rect 37653 254147 37687 254175
rect 37715 254147 37749 254175
rect 37777 254147 37811 254175
rect 37839 254147 46625 254175
rect 46653 254147 46687 254175
rect 46715 254147 46749 254175
rect 46777 254147 46811 254175
rect 46839 254147 52259 254175
rect 52287 254147 52321 254175
rect 52349 254147 67619 254175
rect 67647 254147 67681 254175
rect 67709 254147 82979 254175
rect 83007 254147 83041 254175
rect 83069 254147 98339 254175
rect 98367 254147 98401 254175
rect 98429 254147 113699 254175
rect 113727 254147 113761 254175
rect 113789 254147 129059 254175
rect 129087 254147 129121 254175
rect 129149 254147 144419 254175
rect 144447 254147 144481 254175
rect 144509 254147 154625 254175
rect 154653 254147 154687 254175
rect 154715 254147 154749 254175
rect 154777 254147 154811 254175
rect 154839 254147 163625 254175
rect 163653 254147 163687 254175
rect 163715 254147 163749 254175
rect 163777 254147 163811 254175
rect 163839 254147 172625 254175
rect 172653 254147 172687 254175
rect 172715 254147 172749 254175
rect 172777 254147 172811 254175
rect 172839 254147 181625 254175
rect 181653 254147 181687 254175
rect 181715 254147 181749 254175
rect 181777 254147 181811 254175
rect 181839 254147 190625 254175
rect 190653 254147 190687 254175
rect 190715 254147 190749 254175
rect 190777 254147 190811 254175
rect 190839 254147 199625 254175
rect 199653 254147 199687 254175
rect 199715 254147 199749 254175
rect 199777 254147 199811 254175
rect 199839 254147 208625 254175
rect 208653 254147 208687 254175
rect 208715 254147 208749 254175
rect 208777 254147 208811 254175
rect 208839 254147 217625 254175
rect 217653 254147 217687 254175
rect 217715 254147 217749 254175
rect 217777 254147 217811 254175
rect 217839 254147 226625 254175
rect 226653 254147 226687 254175
rect 226715 254147 226749 254175
rect 226777 254147 226811 254175
rect 226839 254147 235625 254175
rect 235653 254147 235687 254175
rect 235715 254147 235749 254175
rect 235777 254147 235811 254175
rect 235839 254147 244625 254175
rect 244653 254147 244687 254175
rect 244715 254147 244749 254175
rect 244777 254147 244811 254175
rect 244839 254147 253625 254175
rect 253653 254147 253687 254175
rect 253715 254147 253749 254175
rect 253777 254147 253811 254175
rect 253839 254147 262625 254175
rect 262653 254147 262687 254175
rect 262715 254147 262749 254175
rect 262777 254147 262811 254175
rect 262839 254147 271625 254175
rect 271653 254147 271687 254175
rect 271715 254147 271749 254175
rect 271777 254147 271811 254175
rect 271839 254147 280625 254175
rect 280653 254147 280687 254175
rect 280715 254147 280749 254175
rect 280777 254147 280811 254175
rect 280839 254147 289625 254175
rect 289653 254147 289687 254175
rect 289715 254147 289749 254175
rect 289777 254147 289811 254175
rect 289839 254147 298248 254175
rect 298276 254147 298310 254175
rect 298338 254147 298372 254175
rect 298400 254147 298434 254175
rect 298462 254147 298990 254175
rect -958 254113 298990 254147
rect -958 254085 -430 254113
rect -402 254085 -368 254113
rect -340 254085 -306 254113
rect -278 254085 -244 254113
rect -216 254085 1625 254113
rect 1653 254085 1687 254113
rect 1715 254085 1749 254113
rect 1777 254085 1811 254113
rect 1839 254085 10625 254113
rect 10653 254085 10687 254113
rect 10715 254085 10749 254113
rect 10777 254085 10811 254113
rect 10839 254085 19625 254113
rect 19653 254085 19687 254113
rect 19715 254085 19749 254113
rect 19777 254085 19811 254113
rect 19839 254085 28625 254113
rect 28653 254085 28687 254113
rect 28715 254085 28749 254113
rect 28777 254085 28811 254113
rect 28839 254085 37625 254113
rect 37653 254085 37687 254113
rect 37715 254085 37749 254113
rect 37777 254085 37811 254113
rect 37839 254085 46625 254113
rect 46653 254085 46687 254113
rect 46715 254085 46749 254113
rect 46777 254085 46811 254113
rect 46839 254085 52259 254113
rect 52287 254085 52321 254113
rect 52349 254085 67619 254113
rect 67647 254085 67681 254113
rect 67709 254085 82979 254113
rect 83007 254085 83041 254113
rect 83069 254085 98339 254113
rect 98367 254085 98401 254113
rect 98429 254085 113699 254113
rect 113727 254085 113761 254113
rect 113789 254085 129059 254113
rect 129087 254085 129121 254113
rect 129149 254085 144419 254113
rect 144447 254085 144481 254113
rect 144509 254085 154625 254113
rect 154653 254085 154687 254113
rect 154715 254085 154749 254113
rect 154777 254085 154811 254113
rect 154839 254085 163625 254113
rect 163653 254085 163687 254113
rect 163715 254085 163749 254113
rect 163777 254085 163811 254113
rect 163839 254085 172625 254113
rect 172653 254085 172687 254113
rect 172715 254085 172749 254113
rect 172777 254085 172811 254113
rect 172839 254085 181625 254113
rect 181653 254085 181687 254113
rect 181715 254085 181749 254113
rect 181777 254085 181811 254113
rect 181839 254085 190625 254113
rect 190653 254085 190687 254113
rect 190715 254085 190749 254113
rect 190777 254085 190811 254113
rect 190839 254085 199625 254113
rect 199653 254085 199687 254113
rect 199715 254085 199749 254113
rect 199777 254085 199811 254113
rect 199839 254085 208625 254113
rect 208653 254085 208687 254113
rect 208715 254085 208749 254113
rect 208777 254085 208811 254113
rect 208839 254085 217625 254113
rect 217653 254085 217687 254113
rect 217715 254085 217749 254113
rect 217777 254085 217811 254113
rect 217839 254085 226625 254113
rect 226653 254085 226687 254113
rect 226715 254085 226749 254113
rect 226777 254085 226811 254113
rect 226839 254085 235625 254113
rect 235653 254085 235687 254113
rect 235715 254085 235749 254113
rect 235777 254085 235811 254113
rect 235839 254085 244625 254113
rect 244653 254085 244687 254113
rect 244715 254085 244749 254113
rect 244777 254085 244811 254113
rect 244839 254085 253625 254113
rect 253653 254085 253687 254113
rect 253715 254085 253749 254113
rect 253777 254085 253811 254113
rect 253839 254085 262625 254113
rect 262653 254085 262687 254113
rect 262715 254085 262749 254113
rect 262777 254085 262811 254113
rect 262839 254085 271625 254113
rect 271653 254085 271687 254113
rect 271715 254085 271749 254113
rect 271777 254085 271811 254113
rect 271839 254085 280625 254113
rect 280653 254085 280687 254113
rect 280715 254085 280749 254113
rect 280777 254085 280811 254113
rect 280839 254085 289625 254113
rect 289653 254085 289687 254113
rect 289715 254085 289749 254113
rect 289777 254085 289811 254113
rect 289839 254085 298248 254113
rect 298276 254085 298310 254113
rect 298338 254085 298372 254113
rect 298400 254085 298434 254113
rect 298462 254085 298990 254113
rect -958 254051 298990 254085
rect -958 254023 -430 254051
rect -402 254023 -368 254051
rect -340 254023 -306 254051
rect -278 254023 -244 254051
rect -216 254023 1625 254051
rect 1653 254023 1687 254051
rect 1715 254023 1749 254051
rect 1777 254023 1811 254051
rect 1839 254023 10625 254051
rect 10653 254023 10687 254051
rect 10715 254023 10749 254051
rect 10777 254023 10811 254051
rect 10839 254023 19625 254051
rect 19653 254023 19687 254051
rect 19715 254023 19749 254051
rect 19777 254023 19811 254051
rect 19839 254023 28625 254051
rect 28653 254023 28687 254051
rect 28715 254023 28749 254051
rect 28777 254023 28811 254051
rect 28839 254023 37625 254051
rect 37653 254023 37687 254051
rect 37715 254023 37749 254051
rect 37777 254023 37811 254051
rect 37839 254023 46625 254051
rect 46653 254023 46687 254051
rect 46715 254023 46749 254051
rect 46777 254023 46811 254051
rect 46839 254023 52259 254051
rect 52287 254023 52321 254051
rect 52349 254023 67619 254051
rect 67647 254023 67681 254051
rect 67709 254023 82979 254051
rect 83007 254023 83041 254051
rect 83069 254023 98339 254051
rect 98367 254023 98401 254051
rect 98429 254023 113699 254051
rect 113727 254023 113761 254051
rect 113789 254023 129059 254051
rect 129087 254023 129121 254051
rect 129149 254023 144419 254051
rect 144447 254023 144481 254051
rect 144509 254023 154625 254051
rect 154653 254023 154687 254051
rect 154715 254023 154749 254051
rect 154777 254023 154811 254051
rect 154839 254023 163625 254051
rect 163653 254023 163687 254051
rect 163715 254023 163749 254051
rect 163777 254023 163811 254051
rect 163839 254023 172625 254051
rect 172653 254023 172687 254051
rect 172715 254023 172749 254051
rect 172777 254023 172811 254051
rect 172839 254023 181625 254051
rect 181653 254023 181687 254051
rect 181715 254023 181749 254051
rect 181777 254023 181811 254051
rect 181839 254023 190625 254051
rect 190653 254023 190687 254051
rect 190715 254023 190749 254051
rect 190777 254023 190811 254051
rect 190839 254023 199625 254051
rect 199653 254023 199687 254051
rect 199715 254023 199749 254051
rect 199777 254023 199811 254051
rect 199839 254023 208625 254051
rect 208653 254023 208687 254051
rect 208715 254023 208749 254051
rect 208777 254023 208811 254051
rect 208839 254023 217625 254051
rect 217653 254023 217687 254051
rect 217715 254023 217749 254051
rect 217777 254023 217811 254051
rect 217839 254023 226625 254051
rect 226653 254023 226687 254051
rect 226715 254023 226749 254051
rect 226777 254023 226811 254051
rect 226839 254023 235625 254051
rect 235653 254023 235687 254051
rect 235715 254023 235749 254051
rect 235777 254023 235811 254051
rect 235839 254023 244625 254051
rect 244653 254023 244687 254051
rect 244715 254023 244749 254051
rect 244777 254023 244811 254051
rect 244839 254023 253625 254051
rect 253653 254023 253687 254051
rect 253715 254023 253749 254051
rect 253777 254023 253811 254051
rect 253839 254023 262625 254051
rect 262653 254023 262687 254051
rect 262715 254023 262749 254051
rect 262777 254023 262811 254051
rect 262839 254023 271625 254051
rect 271653 254023 271687 254051
rect 271715 254023 271749 254051
rect 271777 254023 271811 254051
rect 271839 254023 280625 254051
rect 280653 254023 280687 254051
rect 280715 254023 280749 254051
rect 280777 254023 280811 254051
rect 280839 254023 289625 254051
rect 289653 254023 289687 254051
rect 289715 254023 289749 254051
rect 289777 254023 289811 254051
rect 289839 254023 298248 254051
rect 298276 254023 298310 254051
rect 298338 254023 298372 254051
rect 298400 254023 298434 254051
rect 298462 254023 298990 254051
rect -958 253989 298990 254023
rect -958 253961 -430 253989
rect -402 253961 -368 253989
rect -340 253961 -306 253989
rect -278 253961 -244 253989
rect -216 253961 1625 253989
rect 1653 253961 1687 253989
rect 1715 253961 1749 253989
rect 1777 253961 1811 253989
rect 1839 253961 10625 253989
rect 10653 253961 10687 253989
rect 10715 253961 10749 253989
rect 10777 253961 10811 253989
rect 10839 253961 19625 253989
rect 19653 253961 19687 253989
rect 19715 253961 19749 253989
rect 19777 253961 19811 253989
rect 19839 253961 28625 253989
rect 28653 253961 28687 253989
rect 28715 253961 28749 253989
rect 28777 253961 28811 253989
rect 28839 253961 37625 253989
rect 37653 253961 37687 253989
rect 37715 253961 37749 253989
rect 37777 253961 37811 253989
rect 37839 253961 46625 253989
rect 46653 253961 46687 253989
rect 46715 253961 46749 253989
rect 46777 253961 46811 253989
rect 46839 253961 52259 253989
rect 52287 253961 52321 253989
rect 52349 253961 67619 253989
rect 67647 253961 67681 253989
rect 67709 253961 82979 253989
rect 83007 253961 83041 253989
rect 83069 253961 98339 253989
rect 98367 253961 98401 253989
rect 98429 253961 113699 253989
rect 113727 253961 113761 253989
rect 113789 253961 129059 253989
rect 129087 253961 129121 253989
rect 129149 253961 144419 253989
rect 144447 253961 144481 253989
rect 144509 253961 154625 253989
rect 154653 253961 154687 253989
rect 154715 253961 154749 253989
rect 154777 253961 154811 253989
rect 154839 253961 163625 253989
rect 163653 253961 163687 253989
rect 163715 253961 163749 253989
rect 163777 253961 163811 253989
rect 163839 253961 172625 253989
rect 172653 253961 172687 253989
rect 172715 253961 172749 253989
rect 172777 253961 172811 253989
rect 172839 253961 181625 253989
rect 181653 253961 181687 253989
rect 181715 253961 181749 253989
rect 181777 253961 181811 253989
rect 181839 253961 190625 253989
rect 190653 253961 190687 253989
rect 190715 253961 190749 253989
rect 190777 253961 190811 253989
rect 190839 253961 199625 253989
rect 199653 253961 199687 253989
rect 199715 253961 199749 253989
rect 199777 253961 199811 253989
rect 199839 253961 208625 253989
rect 208653 253961 208687 253989
rect 208715 253961 208749 253989
rect 208777 253961 208811 253989
rect 208839 253961 217625 253989
rect 217653 253961 217687 253989
rect 217715 253961 217749 253989
rect 217777 253961 217811 253989
rect 217839 253961 226625 253989
rect 226653 253961 226687 253989
rect 226715 253961 226749 253989
rect 226777 253961 226811 253989
rect 226839 253961 235625 253989
rect 235653 253961 235687 253989
rect 235715 253961 235749 253989
rect 235777 253961 235811 253989
rect 235839 253961 244625 253989
rect 244653 253961 244687 253989
rect 244715 253961 244749 253989
rect 244777 253961 244811 253989
rect 244839 253961 253625 253989
rect 253653 253961 253687 253989
rect 253715 253961 253749 253989
rect 253777 253961 253811 253989
rect 253839 253961 262625 253989
rect 262653 253961 262687 253989
rect 262715 253961 262749 253989
rect 262777 253961 262811 253989
rect 262839 253961 271625 253989
rect 271653 253961 271687 253989
rect 271715 253961 271749 253989
rect 271777 253961 271811 253989
rect 271839 253961 280625 253989
rect 280653 253961 280687 253989
rect 280715 253961 280749 253989
rect 280777 253961 280811 253989
rect 280839 253961 289625 253989
rect 289653 253961 289687 253989
rect 289715 253961 289749 253989
rect 289777 253961 289811 253989
rect 289839 253961 298248 253989
rect 298276 253961 298310 253989
rect 298338 253961 298372 253989
rect 298400 253961 298434 253989
rect 298462 253961 298990 253989
rect -958 253913 298990 253961
rect -958 248175 298990 248223
rect -958 248147 -910 248175
rect -882 248147 -848 248175
rect -820 248147 -786 248175
rect -758 248147 -724 248175
rect -696 248147 3485 248175
rect 3513 248147 3547 248175
rect 3575 248147 3609 248175
rect 3637 248147 3671 248175
rect 3699 248147 12485 248175
rect 12513 248147 12547 248175
rect 12575 248147 12609 248175
rect 12637 248147 12671 248175
rect 12699 248147 21485 248175
rect 21513 248147 21547 248175
rect 21575 248147 21609 248175
rect 21637 248147 21671 248175
rect 21699 248147 30485 248175
rect 30513 248147 30547 248175
rect 30575 248147 30609 248175
rect 30637 248147 30671 248175
rect 30699 248147 39485 248175
rect 39513 248147 39547 248175
rect 39575 248147 39609 248175
rect 39637 248147 39671 248175
rect 39699 248147 48485 248175
rect 48513 248147 48547 248175
rect 48575 248147 48609 248175
rect 48637 248147 48671 248175
rect 48699 248147 59939 248175
rect 59967 248147 60001 248175
rect 60029 248147 75299 248175
rect 75327 248147 75361 248175
rect 75389 248147 90659 248175
rect 90687 248147 90721 248175
rect 90749 248147 106019 248175
rect 106047 248147 106081 248175
rect 106109 248147 121379 248175
rect 121407 248147 121441 248175
rect 121469 248147 136739 248175
rect 136767 248147 136801 248175
rect 136829 248147 156485 248175
rect 156513 248147 156547 248175
rect 156575 248147 156609 248175
rect 156637 248147 156671 248175
rect 156699 248147 165485 248175
rect 165513 248147 165547 248175
rect 165575 248147 165609 248175
rect 165637 248147 165671 248175
rect 165699 248147 174485 248175
rect 174513 248147 174547 248175
rect 174575 248147 174609 248175
rect 174637 248147 174671 248175
rect 174699 248147 183485 248175
rect 183513 248147 183547 248175
rect 183575 248147 183609 248175
rect 183637 248147 183671 248175
rect 183699 248147 192485 248175
rect 192513 248147 192547 248175
rect 192575 248147 192609 248175
rect 192637 248147 192671 248175
rect 192699 248147 201485 248175
rect 201513 248147 201547 248175
rect 201575 248147 201609 248175
rect 201637 248147 201671 248175
rect 201699 248147 210485 248175
rect 210513 248147 210547 248175
rect 210575 248147 210609 248175
rect 210637 248147 210671 248175
rect 210699 248147 219485 248175
rect 219513 248147 219547 248175
rect 219575 248147 219609 248175
rect 219637 248147 219671 248175
rect 219699 248147 228485 248175
rect 228513 248147 228547 248175
rect 228575 248147 228609 248175
rect 228637 248147 228671 248175
rect 228699 248147 237485 248175
rect 237513 248147 237547 248175
rect 237575 248147 237609 248175
rect 237637 248147 237671 248175
rect 237699 248147 246485 248175
rect 246513 248147 246547 248175
rect 246575 248147 246609 248175
rect 246637 248147 246671 248175
rect 246699 248147 255485 248175
rect 255513 248147 255547 248175
rect 255575 248147 255609 248175
rect 255637 248147 255671 248175
rect 255699 248147 264485 248175
rect 264513 248147 264547 248175
rect 264575 248147 264609 248175
rect 264637 248147 264671 248175
rect 264699 248147 273485 248175
rect 273513 248147 273547 248175
rect 273575 248147 273609 248175
rect 273637 248147 273671 248175
rect 273699 248147 282485 248175
rect 282513 248147 282547 248175
rect 282575 248147 282609 248175
rect 282637 248147 282671 248175
rect 282699 248147 291485 248175
rect 291513 248147 291547 248175
rect 291575 248147 291609 248175
rect 291637 248147 291671 248175
rect 291699 248147 298728 248175
rect 298756 248147 298790 248175
rect 298818 248147 298852 248175
rect 298880 248147 298914 248175
rect 298942 248147 298990 248175
rect -958 248113 298990 248147
rect -958 248085 -910 248113
rect -882 248085 -848 248113
rect -820 248085 -786 248113
rect -758 248085 -724 248113
rect -696 248085 3485 248113
rect 3513 248085 3547 248113
rect 3575 248085 3609 248113
rect 3637 248085 3671 248113
rect 3699 248085 12485 248113
rect 12513 248085 12547 248113
rect 12575 248085 12609 248113
rect 12637 248085 12671 248113
rect 12699 248085 21485 248113
rect 21513 248085 21547 248113
rect 21575 248085 21609 248113
rect 21637 248085 21671 248113
rect 21699 248085 30485 248113
rect 30513 248085 30547 248113
rect 30575 248085 30609 248113
rect 30637 248085 30671 248113
rect 30699 248085 39485 248113
rect 39513 248085 39547 248113
rect 39575 248085 39609 248113
rect 39637 248085 39671 248113
rect 39699 248085 48485 248113
rect 48513 248085 48547 248113
rect 48575 248085 48609 248113
rect 48637 248085 48671 248113
rect 48699 248085 59939 248113
rect 59967 248085 60001 248113
rect 60029 248085 75299 248113
rect 75327 248085 75361 248113
rect 75389 248085 90659 248113
rect 90687 248085 90721 248113
rect 90749 248085 106019 248113
rect 106047 248085 106081 248113
rect 106109 248085 121379 248113
rect 121407 248085 121441 248113
rect 121469 248085 136739 248113
rect 136767 248085 136801 248113
rect 136829 248085 156485 248113
rect 156513 248085 156547 248113
rect 156575 248085 156609 248113
rect 156637 248085 156671 248113
rect 156699 248085 165485 248113
rect 165513 248085 165547 248113
rect 165575 248085 165609 248113
rect 165637 248085 165671 248113
rect 165699 248085 174485 248113
rect 174513 248085 174547 248113
rect 174575 248085 174609 248113
rect 174637 248085 174671 248113
rect 174699 248085 183485 248113
rect 183513 248085 183547 248113
rect 183575 248085 183609 248113
rect 183637 248085 183671 248113
rect 183699 248085 192485 248113
rect 192513 248085 192547 248113
rect 192575 248085 192609 248113
rect 192637 248085 192671 248113
rect 192699 248085 201485 248113
rect 201513 248085 201547 248113
rect 201575 248085 201609 248113
rect 201637 248085 201671 248113
rect 201699 248085 210485 248113
rect 210513 248085 210547 248113
rect 210575 248085 210609 248113
rect 210637 248085 210671 248113
rect 210699 248085 219485 248113
rect 219513 248085 219547 248113
rect 219575 248085 219609 248113
rect 219637 248085 219671 248113
rect 219699 248085 228485 248113
rect 228513 248085 228547 248113
rect 228575 248085 228609 248113
rect 228637 248085 228671 248113
rect 228699 248085 237485 248113
rect 237513 248085 237547 248113
rect 237575 248085 237609 248113
rect 237637 248085 237671 248113
rect 237699 248085 246485 248113
rect 246513 248085 246547 248113
rect 246575 248085 246609 248113
rect 246637 248085 246671 248113
rect 246699 248085 255485 248113
rect 255513 248085 255547 248113
rect 255575 248085 255609 248113
rect 255637 248085 255671 248113
rect 255699 248085 264485 248113
rect 264513 248085 264547 248113
rect 264575 248085 264609 248113
rect 264637 248085 264671 248113
rect 264699 248085 273485 248113
rect 273513 248085 273547 248113
rect 273575 248085 273609 248113
rect 273637 248085 273671 248113
rect 273699 248085 282485 248113
rect 282513 248085 282547 248113
rect 282575 248085 282609 248113
rect 282637 248085 282671 248113
rect 282699 248085 291485 248113
rect 291513 248085 291547 248113
rect 291575 248085 291609 248113
rect 291637 248085 291671 248113
rect 291699 248085 298728 248113
rect 298756 248085 298790 248113
rect 298818 248085 298852 248113
rect 298880 248085 298914 248113
rect 298942 248085 298990 248113
rect -958 248051 298990 248085
rect -958 248023 -910 248051
rect -882 248023 -848 248051
rect -820 248023 -786 248051
rect -758 248023 -724 248051
rect -696 248023 3485 248051
rect 3513 248023 3547 248051
rect 3575 248023 3609 248051
rect 3637 248023 3671 248051
rect 3699 248023 12485 248051
rect 12513 248023 12547 248051
rect 12575 248023 12609 248051
rect 12637 248023 12671 248051
rect 12699 248023 21485 248051
rect 21513 248023 21547 248051
rect 21575 248023 21609 248051
rect 21637 248023 21671 248051
rect 21699 248023 30485 248051
rect 30513 248023 30547 248051
rect 30575 248023 30609 248051
rect 30637 248023 30671 248051
rect 30699 248023 39485 248051
rect 39513 248023 39547 248051
rect 39575 248023 39609 248051
rect 39637 248023 39671 248051
rect 39699 248023 48485 248051
rect 48513 248023 48547 248051
rect 48575 248023 48609 248051
rect 48637 248023 48671 248051
rect 48699 248023 59939 248051
rect 59967 248023 60001 248051
rect 60029 248023 75299 248051
rect 75327 248023 75361 248051
rect 75389 248023 90659 248051
rect 90687 248023 90721 248051
rect 90749 248023 106019 248051
rect 106047 248023 106081 248051
rect 106109 248023 121379 248051
rect 121407 248023 121441 248051
rect 121469 248023 136739 248051
rect 136767 248023 136801 248051
rect 136829 248023 156485 248051
rect 156513 248023 156547 248051
rect 156575 248023 156609 248051
rect 156637 248023 156671 248051
rect 156699 248023 165485 248051
rect 165513 248023 165547 248051
rect 165575 248023 165609 248051
rect 165637 248023 165671 248051
rect 165699 248023 174485 248051
rect 174513 248023 174547 248051
rect 174575 248023 174609 248051
rect 174637 248023 174671 248051
rect 174699 248023 183485 248051
rect 183513 248023 183547 248051
rect 183575 248023 183609 248051
rect 183637 248023 183671 248051
rect 183699 248023 192485 248051
rect 192513 248023 192547 248051
rect 192575 248023 192609 248051
rect 192637 248023 192671 248051
rect 192699 248023 201485 248051
rect 201513 248023 201547 248051
rect 201575 248023 201609 248051
rect 201637 248023 201671 248051
rect 201699 248023 210485 248051
rect 210513 248023 210547 248051
rect 210575 248023 210609 248051
rect 210637 248023 210671 248051
rect 210699 248023 219485 248051
rect 219513 248023 219547 248051
rect 219575 248023 219609 248051
rect 219637 248023 219671 248051
rect 219699 248023 228485 248051
rect 228513 248023 228547 248051
rect 228575 248023 228609 248051
rect 228637 248023 228671 248051
rect 228699 248023 237485 248051
rect 237513 248023 237547 248051
rect 237575 248023 237609 248051
rect 237637 248023 237671 248051
rect 237699 248023 246485 248051
rect 246513 248023 246547 248051
rect 246575 248023 246609 248051
rect 246637 248023 246671 248051
rect 246699 248023 255485 248051
rect 255513 248023 255547 248051
rect 255575 248023 255609 248051
rect 255637 248023 255671 248051
rect 255699 248023 264485 248051
rect 264513 248023 264547 248051
rect 264575 248023 264609 248051
rect 264637 248023 264671 248051
rect 264699 248023 273485 248051
rect 273513 248023 273547 248051
rect 273575 248023 273609 248051
rect 273637 248023 273671 248051
rect 273699 248023 282485 248051
rect 282513 248023 282547 248051
rect 282575 248023 282609 248051
rect 282637 248023 282671 248051
rect 282699 248023 291485 248051
rect 291513 248023 291547 248051
rect 291575 248023 291609 248051
rect 291637 248023 291671 248051
rect 291699 248023 298728 248051
rect 298756 248023 298790 248051
rect 298818 248023 298852 248051
rect 298880 248023 298914 248051
rect 298942 248023 298990 248051
rect -958 247989 298990 248023
rect -958 247961 -910 247989
rect -882 247961 -848 247989
rect -820 247961 -786 247989
rect -758 247961 -724 247989
rect -696 247961 3485 247989
rect 3513 247961 3547 247989
rect 3575 247961 3609 247989
rect 3637 247961 3671 247989
rect 3699 247961 12485 247989
rect 12513 247961 12547 247989
rect 12575 247961 12609 247989
rect 12637 247961 12671 247989
rect 12699 247961 21485 247989
rect 21513 247961 21547 247989
rect 21575 247961 21609 247989
rect 21637 247961 21671 247989
rect 21699 247961 30485 247989
rect 30513 247961 30547 247989
rect 30575 247961 30609 247989
rect 30637 247961 30671 247989
rect 30699 247961 39485 247989
rect 39513 247961 39547 247989
rect 39575 247961 39609 247989
rect 39637 247961 39671 247989
rect 39699 247961 48485 247989
rect 48513 247961 48547 247989
rect 48575 247961 48609 247989
rect 48637 247961 48671 247989
rect 48699 247961 59939 247989
rect 59967 247961 60001 247989
rect 60029 247961 75299 247989
rect 75327 247961 75361 247989
rect 75389 247961 90659 247989
rect 90687 247961 90721 247989
rect 90749 247961 106019 247989
rect 106047 247961 106081 247989
rect 106109 247961 121379 247989
rect 121407 247961 121441 247989
rect 121469 247961 136739 247989
rect 136767 247961 136801 247989
rect 136829 247961 156485 247989
rect 156513 247961 156547 247989
rect 156575 247961 156609 247989
rect 156637 247961 156671 247989
rect 156699 247961 165485 247989
rect 165513 247961 165547 247989
rect 165575 247961 165609 247989
rect 165637 247961 165671 247989
rect 165699 247961 174485 247989
rect 174513 247961 174547 247989
rect 174575 247961 174609 247989
rect 174637 247961 174671 247989
rect 174699 247961 183485 247989
rect 183513 247961 183547 247989
rect 183575 247961 183609 247989
rect 183637 247961 183671 247989
rect 183699 247961 192485 247989
rect 192513 247961 192547 247989
rect 192575 247961 192609 247989
rect 192637 247961 192671 247989
rect 192699 247961 201485 247989
rect 201513 247961 201547 247989
rect 201575 247961 201609 247989
rect 201637 247961 201671 247989
rect 201699 247961 210485 247989
rect 210513 247961 210547 247989
rect 210575 247961 210609 247989
rect 210637 247961 210671 247989
rect 210699 247961 219485 247989
rect 219513 247961 219547 247989
rect 219575 247961 219609 247989
rect 219637 247961 219671 247989
rect 219699 247961 228485 247989
rect 228513 247961 228547 247989
rect 228575 247961 228609 247989
rect 228637 247961 228671 247989
rect 228699 247961 237485 247989
rect 237513 247961 237547 247989
rect 237575 247961 237609 247989
rect 237637 247961 237671 247989
rect 237699 247961 246485 247989
rect 246513 247961 246547 247989
rect 246575 247961 246609 247989
rect 246637 247961 246671 247989
rect 246699 247961 255485 247989
rect 255513 247961 255547 247989
rect 255575 247961 255609 247989
rect 255637 247961 255671 247989
rect 255699 247961 264485 247989
rect 264513 247961 264547 247989
rect 264575 247961 264609 247989
rect 264637 247961 264671 247989
rect 264699 247961 273485 247989
rect 273513 247961 273547 247989
rect 273575 247961 273609 247989
rect 273637 247961 273671 247989
rect 273699 247961 282485 247989
rect 282513 247961 282547 247989
rect 282575 247961 282609 247989
rect 282637 247961 282671 247989
rect 282699 247961 291485 247989
rect 291513 247961 291547 247989
rect 291575 247961 291609 247989
rect 291637 247961 291671 247989
rect 291699 247961 298728 247989
rect 298756 247961 298790 247989
rect 298818 247961 298852 247989
rect 298880 247961 298914 247989
rect 298942 247961 298990 247989
rect -958 247913 298990 247961
rect -958 245175 298990 245223
rect -958 245147 -430 245175
rect -402 245147 -368 245175
rect -340 245147 -306 245175
rect -278 245147 -244 245175
rect -216 245147 1625 245175
rect 1653 245147 1687 245175
rect 1715 245147 1749 245175
rect 1777 245147 1811 245175
rect 1839 245147 10625 245175
rect 10653 245147 10687 245175
rect 10715 245147 10749 245175
rect 10777 245147 10811 245175
rect 10839 245147 19625 245175
rect 19653 245147 19687 245175
rect 19715 245147 19749 245175
rect 19777 245147 19811 245175
rect 19839 245147 28625 245175
rect 28653 245147 28687 245175
rect 28715 245147 28749 245175
rect 28777 245147 28811 245175
rect 28839 245147 37625 245175
rect 37653 245147 37687 245175
rect 37715 245147 37749 245175
rect 37777 245147 37811 245175
rect 37839 245147 46625 245175
rect 46653 245147 46687 245175
rect 46715 245147 46749 245175
rect 46777 245147 46811 245175
rect 46839 245147 52259 245175
rect 52287 245147 52321 245175
rect 52349 245147 67619 245175
rect 67647 245147 67681 245175
rect 67709 245147 82979 245175
rect 83007 245147 83041 245175
rect 83069 245147 98339 245175
rect 98367 245147 98401 245175
rect 98429 245147 113699 245175
rect 113727 245147 113761 245175
rect 113789 245147 129059 245175
rect 129087 245147 129121 245175
rect 129149 245147 144419 245175
rect 144447 245147 144481 245175
rect 144509 245147 154625 245175
rect 154653 245147 154687 245175
rect 154715 245147 154749 245175
rect 154777 245147 154811 245175
rect 154839 245147 163625 245175
rect 163653 245147 163687 245175
rect 163715 245147 163749 245175
rect 163777 245147 163811 245175
rect 163839 245147 172625 245175
rect 172653 245147 172687 245175
rect 172715 245147 172749 245175
rect 172777 245147 172811 245175
rect 172839 245147 181625 245175
rect 181653 245147 181687 245175
rect 181715 245147 181749 245175
rect 181777 245147 181811 245175
rect 181839 245147 190625 245175
rect 190653 245147 190687 245175
rect 190715 245147 190749 245175
rect 190777 245147 190811 245175
rect 190839 245147 199625 245175
rect 199653 245147 199687 245175
rect 199715 245147 199749 245175
rect 199777 245147 199811 245175
rect 199839 245147 208625 245175
rect 208653 245147 208687 245175
rect 208715 245147 208749 245175
rect 208777 245147 208811 245175
rect 208839 245147 217625 245175
rect 217653 245147 217687 245175
rect 217715 245147 217749 245175
rect 217777 245147 217811 245175
rect 217839 245147 226625 245175
rect 226653 245147 226687 245175
rect 226715 245147 226749 245175
rect 226777 245147 226811 245175
rect 226839 245147 235625 245175
rect 235653 245147 235687 245175
rect 235715 245147 235749 245175
rect 235777 245147 235811 245175
rect 235839 245147 244625 245175
rect 244653 245147 244687 245175
rect 244715 245147 244749 245175
rect 244777 245147 244811 245175
rect 244839 245147 253625 245175
rect 253653 245147 253687 245175
rect 253715 245147 253749 245175
rect 253777 245147 253811 245175
rect 253839 245147 262625 245175
rect 262653 245147 262687 245175
rect 262715 245147 262749 245175
rect 262777 245147 262811 245175
rect 262839 245147 271625 245175
rect 271653 245147 271687 245175
rect 271715 245147 271749 245175
rect 271777 245147 271811 245175
rect 271839 245147 280625 245175
rect 280653 245147 280687 245175
rect 280715 245147 280749 245175
rect 280777 245147 280811 245175
rect 280839 245147 289625 245175
rect 289653 245147 289687 245175
rect 289715 245147 289749 245175
rect 289777 245147 289811 245175
rect 289839 245147 298248 245175
rect 298276 245147 298310 245175
rect 298338 245147 298372 245175
rect 298400 245147 298434 245175
rect 298462 245147 298990 245175
rect -958 245113 298990 245147
rect -958 245085 -430 245113
rect -402 245085 -368 245113
rect -340 245085 -306 245113
rect -278 245085 -244 245113
rect -216 245085 1625 245113
rect 1653 245085 1687 245113
rect 1715 245085 1749 245113
rect 1777 245085 1811 245113
rect 1839 245085 10625 245113
rect 10653 245085 10687 245113
rect 10715 245085 10749 245113
rect 10777 245085 10811 245113
rect 10839 245085 19625 245113
rect 19653 245085 19687 245113
rect 19715 245085 19749 245113
rect 19777 245085 19811 245113
rect 19839 245085 28625 245113
rect 28653 245085 28687 245113
rect 28715 245085 28749 245113
rect 28777 245085 28811 245113
rect 28839 245085 37625 245113
rect 37653 245085 37687 245113
rect 37715 245085 37749 245113
rect 37777 245085 37811 245113
rect 37839 245085 46625 245113
rect 46653 245085 46687 245113
rect 46715 245085 46749 245113
rect 46777 245085 46811 245113
rect 46839 245085 52259 245113
rect 52287 245085 52321 245113
rect 52349 245085 67619 245113
rect 67647 245085 67681 245113
rect 67709 245085 82979 245113
rect 83007 245085 83041 245113
rect 83069 245085 98339 245113
rect 98367 245085 98401 245113
rect 98429 245085 113699 245113
rect 113727 245085 113761 245113
rect 113789 245085 129059 245113
rect 129087 245085 129121 245113
rect 129149 245085 144419 245113
rect 144447 245085 144481 245113
rect 144509 245085 154625 245113
rect 154653 245085 154687 245113
rect 154715 245085 154749 245113
rect 154777 245085 154811 245113
rect 154839 245085 163625 245113
rect 163653 245085 163687 245113
rect 163715 245085 163749 245113
rect 163777 245085 163811 245113
rect 163839 245085 172625 245113
rect 172653 245085 172687 245113
rect 172715 245085 172749 245113
rect 172777 245085 172811 245113
rect 172839 245085 181625 245113
rect 181653 245085 181687 245113
rect 181715 245085 181749 245113
rect 181777 245085 181811 245113
rect 181839 245085 190625 245113
rect 190653 245085 190687 245113
rect 190715 245085 190749 245113
rect 190777 245085 190811 245113
rect 190839 245085 199625 245113
rect 199653 245085 199687 245113
rect 199715 245085 199749 245113
rect 199777 245085 199811 245113
rect 199839 245085 208625 245113
rect 208653 245085 208687 245113
rect 208715 245085 208749 245113
rect 208777 245085 208811 245113
rect 208839 245085 217625 245113
rect 217653 245085 217687 245113
rect 217715 245085 217749 245113
rect 217777 245085 217811 245113
rect 217839 245085 226625 245113
rect 226653 245085 226687 245113
rect 226715 245085 226749 245113
rect 226777 245085 226811 245113
rect 226839 245085 235625 245113
rect 235653 245085 235687 245113
rect 235715 245085 235749 245113
rect 235777 245085 235811 245113
rect 235839 245085 244625 245113
rect 244653 245085 244687 245113
rect 244715 245085 244749 245113
rect 244777 245085 244811 245113
rect 244839 245085 253625 245113
rect 253653 245085 253687 245113
rect 253715 245085 253749 245113
rect 253777 245085 253811 245113
rect 253839 245085 262625 245113
rect 262653 245085 262687 245113
rect 262715 245085 262749 245113
rect 262777 245085 262811 245113
rect 262839 245085 271625 245113
rect 271653 245085 271687 245113
rect 271715 245085 271749 245113
rect 271777 245085 271811 245113
rect 271839 245085 280625 245113
rect 280653 245085 280687 245113
rect 280715 245085 280749 245113
rect 280777 245085 280811 245113
rect 280839 245085 289625 245113
rect 289653 245085 289687 245113
rect 289715 245085 289749 245113
rect 289777 245085 289811 245113
rect 289839 245085 298248 245113
rect 298276 245085 298310 245113
rect 298338 245085 298372 245113
rect 298400 245085 298434 245113
rect 298462 245085 298990 245113
rect -958 245051 298990 245085
rect -958 245023 -430 245051
rect -402 245023 -368 245051
rect -340 245023 -306 245051
rect -278 245023 -244 245051
rect -216 245023 1625 245051
rect 1653 245023 1687 245051
rect 1715 245023 1749 245051
rect 1777 245023 1811 245051
rect 1839 245023 10625 245051
rect 10653 245023 10687 245051
rect 10715 245023 10749 245051
rect 10777 245023 10811 245051
rect 10839 245023 19625 245051
rect 19653 245023 19687 245051
rect 19715 245023 19749 245051
rect 19777 245023 19811 245051
rect 19839 245023 28625 245051
rect 28653 245023 28687 245051
rect 28715 245023 28749 245051
rect 28777 245023 28811 245051
rect 28839 245023 37625 245051
rect 37653 245023 37687 245051
rect 37715 245023 37749 245051
rect 37777 245023 37811 245051
rect 37839 245023 46625 245051
rect 46653 245023 46687 245051
rect 46715 245023 46749 245051
rect 46777 245023 46811 245051
rect 46839 245023 52259 245051
rect 52287 245023 52321 245051
rect 52349 245023 67619 245051
rect 67647 245023 67681 245051
rect 67709 245023 82979 245051
rect 83007 245023 83041 245051
rect 83069 245023 98339 245051
rect 98367 245023 98401 245051
rect 98429 245023 113699 245051
rect 113727 245023 113761 245051
rect 113789 245023 129059 245051
rect 129087 245023 129121 245051
rect 129149 245023 144419 245051
rect 144447 245023 144481 245051
rect 144509 245023 154625 245051
rect 154653 245023 154687 245051
rect 154715 245023 154749 245051
rect 154777 245023 154811 245051
rect 154839 245023 163625 245051
rect 163653 245023 163687 245051
rect 163715 245023 163749 245051
rect 163777 245023 163811 245051
rect 163839 245023 172625 245051
rect 172653 245023 172687 245051
rect 172715 245023 172749 245051
rect 172777 245023 172811 245051
rect 172839 245023 181625 245051
rect 181653 245023 181687 245051
rect 181715 245023 181749 245051
rect 181777 245023 181811 245051
rect 181839 245023 190625 245051
rect 190653 245023 190687 245051
rect 190715 245023 190749 245051
rect 190777 245023 190811 245051
rect 190839 245023 199625 245051
rect 199653 245023 199687 245051
rect 199715 245023 199749 245051
rect 199777 245023 199811 245051
rect 199839 245023 208625 245051
rect 208653 245023 208687 245051
rect 208715 245023 208749 245051
rect 208777 245023 208811 245051
rect 208839 245023 217625 245051
rect 217653 245023 217687 245051
rect 217715 245023 217749 245051
rect 217777 245023 217811 245051
rect 217839 245023 226625 245051
rect 226653 245023 226687 245051
rect 226715 245023 226749 245051
rect 226777 245023 226811 245051
rect 226839 245023 235625 245051
rect 235653 245023 235687 245051
rect 235715 245023 235749 245051
rect 235777 245023 235811 245051
rect 235839 245023 244625 245051
rect 244653 245023 244687 245051
rect 244715 245023 244749 245051
rect 244777 245023 244811 245051
rect 244839 245023 253625 245051
rect 253653 245023 253687 245051
rect 253715 245023 253749 245051
rect 253777 245023 253811 245051
rect 253839 245023 262625 245051
rect 262653 245023 262687 245051
rect 262715 245023 262749 245051
rect 262777 245023 262811 245051
rect 262839 245023 271625 245051
rect 271653 245023 271687 245051
rect 271715 245023 271749 245051
rect 271777 245023 271811 245051
rect 271839 245023 280625 245051
rect 280653 245023 280687 245051
rect 280715 245023 280749 245051
rect 280777 245023 280811 245051
rect 280839 245023 289625 245051
rect 289653 245023 289687 245051
rect 289715 245023 289749 245051
rect 289777 245023 289811 245051
rect 289839 245023 298248 245051
rect 298276 245023 298310 245051
rect 298338 245023 298372 245051
rect 298400 245023 298434 245051
rect 298462 245023 298990 245051
rect -958 244989 298990 245023
rect -958 244961 -430 244989
rect -402 244961 -368 244989
rect -340 244961 -306 244989
rect -278 244961 -244 244989
rect -216 244961 1625 244989
rect 1653 244961 1687 244989
rect 1715 244961 1749 244989
rect 1777 244961 1811 244989
rect 1839 244961 10625 244989
rect 10653 244961 10687 244989
rect 10715 244961 10749 244989
rect 10777 244961 10811 244989
rect 10839 244961 19625 244989
rect 19653 244961 19687 244989
rect 19715 244961 19749 244989
rect 19777 244961 19811 244989
rect 19839 244961 28625 244989
rect 28653 244961 28687 244989
rect 28715 244961 28749 244989
rect 28777 244961 28811 244989
rect 28839 244961 37625 244989
rect 37653 244961 37687 244989
rect 37715 244961 37749 244989
rect 37777 244961 37811 244989
rect 37839 244961 46625 244989
rect 46653 244961 46687 244989
rect 46715 244961 46749 244989
rect 46777 244961 46811 244989
rect 46839 244961 52259 244989
rect 52287 244961 52321 244989
rect 52349 244961 67619 244989
rect 67647 244961 67681 244989
rect 67709 244961 82979 244989
rect 83007 244961 83041 244989
rect 83069 244961 98339 244989
rect 98367 244961 98401 244989
rect 98429 244961 113699 244989
rect 113727 244961 113761 244989
rect 113789 244961 129059 244989
rect 129087 244961 129121 244989
rect 129149 244961 144419 244989
rect 144447 244961 144481 244989
rect 144509 244961 154625 244989
rect 154653 244961 154687 244989
rect 154715 244961 154749 244989
rect 154777 244961 154811 244989
rect 154839 244961 163625 244989
rect 163653 244961 163687 244989
rect 163715 244961 163749 244989
rect 163777 244961 163811 244989
rect 163839 244961 172625 244989
rect 172653 244961 172687 244989
rect 172715 244961 172749 244989
rect 172777 244961 172811 244989
rect 172839 244961 181625 244989
rect 181653 244961 181687 244989
rect 181715 244961 181749 244989
rect 181777 244961 181811 244989
rect 181839 244961 190625 244989
rect 190653 244961 190687 244989
rect 190715 244961 190749 244989
rect 190777 244961 190811 244989
rect 190839 244961 199625 244989
rect 199653 244961 199687 244989
rect 199715 244961 199749 244989
rect 199777 244961 199811 244989
rect 199839 244961 208625 244989
rect 208653 244961 208687 244989
rect 208715 244961 208749 244989
rect 208777 244961 208811 244989
rect 208839 244961 217625 244989
rect 217653 244961 217687 244989
rect 217715 244961 217749 244989
rect 217777 244961 217811 244989
rect 217839 244961 226625 244989
rect 226653 244961 226687 244989
rect 226715 244961 226749 244989
rect 226777 244961 226811 244989
rect 226839 244961 235625 244989
rect 235653 244961 235687 244989
rect 235715 244961 235749 244989
rect 235777 244961 235811 244989
rect 235839 244961 244625 244989
rect 244653 244961 244687 244989
rect 244715 244961 244749 244989
rect 244777 244961 244811 244989
rect 244839 244961 253625 244989
rect 253653 244961 253687 244989
rect 253715 244961 253749 244989
rect 253777 244961 253811 244989
rect 253839 244961 262625 244989
rect 262653 244961 262687 244989
rect 262715 244961 262749 244989
rect 262777 244961 262811 244989
rect 262839 244961 271625 244989
rect 271653 244961 271687 244989
rect 271715 244961 271749 244989
rect 271777 244961 271811 244989
rect 271839 244961 280625 244989
rect 280653 244961 280687 244989
rect 280715 244961 280749 244989
rect 280777 244961 280811 244989
rect 280839 244961 289625 244989
rect 289653 244961 289687 244989
rect 289715 244961 289749 244989
rect 289777 244961 289811 244989
rect 289839 244961 298248 244989
rect 298276 244961 298310 244989
rect 298338 244961 298372 244989
rect 298400 244961 298434 244989
rect 298462 244961 298990 244989
rect -958 244913 298990 244961
rect -958 239175 298990 239223
rect -958 239147 -910 239175
rect -882 239147 -848 239175
rect -820 239147 -786 239175
rect -758 239147 -724 239175
rect -696 239147 3485 239175
rect 3513 239147 3547 239175
rect 3575 239147 3609 239175
rect 3637 239147 3671 239175
rect 3699 239147 12485 239175
rect 12513 239147 12547 239175
rect 12575 239147 12609 239175
rect 12637 239147 12671 239175
rect 12699 239147 21485 239175
rect 21513 239147 21547 239175
rect 21575 239147 21609 239175
rect 21637 239147 21671 239175
rect 21699 239147 30485 239175
rect 30513 239147 30547 239175
rect 30575 239147 30609 239175
rect 30637 239147 30671 239175
rect 30699 239147 39485 239175
rect 39513 239147 39547 239175
rect 39575 239147 39609 239175
rect 39637 239147 39671 239175
rect 39699 239147 48485 239175
rect 48513 239147 48547 239175
rect 48575 239147 48609 239175
rect 48637 239147 48671 239175
rect 48699 239147 59939 239175
rect 59967 239147 60001 239175
rect 60029 239147 75299 239175
rect 75327 239147 75361 239175
rect 75389 239147 90659 239175
rect 90687 239147 90721 239175
rect 90749 239147 106019 239175
rect 106047 239147 106081 239175
rect 106109 239147 121379 239175
rect 121407 239147 121441 239175
rect 121469 239147 136739 239175
rect 136767 239147 136801 239175
rect 136829 239147 156485 239175
rect 156513 239147 156547 239175
rect 156575 239147 156609 239175
rect 156637 239147 156671 239175
rect 156699 239147 165485 239175
rect 165513 239147 165547 239175
rect 165575 239147 165609 239175
rect 165637 239147 165671 239175
rect 165699 239147 174485 239175
rect 174513 239147 174547 239175
rect 174575 239147 174609 239175
rect 174637 239147 174671 239175
rect 174699 239147 183485 239175
rect 183513 239147 183547 239175
rect 183575 239147 183609 239175
rect 183637 239147 183671 239175
rect 183699 239147 192485 239175
rect 192513 239147 192547 239175
rect 192575 239147 192609 239175
rect 192637 239147 192671 239175
rect 192699 239147 201485 239175
rect 201513 239147 201547 239175
rect 201575 239147 201609 239175
rect 201637 239147 201671 239175
rect 201699 239147 210485 239175
rect 210513 239147 210547 239175
rect 210575 239147 210609 239175
rect 210637 239147 210671 239175
rect 210699 239147 219485 239175
rect 219513 239147 219547 239175
rect 219575 239147 219609 239175
rect 219637 239147 219671 239175
rect 219699 239147 228485 239175
rect 228513 239147 228547 239175
rect 228575 239147 228609 239175
rect 228637 239147 228671 239175
rect 228699 239147 237485 239175
rect 237513 239147 237547 239175
rect 237575 239147 237609 239175
rect 237637 239147 237671 239175
rect 237699 239147 246485 239175
rect 246513 239147 246547 239175
rect 246575 239147 246609 239175
rect 246637 239147 246671 239175
rect 246699 239147 255485 239175
rect 255513 239147 255547 239175
rect 255575 239147 255609 239175
rect 255637 239147 255671 239175
rect 255699 239147 264485 239175
rect 264513 239147 264547 239175
rect 264575 239147 264609 239175
rect 264637 239147 264671 239175
rect 264699 239147 273485 239175
rect 273513 239147 273547 239175
rect 273575 239147 273609 239175
rect 273637 239147 273671 239175
rect 273699 239147 282485 239175
rect 282513 239147 282547 239175
rect 282575 239147 282609 239175
rect 282637 239147 282671 239175
rect 282699 239147 291485 239175
rect 291513 239147 291547 239175
rect 291575 239147 291609 239175
rect 291637 239147 291671 239175
rect 291699 239147 298728 239175
rect 298756 239147 298790 239175
rect 298818 239147 298852 239175
rect 298880 239147 298914 239175
rect 298942 239147 298990 239175
rect -958 239113 298990 239147
rect -958 239085 -910 239113
rect -882 239085 -848 239113
rect -820 239085 -786 239113
rect -758 239085 -724 239113
rect -696 239085 3485 239113
rect 3513 239085 3547 239113
rect 3575 239085 3609 239113
rect 3637 239085 3671 239113
rect 3699 239085 12485 239113
rect 12513 239085 12547 239113
rect 12575 239085 12609 239113
rect 12637 239085 12671 239113
rect 12699 239085 21485 239113
rect 21513 239085 21547 239113
rect 21575 239085 21609 239113
rect 21637 239085 21671 239113
rect 21699 239085 30485 239113
rect 30513 239085 30547 239113
rect 30575 239085 30609 239113
rect 30637 239085 30671 239113
rect 30699 239085 39485 239113
rect 39513 239085 39547 239113
rect 39575 239085 39609 239113
rect 39637 239085 39671 239113
rect 39699 239085 48485 239113
rect 48513 239085 48547 239113
rect 48575 239085 48609 239113
rect 48637 239085 48671 239113
rect 48699 239085 59939 239113
rect 59967 239085 60001 239113
rect 60029 239085 75299 239113
rect 75327 239085 75361 239113
rect 75389 239085 90659 239113
rect 90687 239085 90721 239113
rect 90749 239085 106019 239113
rect 106047 239085 106081 239113
rect 106109 239085 121379 239113
rect 121407 239085 121441 239113
rect 121469 239085 136739 239113
rect 136767 239085 136801 239113
rect 136829 239085 156485 239113
rect 156513 239085 156547 239113
rect 156575 239085 156609 239113
rect 156637 239085 156671 239113
rect 156699 239085 165485 239113
rect 165513 239085 165547 239113
rect 165575 239085 165609 239113
rect 165637 239085 165671 239113
rect 165699 239085 174485 239113
rect 174513 239085 174547 239113
rect 174575 239085 174609 239113
rect 174637 239085 174671 239113
rect 174699 239085 183485 239113
rect 183513 239085 183547 239113
rect 183575 239085 183609 239113
rect 183637 239085 183671 239113
rect 183699 239085 192485 239113
rect 192513 239085 192547 239113
rect 192575 239085 192609 239113
rect 192637 239085 192671 239113
rect 192699 239085 201485 239113
rect 201513 239085 201547 239113
rect 201575 239085 201609 239113
rect 201637 239085 201671 239113
rect 201699 239085 210485 239113
rect 210513 239085 210547 239113
rect 210575 239085 210609 239113
rect 210637 239085 210671 239113
rect 210699 239085 219485 239113
rect 219513 239085 219547 239113
rect 219575 239085 219609 239113
rect 219637 239085 219671 239113
rect 219699 239085 228485 239113
rect 228513 239085 228547 239113
rect 228575 239085 228609 239113
rect 228637 239085 228671 239113
rect 228699 239085 237485 239113
rect 237513 239085 237547 239113
rect 237575 239085 237609 239113
rect 237637 239085 237671 239113
rect 237699 239085 246485 239113
rect 246513 239085 246547 239113
rect 246575 239085 246609 239113
rect 246637 239085 246671 239113
rect 246699 239085 255485 239113
rect 255513 239085 255547 239113
rect 255575 239085 255609 239113
rect 255637 239085 255671 239113
rect 255699 239085 264485 239113
rect 264513 239085 264547 239113
rect 264575 239085 264609 239113
rect 264637 239085 264671 239113
rect 264699 239085 273485 239113
rect 273513 239085 273547 239113
rect 273575 239085 273609 239113
rect 273637 239085 273671 239113
rect 273699 239085 282485 239113
rect 282513 239085 282547 239113
rect 282575 239085 282609 239113
rect 282637 239085 282671 239113
rect 282699 239085 291485 239113
rect 291513 239085 291547 239113
rect 291575 239085 291609 239113
rect 291637 239085 291671 239113
rect 291699 239085 298728 239113
rect 298756 239085 298790 239113
rect 298818 239085 298852 239113
rect 298880 239085 298914 239113
rect 298942 239085 298990 239113
rect -958 239051 298990 239085
rect -958 239023 -910 239051
rect -882 239023 -848 239051
rect -820 239023 -786 239051
rect -758 239023 -724 239051
rect -696 239023 3485 239051
rect 3513 239023 3547 239051
rect 3575 239023 3609 239051
rect 3637 239023 3671 239051
rect 3699 239023 12485 239051
rect 12513 239023 12547 239051
rect 12575 239023 12609 239051
rect 12637 239023 12671 239051
rect 12699 239023 21485 239051
rect 21513 239023 21547 239051
rect 21575 239023 21609 239051
rect 21637 239023 21671 239051
rect 21699 239023 30485 239051
rect 30513 239023 30547 239051
rect 30575 239023 30609 239051
rect 30637 239023 30671 239051
rect 30699 239023 39485 239051
rect 39513 239023 39547 239051
rect 39575 239023 39609 239051
rect 39637 239023 39671 239051
rect 39699 239023 48485 239051
rect 48513 239023 48547 239051
rect 48575 239023 48609 239051
rect 48637 239023 48671 239051
rect 48699 239023 59939 239051
rect 59967 239023 60001 239051
rect 60029 239023 75299 239051
rect 75327 239023 75361 239051
rect 75389 239023 90659 239051
rect 90687 239023 90721 239051
rect 90749 239023 106019 239051
rect 106047 239023 106081 239051
rect 106109 239023 121379 239051
rect 121407 239023 121441 239051
rect 121469 239023 136739 239051
rect 136767 239023 136801 239051
rect 136829 239023 156485 239051
rect 156513 239023 156547 239051
rect 156575 239023 156609 239051
rect 156637 239023 156671 239051
rect 156699 239023 165485 239051
rect 165513 239023 165547 239051
rect 165575 239023 165609 239051
rect 165637 239023 165671 239051
rect 165699 239023 174485 239051
rect 174513 239023 174547 239051
rect 174575 239023 174609 239051
rect 174637 239023 174671 239051
rect 174699 239023 183485 239051
rect 183513 239023 183547 239051
rect 183575 239023 183609 239051
rect 183637 239023 183671 239051
rect 183699 239023 192485 239051
rect 192513 239023 192547 239051
rect 192575 239023 192609 239051
rect 192637 239023 192671 239051
rect 192699 239023 201485 239051
rect 201513 239023 201547 239051
rect 201575 239023 201609 239051
rect 201637 239023 201671 239051
rect 201699 239023 210485 239051
rect 210513 239023 210547 239051
rect 210575 239023 210609 239051
rect 210637 239023 210671 239051
rect 210699 239023 219485 239051
rect 219513 239023 219547 239051
rect 219575 239023 219609 239051
rect 219637 239023 219671 239051
rect 219699 239023 228485 239051
rect 228513 239023 228547 239051
rect 228575 239023 228609 239051
rect 228637 239023 228671 239051
rect 228699 239023 237485 239051
rect 237513 239023 237547 239051
rect 237575 239023 237609 239051
rect 237637 239023 237671 239051
rect 237699 239023 246485 239051
rect 246513 239023 246547 239051
rect 246575 239023 246609 239051
rect 246637 239023 246671 239051
rect 246699 239023 255485 239051
rect 255513 239023 255547 239051
rect 255575 239023 255609 239051
rect 255637 239023 255671 239051
rect 255699 239023 264485 239051
rect 264513 239023 264547 239051
rect 264575 239023 264609 239051
rect 264637 239023 264671 239051
rect 264699 239023 273485 239051
rect 273513 239023 273547 239051
rect 273575 239023 273609 239051
rect 273637 239023 273671 239051
rect 273699 239023 282485 239051
rect 282513 239023 282547 239051
rect 282575 239023 282609 239051
rect 282637 239023 282671 239051
rect 282699 239023 291485 239051
rect 291513 239023 291547 239051
rect 291575 239023 291609 239051
rect 291637 239023 291671 239051
rect 291699 239023 298728 239051
rect 298756 239023 298790 239051
rect 298818 239023 298852 239051
rect 298880 239023 298914 239051
rect 298942 239023 298990 239051
rect -958 238989 298990 239023
rect -958 238961 -910 238989
rect -882 238961 -848 238989
rect -820 238961 -786 238989
rect -758 238961 -724 238989
rect -696 238961 3485 238989
rect 3513 238961 3547 238989
rect 3575 238961 3609 238989
rect 3637 238961 3671 238989
rect 3699 238961 12485 238989
rect 12513 238961 12547 238989
rect 12575 238961 12609 238989
rect 12637 238961 12671 238989
rect 12699 238961 21485 238989
rect 21513 238961 21547 238989
rect 21575 238961 21609 238989
rect 21637 238961 21671 238989
rect 21699 238961 30485 238989
rect 30513 238961 30547 238989
rect 30575 238961 30609 238989
rect 30637 238961 30671 238989
rect 30699 238961 39485 238989
rect 39513 238961 39547 238989
rect 39575 238961 39609 238989
rect 39637 238961 39671 238989
rect 39699 238961 48485 238989
rect 48513 238961 48547 238989
rect 48575 238961 48609 238989
rect 48637 238961 48671 238989
rect 48699 238961 59939 238989
rect 59967 238961 60001 238989
rect 60029 238961 75299 238989
rect 75327 238961 75361 238989
rect 75389 238961 90659 238989
rect 90687 238961 90721 238989
rect 90749 238961 106019 238989
rect 106047 238961 106081 238989
rect 106109 238961 121379 238989
rect 121407 238961 121441 238989
rect 121469 238961 136739 238989
rect 136767 238961 136801 238989
rect 136829 238961 156485 238989
rect 156513 238961 156547 238989
rect 156575 238961 156609 238989
rect 156637 238961 156671 238989
rect 156699 238961 165485 238989
rect 165513 238961 165547 238989
rect 165575 238961 165609 238989
rect 165637 238961 165671 238989
rect 165699 238961 174485 238989
rect 174513 238961 174547 238989
rect 174575 238961 174609 238989
rect 174637 238961 174671 238989
rect 174699 238961 183485 238989
rect 183513 238961 183547 238989
rect 183575 238961 183609 238989
rect 183637 238961 183671 238989
rect 183699 238961 192485 238989
rect 192513 238961 192547 238989
rect 192575 238961 192609 238989
rect 192637 238961 192671 238989
rect 192699 238961 201485 238989
rect 201513 238961 201547 238989
rect 201575 238961 201609 238989
rect 201637 238961 201671 238989
rect 201699 238961 210485 238989
rect 210513 238961 210547 238989
rect 210575 238961 210609 238989
rect 210637 238961 210671 238989
rect 210699 238961 219485 238989
rect 219513 238961 219547 238989
rect 219575 238961 219609 238989
rect 219637 238961 219671 238989
rect 219699 238961 228485 238989
rect 228513 238961 228547 238989
rect 228575 238961 228609 238989
rect 228637 238961 228671 238989
rect 228699 238961 237485 238989
rect 237513 238961 237547 238989
rect 237575 238961 237609 238989
rect 237637 238961 237671 238989
rect 237699 238961 246485 238989
rect 246513 238961 246547 238989
rect 246575 238961 246609 238989
rect 246637 238961 246671 238989
rect 246699 238961 255485 238989
rect 255513 238961 255547 238989
rect 255575 238961 255609 238989
rect 255637 238961 255671 238989
rect 255699 238961 264485 238989
rect 264513 238961 264547 238989
rect 264575 238961 264609 238989
rect 264637 238961 264671 238989
rect 264699 238961 273485 238989
rect 273513 238961 273547 238989
rect 273575 238961 273609 238989
rect 273637 238961 273671 238989
rect 273699 238961 282485 238989
rect 282513 238961 282547 238989
rect 282575 238961 282609 238989
rect 282637 238961 282671 238989
rect 282699 238961 291485 238989
rect 291513 238961 291547 238989
rect 291575 238961 291609 238989
rect 291637 238961 291671 238989
rect 291699 238961 298728 238989
rect 298756 238961 298790 238989
rect 298818 238961 298852 238989
rect 298880 238961 298914 238989
rect 298942 238961 298990 238989
rect -958 238913 298990 238961
rect -958 236175 298990 236223
rect -958 236147 -430 236175
rect -402 236147 -368 236175
rect -340 236147 -306 236175
rect -278 236147 -244 236175
rect -216 236147 1625 236175
rect 1653 236147 1687 236175
rect 1715 236147 1749 236175
rect 1777 236147 1811 236175
rect 1839 236147 10625 236175
rect 10653 236147 10687 236175
rect 10715 236147 10749 236175
rect 10777 236147 10811 236175
rect 10839 236147 19625 236175
rect 19653 236147 19687 236175
rect 19715 236147 19749 236175
rect 19777 236147 19811 236175
rect 19839 236147 28625 236175
rect 28653 236147 28687 236175
rect 28715 236147 28749 236175
rect 28777 236147 28811 236175
rect 28839 236147 37625 236175
rect 37653 236147 37687 236175
rect 37715 236147 37749 236175
rect 37777 236147 37811 236175
rect 37839 236147 46625 236175
rect 46653 236147 46687 236175
rect 46715 236147 46749 236175
rect 46777 236147 46811 236175
rect 46839 236147 52259 236175
rect 52287 236147 52321 236175
rect 52349 236147 67619 236175
rect 67647 236147 67681 236175
rect 67709 236147 82979 236175
rect 83007 236147 83041 236175
rect 83069 236147 98339 236175
rect 98367 236147 98401 236175
rect 98429 236147 113699 236175
rect 113727 236147 113761 236175
rect 113789 236147 129059 236175
rect 129087 236147 129121 236175
rect 129149 236147 144419 236175
rect 144447 236147 144481 236175
rect 144509 236147 154625 236175
rect 154653 236147 154687 236175
rect 154715 236147 154749 236175
rect 154777 236147 154811 236175
rect 154839 236147 163625 236175
rect 163653 236147 163687 236175
rect 163715 236147 163749 236175
rect 163777 236147 163811 236175
rect 163839 236147 172625 236175
rect 172653 236147 172687 236175
rect 172715 236147 172749 236175
rect 172777 236147 172811 236175
rect 172839 236147 181625 236175
rect 181653 236147 181687 236175
rect 181715 236147 181749 236175
rect 181777 236147 181811 236175
rect 181839 236147 190625 236175
rect 190653 236147 190687 236175
rect 190715 236147 190749 236175
rect 190777 236147 190811 236175
rect 190839 236147 199625 236175
rect 199653 236147 199687 236175
rect 199715 236147 199749 236175
rect 199777 236147 199811 236175
rect 199839 236147 208625 236175
rect 208653 236147 208687 236175
rect 208715 236147 208749 236175
rect 208777 236147 208811 236175
rect 208839 236147 217625 236175
rect 217653 236147 217687 236175
rect 217715 236147 217749 236175
rect 217777 236147 217811 236175
rect 217839 236147 226625 236175
rect 226653 236147 226687 236175
rect 226715 236147 226749 236175
rect 226777 236147 226811 236175
rect 226839 236147 235625 236175
rect 235653 236147 235687 236175
rect 235715 236147 235749 236175
rect 235777 236147 235811 236175
rect 235839 236147 244625 236175
rect 244653 236147 244687 236175
rect 244715 236147 244749 236175
rect 244777 236147 244811 236175
rect 244839 236147 253625 236175
rect 253653 236147 253687 236175
rect 253715 236147 253749 236175
rect 253777 236147 253811 236175
rect 253839 236147 262625 236175
rect 262653 236147 262687 236175
rect 262715 236147 262749 236175
rect 262777 236147 262811 236175
rect 262839 236147 271625 236175
rect 271653 236147 271687 236175
rect 271715 236147 271749 236175
rect 271777 236147 271811 236175
rect 271839 236147 280625 236175
rect 280653 236147 280687 236175
rect 280715 236147 280749 236175
rect 280777 236147 280811 236175
rect 280839 236147 289625 236175
rect 289653 236147 289687 236175
rect 289715 236147 289749 236175
rect 289777 236147 289811 236175
rect 289839 236147 298248 236175
rect 298276 236147 298310 236175
rect 298338 236147 298372 236175
rect 298400 236147 298434 236175
rect 298462 236147 298990 236175
rect -958 236113 298990 236147
rect -958 236085 -430 236113
rect -402 236085 -368 236113
rect -340 236085 -306 236113
rect -278 236085 -244 236113
rect -216 236085 1625 236113
rect 1653 236085 1687 236113
rect 1715 236085 1749 236113
rect 1777 236085 1811 236113
rect 1839 236085 10625 236113
rect 10653 236085 10687 236113
rect 10715 236085 10749 236113
rect 10777 236085 10811 236113
rect 10839 236085 19625 236113
rect 19653 236085 19687 236113
rect 19715 236085 19749 236113
rect 19777 236085 19811 236113
rect 19839 236085 28625 236113
rect 28653 236085 28687 236113
rect 28715 236085 28749 236113
rect 28777 236085 28811 236113
rect 28839 236085 37625 236113
rect 37653 236085 37687 236113
rect 37715 236085 37749 236113
rect 37777 236085 37811 236113
rect 37839 236085 46625 236113
rect 46653 236085 46687 236113
rect 46715 236085 46749 236113
rect 46777 236085 46811 236113
rect 46839 236085 52259 236113
rect 52287 236085 52321 236113
rect 52349 236085 67619 236113
rect 67647 236085 67681 236113
rect 67709 236085 82979 236113
rect 83007 236085 83041 236113
rect 83069 236085 98339 236113
rect 98367 236085 98401 236113
rect 98429 236085 113699 236113
rect 113727 236085 113761 236113
rect 113789 236085 129059 236113
rect 129087 236085 129121 236113
rect 129149 236085 144419 236113
rect 144447 236085 144481 236113
rect 144509 236085 154625 236113
rect 154653 236085 154687 236113
rect 154715 236085 154749 236113
rect 154777 236085 154811 236113
rect 154839 236085 163625 236113
rect 163653 236085 163687 236113
rect 163715 236085 163749 236113
rect 163777 236085 163811 236113
rect 163839 236085 172625 236113
rect 172653 236085 172687 236113
rect 172715 236085 172749 236113
rect 172777 236085 172811 236113
rect 172839 236085 181625 236113
rect 181653 236085 181687 236113
rect 181715 236085 181749 236113
rect 181777 236085 181811 236113
rect 181839 236085 190625 236113
rect 190653 236085 190687 236113
rect 190715 236085 190749 236113
rect 190777 236085 190811 236113
rect 190839 236085 199625 236113
rect 199653 236085 199687 236113
rect 199715 236085 199749 236113
rect 199777 236085 199811 236113
rect 199839 236085 208625 236113
rect 208653 236085 208687 236113
rect 208715 236085 208749 236113
rect 208777 236085 208811 236113
rect 208839 236085 217625 236113
rect 217653 236085 217687 236113
rect 217715 236085 217749 236113
rect 217777 236085 217811 236113
rect 217839 236085 226625 236113
rect 226653 236085 226687 236113
rect 226715 236085 226749 236113
rect 226777 236085 226811 236113
rect 226839 236085 235625 236113
rect 235653 236085 235687 236113
rect 235715 236085 235749 236113
rect 235777 236085 235811 236113
rect 235839 236085 244625 236113
rect 244653 236085 244687 236113
rect 244715 236085 244749 236113
rect 244777 236085 244811 236113
rect 244839 236085 253625 236113
rect 253653 236085 253687 236113
rect 253715 236085 253749 236113
rect 253777 236085 253811 236113
rect 253839 236085 262625 236113
rect 262653 236085 262687 236113
rect 262715 236085 262749 236113
rect 262777 236085 262811 236113
rect 262839 236085 271625 236113
rect 271653 236085 271687 236113
rect 271715 236085 271749 236113
rect 271777 236085 271811 236113
rect 271839 236085 280625 236113
rect 280653 236085 280687 236113
rect 280715 236085 280749 236113
rect 280777 236085 280811 236113
rect 280839 236085 289625 236113
rect 289653 236085 289687 236113
rect 289715 236085 289749 236113
rect 289777 236085 289811 236113
rect 289839 236085 298248 236113
rect 298276 236085 298310 236113
rect 298338 236085 298372 236113
rect 298400 236085 298434 236113
rect 298462 236085 298990 236113
rect -958 236051 298990 236085
rect -958 236023 -430 236051
rect -402 236023 -368 236051
rect -340 236023 -306 236051
rect -278 236023 -244 236051
rect -216 236023 1625 236051
rect 1653 236023 1687 236051
rect 1715 236023 1749 236051
rect 1777 236023 1811 236051
rect 1839 236023 10625 236051
rect 10653 236023 10687 236051
rect 10715 236023 10749 236051
rect 10777 236023 10811 236051
rect 10839 236023 19625 236051
rect 19653 236023 19687 236051
rect 19715 236023 19749 236051
rect 19777 236023 19811 236051
rect 19839 236023 28625 236051
rect 28653 236023 28687 236051
rect 28715 236023 28749 236051
rect 28777 236023 28811 236051
rect 28839 236023 37625 236051
rect 37653 236023 37687 236051
rect 37715 236023 37749 236051
rect 37777 236023 37811 236051
rect 37839 236023 46625 236051
rect 46653 236023 46687 236051
rect 46715 236023 46749 236051
rect 46777 236023 46811 236051
rect 46839 236023 52259 236051
rect 52287 236023 52321 236051
rect 52349 236023 67619 236051
rect 67647 236023 67681 236051
rect 67709 236023 82979 236051
rect 83007 236023 83041 236051
rect 83069 236023 98339 236051
rect 98367 236023 98401 236051
rect 98429 236023 113699 236051
rect 113727 236023 113761 236051
rect 113789 236023 129059 236051
rect 129087 236023 129121 236051
rect 129149 236023 144419 236051
rect 144447 236023 144481 236051
rect 144509 236023 154625 236051
rect 154653 236023 154687 236051
rect 154715 236023 154749 236051
rect 154777 236023 154811 236051
rect 154839 236023 163625 236051
rect 163653 236023 163687 236051
rect 163715 236023 163749 236051
rect 163777 236023 163811 236051
rect 163839 236023 172625 236051
rect 172653 236023 172687 236051
rect 172715 236023 172749 236051
rect 172777 236023 172811 236051
rect 172839 236023 181625 236051
rect 181653 236023 181687 236051
rect 181715 236023 181749 236051
rect 181777 236023 181811 236051
rect 181839 236023 190625 236051
rect 190653 236023 190687 236051
rect 190715 236023 190749 236051
rect 190777 236023 190811 236051
rect 190839 236023 199625 236051
rect 199653 236023 199687 236051
rect 199715 236023 199749 236051
rect 199777 236023 199811 236051
rect 199839 236023 208625 236051
rect 208653 236023 208687 236051
rect 208715 236023 208749 236051
rect 208777 236023 208811 236051
rect 208839 236023 217625 236051
rect 217653 236023 217687 236051
rect 217715 236023 217749 236051
rect 217777 236023 217811 236051
rect 217839 236023 226625 236051
rect 226653 236023 226687 236051
rect 226715 236023 226749 236051
rect 226777 236023 226811 236051
rect 226839 236023 235625 236051
rect 235653 236023 235687 236051
rect 235715 236023 235749 236051
rect 235777 236023 235811 236051
rect 235839 236023 244625 236051
rect 244653 236023 244687 236051
rect 244715 236023 244749 236051
rect 244777 236023 244811 236051
rect 244839 236023 253625 236051
rect 253653 236023 253687 236051
rect 253715 236023 253749 236051
rect 253777 236023 253811 236051
rect 253839 236023 262625 236051
rect 262653 236023 262687 236051
rect 262715 236023 262749 236051
rect 262777 236023 262811 236051
rect 262839 236023 271625 236051
rect 271653 236023 271687 236051
rect 271715 236023 271749 236051
rect 271777 236023 271811 236051
rect 271839 236023 280625 236051
rect 280653 236023 280687 236051
rect 280715 236023 280749 236051
rect 280777 236023 280811 236051
rect 280839 236023 289625 236051
rect 289653 236023 289687 236051
rect 289715 236023 289749 236051
rect 289777 236023 289811 236051
rect 289839 236023 298248 236051
rect 298276 236023 298310 236051
rect 298338 236023 298372 236051
rect 298400 236023 298434 236051
rect 298462 236023 298990 236051
rect -958 235989 298990 236023
rect -958 235961 -430 235989
rect -402 235961 -368 235989
rect -340 235961 -306 235989
rect -278 235961 -244 235989
rect -216 235961 1625 235989
rect 1653 235961 1687 235989
rect 1715 235961 1749 235989
rect 1777 235961 1811 235989
rect 1839 235961 10625 235989
rect 10653 235961 10687 235989
rect 10715 235961 10749 235989
rect 10777 235961 10811 235989
rect 10839 235961 19625 235989
rect 19653 235961 19687 235989
rect 19715 235961 19749 235989
rect 19777 235961 19811 235989
rect 19839 235961 28625 235989
rect 28653 235961 28687 235989
rect 28715 235961 28749 235989
rect 28777 235961 28811 235989
rect 28839 235961 37625 235989
rect 37653 235961 37687 235989
rect 37715 235961 37749 235989
rect 37777 235961 37811 235989
rect 37839 235961 46625 235989
rect 46653 235961 46687 235989
rect 46715 235961 46749 235989
rect 46777 235961 46811 235989
rect 46839 235961 52259 235989
rect 52287 235961 52321 235989
rect 52349 235961 67619 235989
rect 67647 235961 67681 235989
rect 67709 235961 82979 235989
rect 83007 235961 83041 235989
rect 83069 235961 98339 235989
rect 98367 235961 98401 235989
rect 98429 235961 113699 235989
rect 113727 235961 113761 235989
rect 113789 235961 129059 235989
rect 129087 235961 129121 235989
rect 129149 235961 144419 235989
rect 144447 235961 144481 235989
rect 144509 235961 154625 235989
rect 154653 235961 154687 235989
rect 154715 235961 154749 235989
rect 154777 235961 154811 235989
rect 154839 235961 163625 235989
rect 163653 235961 163687 235989
rect 163715 235961 163749 235989
rect 163777 235961 163811 235989
rect 163839 235961 172625 235989
rect 172653 235961 172687 235989
rect 172715 235961 172749 235989
rect 172777 235961 172811 235989
rect 172839 235961 181625 235989
rect 181653 235961 181687 235989
rect 181715 235961 181749 235989
rect 181777 235961 181811 235989
rect 181839 235961 190625 235989
rect 190653 235961 190687 235989
rect 190715 235961 190749 235989
rect 190777 235961 190811 235989
rect 190839 235961 199625 235989
rect 199653 235961 199687 235989
rect 199715 235961 199749 235989
rect 199777 235961 199811 235989
rect 199839 235961 208625 235989
rect 208653 235961 208687 235989
rect 208715 235961 208749 235989
rect 208777 235961 208811 235989
rect 208839 235961 217625 235989
rect 217653 235961 217687 235989
rect 217715 235961 217749 235989
rect 217777 235961 217811 235989
rect 217839 235961 226625 235989
rect 226653 235961 226687 235989
rect 226715 235961 226749 235989
rect 226777 235961 226811 235989
rect 226839 235961 235625 235989
rect 235653 235961 235687 235989
rect 235715 235961 235749 235989
rect 235777 235961 235811 235989
rect 235839 235961 244625 235989
rect 244653 235961 244687 235989
rect 244715 235961 244749 235989
rect 244777 235961 244811 235989
rect 244839 235961 253625 235989
rect 253653 235961 253687 235989
rect 253715 235961 253749 235989
rect 253777 235961 253811 235989
rect 253839 235961 262625 235989
rect 262653 235961 262687 235989
rect 262715 235961 262749 235989
rect 262777 235961 262811 235989
rect 262839 235961 271625 235989
rect 271653 235961 271687 235989
rect 271715 235961 271749 235989
rect 271777 235961 271811 235989
rect 271839 235961 280625 235989
rect 280653 235961 280687 235989
rect 280715 235961 280749 235989
rect 280777 235961 280811 235989
rect 280839 235961 289625 235989
rect 289653 235961 289687 235989
rect 289715 235961 289749 235989
rect 289777 235961 289811 235989
rect 289839 235961 298248 235989
rect 298276 235961 298310 235989
rect 298338 235961 298372 235989
rect 298400 235961 298434 235989
rect 298462 235961 298990 235989
rect -958 235913 298990 235961
rect -958 230175 298990 230223
rect -958 230147 -910 230175
rect -882 230147 -848 230175
rect -820 230147 -786 230175
rect -758 230147 -724 230175
rect -696 230147 3485 230175
rect 3513 230147 3547 230175
rect 3575 230147 3609 230175
rect 3637 230147 3671 230175
rect 3699 230147 12485 230175
rect 12513 230147 12547 230175
rect 12575 230147 12609 230175
rect 12637 230147 12671 230175
rect 12699 230147 21485 230175
rect 21513 230147 21547 230175
rect 21575 230147 21609 230175
rect 21637 230147 21671 230175
rect 21699 230147 30485 230175
rect 30513 230147 30547 230175
rect 30575 230147 30609 230175
rect 30637 230147 30671 230175
rect 30699 230147 39485 230175
rect 39513 230147 39547 230175
rect 39575 230147 39609 230175
rect 39637 230147 39671 230175
rect 39699 230147 48485 230175
rect 48513 230147 48547 230175
rect 48575 230147 48609 230175
rect 48637 230147 48671 230175
rect 48699 230147 59939 230175
rect 59967 230147 60001 230175
rect 60029 230147 75299 230175
rect 75327 230147 75361 230175
rect 75389 230147 90659 230175
rect 90687 230147 90721 230175
rect 90749 230147 106019 230175
rect 106047 230147 106081 230175
rect 106109 230147 121379 230175
rect 121407 230147 121441 230175
rect 121469 230147 136739 230175
rect 136767 230147 136801 230175
rect 136829 230147 156485 230175
rect 156513 230147 156547 230175
rect 156575 230147 156609 230175
rect 156637 230147 156671 230175
rect 156699 230147 165485 230175
rect 165513 230147 165547 230175
rect 165575 230147 165609 230175
rect 165637 230147 165671 230175
rect 165699 230147 174485 230175
rect 174513 230147 174547 230175
rect 174575 230147 174609 230175
rect 174637 230147 174671 230175
rect 174699 230147 183485 230175
rect 183513 230147 183547 230175
rect 183575 230147 183609 230175
rect 183637 230147 183671 230175
rect 183699 230147 192485 230175
rect 192513 230147 192547 230175
rect 192575 230147 192609 230175
rect 192637 230147 192671 230175
rect 192699 230147 201485 230175
rect 201513 230147 201547 230175
rect 201575 230147 201609 230175
rect 201637 230147 201671 230175
rect 201699 230147 210485 230175
rect 210513 230147 210547 230175
rect 210575 230147 210609 230175
rect 210637 230147 210671 230175
rect 210699 230147 219485 230175
rect 219513 230147 219547 230175
rect 219575 230147 219609 230175
rect 219637 230147 219671 230175
rect 219699 230147 228485 230175
rect 228513 230147 228547 230175
rect 228575 230147 228609 230175
rect 228637 230147 228671 230175
rect 228699 230147 237485 230175
rect 237513 230147 237547 230175
rect 237575 230147 237609 230175
rect 237637 230147 237671 230175
rect 237699 230147 246485 230175
rect 246513 230147 246547 230175
rect 246575 230147 246609 230175
rect 246637 230147 246671 230175
rect 246699 230147 255485 230175
rect 255513 230147 255547 230175
rect 255575 230147 255609 230175
rect 255637 230147 255671 230175
rect 255699 230147 264485 230175
rect 264513 230147 264547 230175
rect 264575 230147 264609 230175
rect 264637 230147 264671 230175
rect 264699 230147 273485 230175
rect 273513 230147 273547 230175
rect 273575 230147 273609 230175
rect 273637 230147 273671 230175
rect 273699 230147 282485 230175
rect 282513 230147 282547 230175
rect 282575 230147 282609 230175
rect 282637 230147 282671 230175
rect 282699 230147 291485 230175
rect 291513 230147 291547 230175
rect 291575 230147 291609 230175
rect 291637 230147 291671 230175
rect 291699 230147 298728 230175
rect 298756 230147 298790 230175
rect 298818 230147 298852 230175
rect 298880 230147 298914 230175
rect 298942 230147 298990 230175
rect -958 230113 298990 230147
rect -958 230085 -910 230113
rect -882 230085 -848 230113
rect -820 230085 -786 230113
rect -758 230085 -724 230113
rect -696 230085 3485 230113
rect 3513 230085 3547 230113
rect 3575 230085 3609 230113
rect 3637 230085 3671 230113
rect 3699 230085 12485 230113
rect 12513 230085 12547 230113
rect 12575 230085 12609 230113
rect 12637 230085 12671 230113
rect 12699 230085 21485 230113
rect 21513 230085 21547 230113
rect 21575 230085 21609 230113
rect 21637 230085 21671 230113
rect 21699 230085 30485 230113
rect 30513 230085 30547 230113
rect 30575 230085 30609 230113
rect 30637 230085 30671 230113
rect 30699 230085 39485 230113
rect 39513 230085 39547 230113
rect 39575 230085 39609 230113
rect 39637 230085 39671 230113
rect 39699 230085 48485 230113
rect 48513 230085 48547 230113
rect 48575 230085 48609 230113
rect 48637 230085 48671 230113
rect 48699 230085 59939 230113
rect 59967 230085 60001 230113
rect 60029 230085 75299 230113
rect 75327 230085 75361 230113
rect 75389 230085 90659 230113
rect 90687 230085 90721 230113
rect 90749 230085 106019 230113
rect 106047 230085 106081 230113
rect 106109 230085 121379 230113
rect 121407 230085 121441 230113
rect 121469 230085 136739 230113
rect 136767 230085 136801 230113
rect 136829 230085 156485 230113
rect 156513 230085 156547 230113
rect 156575 230085 156609 230113
rect 156637 230085 156671 230113
rect 156699 230085 165485 230113
rect 165513 230085 165547 230113
rect 165575 230085 165609 230113
rect 165637 230085 165671 230113
rect 165699 230085 174485 230113
rect 174513 230085 174547 230113
rect 174575 230085 174609 230113
rect 174637 230085 174671 230113
rect 174699 230085 183485 230113
rect 183513 230085 183547 230113
rect 183575 230085 183609 230113
rect 183637 230085 183671 230113
rect 183699 230085 192485 230113
rect 192513 230085 192547 230113
rect 192575 230085 192609 230113
rect 192637 230085 192671 230113
rect 192699 230085 201485 230113
rect 201513 230085 201547 230113
rect 201575 230085 201609 230113
rect 201637 230085 201671 230113
rect 201699 230085 210485 230113
rect 210513 230085 210547 230113
rect 210575 230085 210609 230113
rect 210637 230085 210671 230113
rect 210699 230085 219485 230113
rect 219513 230085 219547 230113
rect 219575 230085 219609 230113
rect 219637 230085 219671 230113
rect 219699 230085 228485 230113
rect 228513 230085 228547 230113
rect 228575 230085 228609 230113
rect 228637 230085 228671 230113
rect 228699 230085 237485 230113
rect 237513 230085 237547 230113
rect 237575 230085 237609 230113
rect 237637 230085 237671 230113
rect 237699 230085 246485 230113
rect 246513 230085 246547 230113
rect 246575 230085 246609 230113
rect 246637 230085 246671 230113
rect 246699 230085 255485 230113
rect 255513 230085 255547 230113
rect 255575 230085 255609 230113
rect 255637 230085 255671 230113
rect 255699 230085 264485 230113
rect 264513 230085 264547 230113
rect 264575 230085 264609 230113
rect 264637 230085 264671 230113
rect 264699 230085 273485 230113
rect 273513 230085 273547 230113
rect 273575 230085 273609 230113
rect 273637 230085 273671 230113
rect 273699 230085 282485 230113
rect 282513 230085 282547 230113
rect 282575 230085 282609 230113
rect 282637 230085 282671 230113
rect 282699 230085 291485 230113
rect 291513 230085 291547 230113
rect 291575 230085 291609 230113
rect 291637 230085 291671 230113
rect 291699 230085 298728 230113
rect 298756 230085 298790 230113
rect 298818 230085 298852 230113
rect 298880 230085 298914 230113
rect 298942 230085 298990 230113
rect -958 230051 298990 230085
rect -958 230023 -910 230051
rect -882 230023 -848 230051
rect -820 230023 -786 230051
rect -758 230023 -724 230051
rect -696 230023 3485 230051
rect 3513 230023 3547 230051
rect 3575 230023 3609 230051
rect 3637 230023 3671 230051
rect 3699 230023 12485 230051
rect 12513 230023 12547 230051
rect 12575 230023 12609 230051
rect 12637 230023 12671 230051
rect 12699 230023 21485 230051
rect 21513 230023 21547 230051
rect 21575 230023 21609 230051
rect 21637 230023 21671 230051
rect 21699 230023 30485 230051
rect 30513 230023 30547 230051
rect 30575 230023 30609 230051
rect 30637 230023 30671 230051
rect 30699 230023 39485 230051
rect 39513 230023 39547 230051
rect 39575 230023 39609 230051
rect 39637 230023 39671 230051
rect 39699 230023 48485 230051
rect 48513 230023 48547 230051
rect 48575 230023 48609 230051
rect 48637 230023 48671 230051
rect 48699 230023 59939 230051
rect 59967 230023 60001 230051
rect 60029 230023 75299 230051
rect 75327 230023 75361 230051
rect 75389 230023 90659 230051
rect 90687 230023 90721 230051
rect 90749 230023 106019 230051
rect 106047 230023 106081 230051
rect 106109 230023 121379 230051
rect 121407 230023 121441 230051
rect 121469 230023 136739 230051
rect 136767 230023 136801 230051
rect 136829 230023 156485 230051
rect 156513 230023 156547 230051
rect 156575 230023 156609 230051
rect 156637 230023 156671 230051
rect 156699 230023 165485 230051
rect 165513 230023 165547 230051
rect 165575 230023 165609 230051
rect 165637 230023 165671 230051
rect 165699 230023 174485 230051
rect 174513 230023 174547 230051
rect 174575 230023 174609 230051
rect 174637 230023 174671 230051
rect 174699 230023 183485 230051
rect 183513 230023 183547 230051
rect 183575 230023 183609 230051
rect 183637 230023 183671 230051
rect 183699 230023 192485 230051
rect 192513 230023 192547 230051
rect 192575 230023 192609 230051
rect 192637 230023 192671 230051
rect 192699 230023 201485 230051
rect 201513 230023 201547 230051
rect 201575 230023 201609 230051
rect 201637 230023 201671 230051
rect 201699 230023 210485 230051
rect 210513 230023 210547 230051
rect 210575 230023 210609 230051
rect 210637 230023 210671 230051
rect 210699 230023 219485 230051
rect 219513 230023 219547 230051
rect 219575 230023 219609 230051
rect 219637 230023 219671 230051
rect 219699 230023 228485 230051
rect 228513 230023 228547 230051
rect 228575 230023 228609 230051
rect 228637 230023 228671 230051
rect 228699 230023 237485 230051
rect 237513 230023 237547 230051
rect 237575 230023 237609 230051
rect 237637 230023 237671 230051
rect 237699 230023 246485 230051
rect 246513 230023 246547 230051
rect 246575 230023 246609 230051
rect 246637 230023 246671 230051
rect 246699 230023 255485 230051
rect 255513 230023 255547 230051
rect 255575 230023 255609 230051
rect 255637 230023 255671 230051
rect 255699 230023 264485 230051
rect 264513 230023 264547 230051
rect 264575 230023 264609 230051
rect 264637 230023 264671 230051
rect 264699 230023 273485 230051
rect 273513 230023 273547 230051
rect 273575 230023 273609 230051
rect 273637 230023 273671 230051
rect 273699 230023 282485 230051
rect 282513 230023 282547 230051
rect 282575 230023 282609 230051
rect 282637 230023 282671 230051
rect 282699 230023 291485 230051
rect 291513 230023 291547 230051
rect 291575 230023 291609 230051
rect 291637 230023 291671 230051
rect 291699 230023 298728 230051
rect 298756 230023 298790 230051
rect 298818 230023 298852 230051
rect 298880 230023 298914 230051
rect 298942 230023 298990 230051
rect -958 229989 298990 230023
rect -958 229961 -910 229989
rect -882 229961 -848 229989
rect -820 229961 -786 229989
rect -758 229961 -724 229989
rect -696 229961 3485 229989
rect 3513 229961 3547 229989
rect 3575 229961 3609 229989
rect 3637 229961 3671 229989
rect 3699 229961 12485 229989
rect 12513 229961 12547 229989
rect 12575 229961 12609 229989
rect 12637 229961 12671 229989
rect 12699 229961 21485 229989
rect 21513 229961 21547 229989
rect 21575 229961 21609 229989
rect 21637 229961 21671 229989
rect 21699 229961 30485 229989
rect 30513 229961 30547 229989
rect 30575 229961 30609 229989
rect 30637 229961 30671 229989
rect 30699 229961 39485 229989
rect 39513 229961 39547 229989
rect 39575 229961 39609 229989
rect 39637 229961 39671 229989
rect 39699 229961 48485 229989
rect 48513 229961 48547 229989
rect 48575 229961 48609 229989
rect 48637 229961 48671 229989
rect 48699 229961 59939 229989
rect 59967 229961 60001 229989
rect 60029 229961 75299 229989
rect 75327 229961 75361 229989
rect 75389 229961 90659 229989
rect 90687 229961 90721 229989
rect 90749 229961 106019 229989
rect 106047 229961 106081 229989
rect 106109 229961 121379 229989
rect 121407 229961 121441 229989
rect 121469 229961 136739 229989
rect 136767 229961 136801 229989
rect 136829 229961 156485 229989
rect 156513 229961 156547 229989
rect 156575 229961 156609 229989
rect 156637 229961 156671 229989
rect 156699 229961 165485 229989
rect 165513 229961 165547 229989
rect 165575 229961 165609 229989
rect 165637 229961 165671 229989
rect 165699 229961 174485 229989
rect 174513 229961 174547 229989
rect 174575 229961 174609 229989
rect 174637 229961 174671 229989
rect 174699 229961 183485 229989
rect 183513 229961 183547 229989
rect 183575 229961 183609 229989
rect 183637 229961 183671 229989
rect 183699 229961 192485 229989
rect 192513 229961 192547 229989
rect 192575 229961 192609 229989
rect 192637 229961 192671 229989
rect 192699 229961 201485 229989
rect 201513 229961 201547 229989
rect 201575 229961 201609 229989
rect 201637 229961 201671 229989
rect 201699 229961 210485 229989
rect 210513 229961 210547 229989
rect 210575 229961 210609 229989
rect 210637 229961 210671 229989
rect 210699 229961 219485 229989
rect 219513 229961 219547 229989
rect 219575 229961 219609 229989
rect 219637 229961 219671 229989
rect 219699 229961 228485 229989
rect 228513 229961 228547 229989
rect 228575 229961 228609 229989
rect 228637 229961 228671 229989
rect 228699 229961 237485 229989
rect 237513 229961 237547 229989
rect 237575 229961 237609 229989
rect 237637 229961 237671 229989
rect 237699 229961 246485 229989
rect 246513 229961 246547 229989
rect 246575 229961 246609 229989
rect 246637 229961 246671 229989
rect 246699 229961 255485 229989
rect 255513 229961 255547 229989
rect 255575 229961 255609 229989
rect 255637 229961 255671 229989
rect 255699 229961 264485 229989
rect 264513 229961 264547 229989
rect 264575 229961 264609 229989
rect 264637 229961 264671 229989
rect 264699 229961 273485 229989
rect 273513 229961 273547 229989
rect 273575 229961 273609 229989
rect 273637 229961 273671 229989
rect 273699 229961 282485 229989
rect 282513 229961 282547 229989
rect 282575 229961 282609 229989
rect 282637 229961 282671 229989
rect 282699 229961 291485 229989
rect 291513 229961 291547 229989
rect 291575 229961 291609 229989
rect 291637 229961 291671 229989
rect 291699 229961 298728 229989
rect 298756 229961 298790 229989
rect 298818 229961 298852 229989
rect 298880 229961 298914 229989
rect 298942 229961 298990 229989
rect -958 229913 298990 229961
rect -958 227175 298990 227223
rect -958 227147 -430 227175
rect -402 227147 -368 227175
rect -340 227147 -306 227175
rect -278 227147 -244 227175
rect -216 227147 1625 227175
rect 1653 227147 1687 227175
rect 1715 227147 1749 227175
rect 1777 227147 1811 227175
rect 1839 227147 10625 227175
rect 10653 227147 10687 227175
rect 10715 227147 10749 227175
rect 10777 227147 10811 227175
rect 10839 227147 19625 227175
rect 19653 227147 19687 227175
rect 19715 227147 19749 227175
rect 19777 227147 19811 227175
rect 19839 227147 28625 227175
rect 28653 227147 28687 227175
rect 28715 227147 28749 227175
rect 28777 227147 28811 227175
rect 28839 227147 37625 227175
rect 37653 227147 37687 227175
rect 37715 227147 37749 227175
rect 37777 227147 37811 227175
rect 37839 227147 46625 227175
rect 46653 227147 46687 227175
rect 46715 227147 46749 227175
rect 46777 227147 46811 227175
rect 46839 227147 52259 227175
rect 52287 227147 52321 227175
rect 52349 227147 67619 227175
rect 67647 227147 67681 227175
rect 67709 227147 82979 227175
rect 83007 227147 83041 227175
rect 83069 227147 98339 227175
rect 98367 227147 98401 227175
rect 98429 227147 113699 227175
rect 113727 227147 113761 227175
rect 113789 227147 129059 227175
rect 129087 227147 129121 227175
rect 129149 227147 144419 227175
rect 144447 227147 144481 227175
rect 144509 227147 154625 227175
rect 154653 227147 154687 227175
rect 154715 227147 154749 227175
rect 154777 227147 154811 227175
rect 154839 227147 163625 227175
rect 163653 227147 163687 227175
rect 163715 227147 163749 227175
rect 163777 227147 163811 227175
rect 163839 227147 172625 227175
rect 172653 227147 172687 227175
rect 172715 227147 172749 227175
rect 172777 227147 172811 227175
rect 172839 227147 181625 227175
rect 181653 227147 181687 227175
rect 181715 227147 181749 227175
rect 181777 227147 181811 227175
rect 181839 227147 190625 227175
rect 190653 227147 190687 227175
rect 190715 227147 190749 227175
rect 190777 227147 190811 227175
rect 190839 227147 199625 227175
rect 199653 227147 199687 227175
rect 199715 227147 199749 227175
rect 199777 227147 199811 227175
rect 199839 227147 208625 227175
rect 208653 227147 208687 227175
rect 208715 227147 208749 227175
rect 208777 227147 208811 227175
rect 208839 227147 217625 227175
rect 217653 227147 217687 227175
rect 217715 227147 217749 227175
rect 217777 227147 217811 227175
rect 217839 227147 226625 227175
rect 226653 227147 226687 227175
rect 226715 227147 226749 227175
rect 226777 227147 226811 227175
rect 226839 227147 235625 227175
rect 235653 227147 235687 227175
rect 235715 227147 235749 227175
rect 235777 227147 235811 227175
rect 235839 227147 244625 227175
rect 244653 227147 244687 227175
rect 244715 227147 244749 227175
rect 244777 227147 244811 227175
rect 244839 227147 253625 227175
rect 253653 227147 253687 227175
rect 253715 227147 253749 227175
rect 253777 227147 253811 227175
rect 253839 227147 262625 227175
rect 262653 227147 262687 227175
rect 262715 227147 262749 227175
rect 262777 227147 262811 227175
rect 262839 227147 271625 227175
rect 271653 227147 271687 227175
rect 271715 227147 271749 227175
rect 271777 227147 271811 227175
rect 271839 227147 280625 227175
rect 280653 227147 280687 227175
rect 280715 227147 280749 227175
rect 280777 227147 280811 227175
rect 280839 227147 289625 227175
rect 289653 227147 289687 227175
rect 289715 227147 289749 227175
rect 289777 227147 289811 227175
rect 289839 227147 298248 227175
rect 298276 227147 298310 227175
rect 298338 227147 298372 227175
rect 298400 227147 298434 227175
rect 298462 227147 298990 227175
rect -958 227113 298990 227147
rect -958 227085 -430 227113
rect -402 227085 -368 227113
rect -340 227085 -306 227113
rect -278 227085 -244 227113
rect -216 227085 1625 227113
rect 1653 227085 1687 227113
rect 1715 227085 1749 227113
rect 1777 227085 1811 227113
rect 1839 227085 10625 227113
rect 10653 227085 10687 227113
rect 10715 227085 10749 227113
rect 10777 227085 10811 227113
rect 10839 227085 19625 227113
rect 19653 227085 19687 227113
rect 19715 227085 19749 227113
rect 19777 227085 19811 227113
rect 19839 227085 28625 227113
rect 28653 227085 28687 227113
rect 28715 227085 28749 227113
rect 28777 227085 28811 227113
rect 28839 227085 37625 227113
rect 37653 227085 37687 227113
rect 37715 227085 37749 227113
rect 37777 227085 37811 227113
rect 37839 227085 46625 227113
rect 46653 227085 46687 227113
rect 46715 227085 46749 227113
rect 46777 227085 46811 227113
rect 46839 227085 52259 227113
rect 52287 227085 52321 227113
rect 52349 227085 67619 227113
rect 67647 227085 67681 227113
rect 67709 227085 82979 227113
rect 83007 227085 83041 227113
rect 83069 227085 98339 227113
rect 98367 227085 98401 227113
rect 98429 227085 113699 227113
rect 113727 227085 113761 227113
rect 113789 227085 129059 227113
rect 129087 227085 129121 227113
rect 129149 227085 144419 227113
rect 144447 227085 144481 227113
rect 144509 227085 154625 227113
rect 154653 227085 154687 227113
rect 154715 227085 154749 227113
rect 154777 227085 154811 227113
rect 154839 227085 163625 227113
rect 163653 227085 163687 227113
rect 163715 227085 163749 227113
rect 163777 227085 163811 227113
rect 163839 227085 172625 227113
rect 172653 227085 172687 227113
rect 172715 227085 172749 227113
rect 172777 227085 172811 227113
rect 172839 227085 181625 227113
rect 181653 227085 181687 227113
rect 181715 227085 181749 227113
rect 181777 227085 181811 227113
rect 181839 227085 190625 227113
rect 190653 227085 190687 227113
rect 190715 227085 190749 227113
rect 190777 227085 190811 227113
rect 190839 227085 199625 227113
rect 199653 227085 199687 227113
rect 199715 227085 199749 227113
rect 199777 227085 199811 227113
rect 199839 227085 208625 227113
rect 208653 227085 208687 227113
rect 208715 227085 208749 227113
rect 208777 227085 208811 227113
rect 208839 227085 217625 227113
rect 217653 227085 217687 227113
rect 217715 227085 217749 227113
rect 217777 227085 217811 227113
rect 217839 227085 226625 227113
rect 226653 227085 226687 227113
rect 226715 227085 226749 227113
rect 226777 227085 226811 227113
rect 226839 227085 235625 227113
rect 235653 227085 235687 227113
rect 235715 227085 235749 227113
rect 235777 227085 235811 227113
rect 235839 227085 244625 227113
rect 244653 227085 244687 227113
rect 244715 227085 244749 227113
rect 244777 227085 244811 227113
rect 244839 227085 253625 227113
rect 253653 227085 253687 227113
rect 253715 227085 253749 227113
rect 253777 227085 253811 227113
rect 253839 227085 262625 227113
rect 262653 227085 262687 227113
rect 262715 227085 262749 227113
rect 262777 227085 262811 227113
rect 262839 227085 271625 227113
rect 271653 227085 271687 227113
rect 271715 227085 271749 227113
rect 271777 227085 271811 227113
rect 271839 227085 280625 227113
rect 280653 227085 280687 227113
rect 280715 227085 280749 227113
rect 280777 227085 280811 227113
rect 280839 227085 289625 227113
rect 289653 227085 289687 227113
rect 289715 227085 289749 227113
rect 289777 227085 289811 227113
rect 289839 227085 298248 227113
rect 298276 227085 298310 227113
rect 298338 227085 298372 227113
rect 298400 227085 298434 227113
rect 298462 227085 298990 227113
rect -958 227051 298990 227085
rect -958 227023 -430 227051
rect -402 227023 -368 227051
rect -340 227023 -306 227051
rect -278 227023 -244 227051
rect -216 227023 1625 227051
rect 1653 227023 1687 227051
rect 1715 227023 1749 227051
rect 1777 227023 1811 227051
rect 1839 227023 10625 227051
rect 10653 227023 10687 227051
rect 10715 227023 10749 227051
rect 10777 227023 10811 227051
rect 10839 227023 19625 227051
rect 19653 227023 19687 227051
rect 19715 227023 19749 227051
rect 19777 227023 19811 227051
rect 19839 227023 28625 227051
rect 28653 227023 28687 227051
rect 28715 227023 28749 227051
rect 28777 227023 28811 227051
rect 28839 227023 37625 227051
rect 37653 227023 37687 227051
rect 37715 227023 37749 227051
rect 37777 227023 37811 227051
rect 37839 227023 46625 227051
rect 46653 227023 46687 227051
rect 46715 227023 46749 227051
rect 46777 227023 46811 227051
rect 46839 227023 52259 227051
rect 52287 227023 52321 227051
rect 52349 227023 67619 227051
rect 67647 227023 67681 227051
rect 67709 227023 82979 227051
rect 83007 227023 83041 227051
rect 83069 227023 98339 227051
rect 98367 227023 98401 227051
rect 98429 227023 113699 227051
rect 113727 227023 113761 227051
rect 113789 227023 129059 227051
rect 129087 227023 129121 227051
rect 129149 227023 144419 227051
rect 144447 227023 144481 227051
rect 144509 227023 154625 227051
rect 154653 227023 154687 227051
rect 154715 227023 154749 227051
rect 154777 227023 154811 227051
rect 154839 227023 163625 227051
rect 163653 227023 163687 227051
rect 163715 227023 163749 227051
rect 163777 227023 163811 227051
rect 163839 227023 172625 227051
rect 172653 227023 172687 227051
rect 172715 227023 172749 227051
rect 172777 227023 172811 227051
rect 172839 227023 181625 227051
rect 181653 227023 181687 227051
rect 181715 227023 181749 227051
rect 181777 227023 181811 227051
rect 181839 227023 190625 227051
rect 190653 227023 190687 227051
rect 190715 227023 190749 227051
rect 190777 227023 190811 227051
rect 190839 227023 199625 227051
rect 199653 227023 199687 227051
rect 199715 227023 199749 227051
rect 199777 227023 199811 227051
rect 199839 227023 208625 227051
rect 208653 227023 208687 227051
rect 208715 227023 208749 227051
rect 208777 227023 208811 227051
rect 208839 227023 217625 227051
rect 217653 227023 217687 227051
rect 217715 227023 217749 227051
rect 217777 227023 217811 227051
rect 217839 227023 226625 227051
rect 226653 227023 226687 227051
rect 226715 227023 226749 227051
rect 226777 227023 226811 227051
rect 226839 227023 235625 227051
rect 235653 227023 235687 227051
rect 235715 227023 235749 227051
rect 235777 227023 235811 227051
rect 235839 227023 244625 227051
rect 244653 227023 244687 227051
rect 244715 227023 244749 227051
rect 244777 227023 244811 227051
rect 244839 227023 253625 227051
rect 253653 227023 253687 227051
rect 253715 227023 253749 227051
rect 253777 227023 253811 227051
rect 253839 227023 262625 227051
rect 262653 227023 262687 227051
rect 262715 227023 262749 227051
rect 262777 227023 262811 227051
rect 262839 227023 271625 227051
rect 271653 227023 271687 227051
rect 271715 227023 271749 227051
rect 271777 227023 271811 227051
rect 271839 227023 280625 227051
rect 280653 227023 280687 227051
rect 280715 227023 280749 227051
rect 280777 227023 280811 227051
rect 280839 227023 289625 227051
rect 289653 227023 289687 227051
rect 289715 227023 289749 227051
rect 289777 227023 289811 227051
rect 289839 227023 298248 227051
rect 298276 227023 298310 227051
rect 298338 227023 298372 227051
rect 298400 227023 298434 227051
rect 298462 227023 298990 227051
rect -958 226989 298990 227023
rect -958 226961 -430 226989
rect -402 226961 -368 226989
rect -340 226961 -306 226989
rect -278 226961 -244 226989
rect -216 226961 1625 226989
rect 1653 226961 1687 226989
rect 1715 226961 1749 226989
rect 1777 226961 1811 226989
rect 1839 226961 10625 226989
rect 10653 226961 10687 226989
rect 10715 226961 10749 226989
rect 10777 226961 10811 226989
rect 10839 226961 19625 226989
rect 19653 226961 19687 226989
rect 19715 226961 19749 226989
rect 19777 226961 19811 226989
rect 19839 226961 28625 226989
rect 28653 226961 28687 226989
rect 28715 226961 28749 226989
rect 28777 226961 28811 226989
rect 28839 226961 37625 226989
rect 37653 226961 37687 226989
rect 37715 226961 37749 226989
rect 37777 226961 37811 226989
rect 37839 226961 46625 226989
rect 46653 226961 46687 226989
rect 46715 226961 46749 226989
rect 46777 226961 46811 226989
rect 46839 226961 52259 226989
rect 52287 226961 52321 226989
rect 52349 226961 67619 226989
rect 67647 226961 67681 226989
rect 67709 226961 82979 226989
rect 83007 226961 83041 226989
rect 83069 226961 98339 226989
rect 98367 226961 98401 226989
rect 98429 226961 113699 226989
rect 113727 226961 113761 226989
rect 113789 226961 129059 226989
rect 129087 226961 129121 226989
rect 129149 226961 144419 226989
rect 144447 226961 144481 226989
rect 144509 226961 154625 226989
rect 154653 226961 154687 226989
rect 154715 226961 154749 226989
rect 154777 226961 154811 226989
rect 154839 226961 163625 226989
rect 163653 226961 163687 226989
rect 163715 226961 163749 226989
rect 163777 226961 163811 226989
rect 163839 226961 172625 226989
rect 172653 226961 172687 226989
rect 172715 226961 172749 226989
rect 172777 226961 172811 226989
rect 172839 226961 181625 226989
rect 181653 226961 181687 226989
rect 181715 226961 181749 226989
rect 181777 226961 181811 226989
rect 181839 226961 190625 226989
rect 190653 226961 190687 226989
rect 190715 226961 190749 226989
rect 190777 226961 190811 226989
rect 190839 226961 199625 226989
rect 199653 226961 199687 226989
rect 199715 226961 199749 226989
rect 199777 226961 199811 226989
rect 199839 226961 208625 226989
rect 208653 226961 208687 226989
rect 208715 226961 208749 226989
rect 208777 226961 208811 226989
rect 208839 226961 217625 226989
rect 217653 226961 217687 226989
rect 217715 226961 217749 226989
rect 217777 226961 217811 226989
rect 217839 226961 226625 226989
rect 226653 226961 226687 226989
rect 226715 226961 226749 226989
rect 226777 226961 226811 226989
rect 226839 226961 235625 226989
rect 235653 226961 235687 226989
rect 235715 226961 235749 226989
rect 235777 226961 235811 226989
rect 235839 226961 244625 226989
rect 244653 226961 244687 226989
rect 244715 226961 244749 226989
rect 244777 226961 244811 226989
rect 244839 226961 253625 226989
rect 253653 226961 253687 226989
rect 253715 226961 253749 226989
rect 253777 226961 253811 226989
rect 253839 226961 262625 226989
rect 262653 226961 262687 226989
rect 262715 226961 262749 226989
rect 262777 226961 262811 226989
rect 262839 226961 271625 226989
rect 271653 226961 271687 226989
rect 271715 226961 271749 226989
rect 271777 226961 271811 226989
rect 271839 226961 280625 226989
rect 280653 226961 280687 226989
rect 280715 226961 280749 226989
rect 280777 226961 280811 226989
rect 280839 226961 289625 226989
rect 289653 226961 289687 226989
rect 289715 226961 289749 226989
rect 289777 226961 289811 226989
rect 289839 226961 298248 226989
rect 298276 226961 298310 226989
rect 298338 226961 298372 226989
rect 298400 226961 298434 226989
rect 298462 226961 298990 226989
rect -958 226913 298990 226961
rect -958 221175 298990 221223
rect -958 221147 -910 221175
rect -882 221147 -848 221175
rect -820 221147 -786 221175
rect -758 221147 -724 221175
rect -696 221147 3485 221175
rect 3513 221147 3547 221175
rect 3575 221147 3609 221175
rect 3637 221147 3671 221175
rect 3699 221147 12485 221175
rect 12513 221147 12547 221175
rect 12575 221147 12609 221175
rect 12637 221147 12671 221175
rect 12699 221147 21485 221175
rect 21513 221147 21547 221175
rect 21575 221147 21609 221175
rect 21637 221147 21671 221175
rect 21699 221147 30485 221175
rect 30513 221147 30547 221175
rect 30575 221147 30609 221175
rect 30637 221147 30671 221175
rect 30699 221147 39485 221175
rect 39513 221147 39547 221175
rect 39575 221147 39609 221175
rect 39637 221147 39671 221175
rect 39699 221147 48485 221175
rect 48513 221147 48547 221175
rect 48575 221147 48609 221175
rect 48637 221147 48671 221175
rect 48699 221147 59939 221175
rect 59967 221147 60001 221175
rect 60029 221147 75299 221175
rect 75327 221147 75361 221175
rect 75389 221147 90659 221175
rect 90687 221147 90721 221175
rect 90749 221147 106019 221175
rect 106047 221147 106081 221175
rect 106109 221147 121379 221175
rect 121407 221147 121441 221175
rect 121469 221147 136739 221175
rect 136767 221147 136801 221175
rect 136829 221147 156485 221175
rect 156513 221147 156547 221175
rect 156575 221147 156609 221175
rect 156637 221147 156671 221175
rect 156699 221147 165485 221175
rect 165513 221147 165547 221175
rect 165575 221147 165609 221175
rect 165637 221147 165671 221175
rect 165699 221147 174485 221175
rect 174513 221147 174547 221175
rect 174575 221147 174609 221175
rect 174637 221147 174671 221175
rect 174699 221147 183485 221175
rect 183513 221147 183547 221175
rect 183575 221147 183609 221175
rect 183637 221147 183671 221175
rect 183699 221147 192485 221175
rect 192513 221147 192547 221175
rect 192575 221147 192609 221175
rect 192637 221147 192671 221175
rect 192699 221147 201485 221175
rect 201513 221147 201547 221175
rect 201575 221147 201609 221175
rect 201637 221147 201671 221175
rect 201699 221147 210485 221175
rect 210513 221147 210547 221175
rect 210575 221147 210609 221175
rect 210637 221147 210671 221175
rect 210699 221147 219485 221175
rect 219513 221147 219547 221175
rect 219575 221147 219609 221175
rect 219637 221147 219671 221175
rect 219699 221147 228485 221175
rect 228513 221147 228547 221175
rect 228575 221147 228609 221175
rect 228637 221147 228671 221175
rect 228699 221147 237485 221175
rect 237513 221147 237547 221175
rect 237575 221147 237609 221175
rect 237637 221147 237671 221175
rect 237699 221147 246485 221175
rect 246513 221147 246547 221175
rect 246575 221147 246609 221175
rect 246637 221147 246671 221175
rect 246699 221147 255485 221175
rect 255513 221147 255547 221175
rect 255575 221147 255609 221175
rect 255637 221147 255671 221175
rect 255699 221147 264485 221175
rect 264513 221147 264547 221175
rect 264575 221147 264609 221175
rect 264637 221147 264671 221175
rect 264699 221147 273485 221175
rect 273513 221147 273547 221175
rect 273575 221147 273609 221175
rect 273637 221147 273671 221175
rect 273699 221147 282485 221175
rect 282513 221147 282547 221175
rect 282575 221147 282609 221175
rect 282637 221147 282671 221175
rect 282699 221147 291485 221175
rect 291513 221147 291547 221175
rect 291575 221147 291609 221175
rect 291637 221147 291671 221175
rect 291699 221147 298728 221175
rect 298756 221147 298790 221175
rect 298818 221147 298852 221175
rect 298880 221147 298914 221175
rect 298942 221147 298990 221175
rect -958 221113 298990 221147
rect -958 221085 -910 221113
rect -882 221085 -848 221113
rect -820 221085 -786 221113
rect -758 221085 -724 221113
rect -696 221085 3485 221113
rect 3513 221085 3547 221113
rect 3575 221085 3609 221113
rect 3637 221085 3671 221113
rect 3699 221085 12485 221113
rect 12513 221085 12547 221113
rect 12575 221085 12609 221113
rect 12637 221085 12671 221113
rect 12699 221085 21485 221113
rect 21513 221085 21547 221113
rect 21575 221085 21609 221113
rect 21637 221085 21671 221113
rect 21699 221085 30485 221113
rect 30513 221085 30547 221113
rect 30575 221085 30609 221113
rect 30637 221085 30671 221113
rect 30699 221085 39485 221113
rect 39513 221085 39547 221113
rect 39575 221085 39609 221113
rect 39637 221085 39671 221113
rect 39699 221085 48485 221113
rect 48513 221085 48547 221113
rect 48575 221085 48609 221113
rect 48637 221085 48671 221113
rect 48699 221085 59939 221113
rect 59967 221085 60001 221113
rect 60029 221085 75299 221113
rect 75327 221085 75361 221113
rect 75389 221085 90659 221113
rect 90687 221085 90721 221113
rect 90749 221085 106019 221113
rect 106047 221085 106081 221113
rect 106109 221085 121379 221113
rect 121407 221085 121441 221113
rect 121469 221085 136739 221113
rect 136767 221085 136801 221113
rect 136829 221085 156485 221113
rect 156513 221085 156547 221113
rect 156575 221085 156609 221113
rect 156637 221085 156671 221113
rect 156699 221085 165485 221113
rect 165513 221085 165547 221113
rect 165575 221085 165609 221113
rect 165637 221085 165671 221113
rect 165699 221085 174485 221113
rect 174513 221085 174547 221113
rect 174575 221085 174609 221113
rect 174637 221085 174671 221113
rect 174699 221085 183485 221113
rect 183513 221085 183547 221113
rect 183575 221085 183609 221113
rect 183637 221085 183671 221113
rect 183699 221085 192485 221113
rect 192513 221085 192547 221113
rect 192575 221085 192609 221113
rect 192637 221085 192671 221113
rect 192699 221085 201485 221113
rect 201513 221085 201547 221113
rect 201575 221085 201609 221113
rect 201637 221085 201671 221113
rect 201699 221085 210485 221113
rect 210513 221085 210547 221113
rect 210575 221085 210609 221113
rect 210637 221085 210671 221113
rect 210699 221085 219485 221113
rect 219513 221085 219547 221113
rect 219575 221085 219609 221113
rect 219637 221085 219671 221113
rect 219699 221085 228485 221113
rect 228513 221085 228547 221113
rect 228575 221085 228609 221113
rect 228637 221085 228671 221113
rect 228699 221085 237485 221113
rect 237513 221085 237547 221113
rect 237575 221085 237609 221113
rect 237637 221085 237671 221113
rect 237699 221085 246485 221113
rect 246513 221085 246547 221113
rect 246575 221085 246609 221113
rect 246637 221085 246671 221113
rect 246699 221085 255485 221113
rect 255513 221085 255547 221113
rect 255575 221085 255609 221113
rect 255637 221085 255671 221113
rect 255699 221085 264485 221113
rect 264513 221085 264547 221113
rect 264575 221085 264609 221113
rect 264637 221085 264671 221113
rect 264699 221085 273485 221113
rect 273513 221085 273547 221113
rect 273575 221085 273609 221113
rect 273637 221085 273671 221113
rect 273699 221085 282485 221113
rect 282513 221085 282547 221113
rect 282575 221085 282609 221113
rect 282637 221085 282671 221113
rect 282699 221085 291485 221113
rect 291513 221085 291547 221113
rect 291575 221085 291609 221113
rect 291637 221085 291671 221113
rect 291699 221085 298728 221113
rect 298756 221085 298790 221113
rect 298818 221085 298852 221113
rect 298880 221085 298914 221113
rect 298942 221085 298990 221113
rect -958 221051 298990 221085
rect -958 221023 -910 221051
rect -882 221023 -848 221051
rect -820 221023 -786 221051
rect -758 221023 -724 221051
rect -696 221023 3485 221051
rect 3513 221023 3547 221051
rect 3575 221023 3609 221051
rect 3637 221023 3671 221051
rect 3699 221023 12485 221051
rect 12513 221023 12547 221051
rect 12575 221023 12609 221051
rect 12637 221023 12671 221051
rect 12699 221023 21485 221051
rect 21513 221023 21547 221051
rect 21575 221023 21609 221051
rect 21637 221023 21671 221051
rect 21699 221023 30485 221051
rect 30513 221023 30547 221051
rect 30575 221023 30609 221051
rect 30637 221023 30671 221051
rect 30699 221023 39485 221051
rect 39513 221023 39547 221051
rect 39575 221023 39609 221051
rect 39637 221023 39671 221051
rect 39699 221023 48485 221051
rect 48513 221023 48547 221051
rect 48575 221023 48609 221051
rect 48637 221023 48671 221051
rect 48699 221023 59939 221051
rect 59967 221023 60001 221051
rect 60029 221023 75299 221051
rect 75327 221023 75361 221051
rect 75389 221023 90659 221051
rect 90687 221023 90721 221051
rect 90749 221023 106019 221051
rect 106047 221023 106081 221051
rect 106109 221023 121379 221051
rect 121407 221023 121441 221051
rect 121469 221023 136739 221051
rect 136767 221023 136801 221051
rect 136829 221023 156485 221051
rect 156513 221023 156547 221051
rect 156575 221023 156609 221051
rect 156637 221023 156671 221051
rect 156699 221023 165485 221051
rect 165513 221023 165547 221051
rect 165575 221023 165609 221051
rect 165637 221023 165671 221051
rect 165699 221023 174485 221051
rect 174513 221023 174547 221051
rect 174575 221023 174609 221051
rect 174637 221023 174671 221051
rect 174699 221023 183485 221051
rect 183513 221023 183547 221051
rect 183575 221023 183609 221051
rect 183637 221023 183671 221051
rect 183699 221023 192485 221051
rect 192513 221023 192547 221051
rect 192575 221023 192609 221051
rect 192637 221023 192671 221051
rect 192699 221023 201485 221051
rect 201513 221023 201547 221051
rect 201575 221023 201609 221051
rect 201637 221023 201671 221051
rect 201699 221023 210485 221051
rect 210513 221023 210547 221051
rect 210575 221023 210609 221051
rect 210637 221023 210671 221051
rect 210699 221023 219485 221051
rect 219513 221023 219547 221051
rect 219575 221023 219609 221051
rect 219637 221023 219671 221051
rect 219699 221023 228485 221051
rect 228513 221023 228547 221051
rect 228575 221023 228609 221051
rect 228637 221023 228671 221051
rect 228699 221023 237485 221051
rect 237513 221023 237547 221051
rect 237575 221023 237609 221051
rect 237637 221023 237671 221051
rect 237699 221023 246485 221051
rect 246513 221023 246547 221051
rect 246575 221023 246609 221051
rect 246637 221023 246671 221051
rect 246699 221023 255485 221051
rect 255513 221023 255547 221051
rect 255575 221023 255609 221051
rect 255637 221023 255671 221051
rect 255699 221023 264485 221051
rect 264513 221023 264547 221051
rect 264575 221023 264609 221051
rect 264637 221023 264671 221051
rect 264699 221023 273485 221051
rect 273513 221023 273547 221051
rect 273575 221023 273609 221051
rect 273637 221023 273671 221051
rect 273699 221023 282485 221051
rect 282513 221023 282547 221051
rect 282575 221023 282609 221051
rect 282637 221023 282671 221051
rect 282699 221023 291485 221051
rect 291513 221023 291547 221051
rect 291575 221023 291609 221051
rect 291637 221023 291671 221051
rect 291699 221023 298728 221051
rect 298756 221023 298790 221051
rect 298818 221023 298852 221051
rect 298880 221023 298914 221051
rect 298942 221023 298990 221051
rect -958 220989 298990 221023
rect -958 220961 -910 220989
rect -882 220961 -848 220989
rect -820 220961 -786 220989
rect -758 220961 -724 220989
rect -696 220961 3485 220989
rect 3513 220961 3547 220989
rect 3575 220961 3609 220989
rect 3637 220961 3671 220989
rect 3699 220961 12485 220989
rect 12513 220961 12547 220989
rect 12575 220961 12609 220989
rect 12637 220961 12671 220989
rect 12699 220961 21485 220989
rect 21513 220961 21547 220989
rect 21575 220961 21609 220989
rect 21637 220961 21671 220989
rect 21699 220961 30485 220989
rect 30513 220961 30547 220989
rect 30575 220961 30609 220989
rect 30637 220961 30671 220989
rect 30699 220961 39485 220989
rect 39513 220961 39547 220989
rect 39575 220961 39609 220989
rect 39637 220961 39671 220989
rect 39699 220961 48485 220989
rect 48513 220961 48547 220989
rect 48575 220961 48609 220989
rect 48637 220961 48671 220989
rect 48699 220961 59939 220989
rect 59967 220961 60001 220989
rect 60029 220961 75299 220989
rect 75327 220961 75361 220989
rect 75389 220961 90659 220989
rect 90687 220961 90721 220989
rect 90749 220961 106019 220989
rect 106047 220961 106081 220989
rect 106109 220961 121379 220989
rect 121407 220961 121441 220989
rect 121469 220961 136739 220989
rect 136767 220961 136801 220989
rect 136829 220961 156485 220989
rect 156513 220961 156547 220989
rect 156575 220961 156609 220989
rect 156637 220961 156671 220989
rect 156699 220961 165485 220989
rect 165513 220961 165547 220989
rect 165575 220961 165609 220989
rect 165637 220961 165671 220989
rect 165699 220961 174485 220989
rect 174513 220961 174547 220989
rect 174575 220961 174609 220989
rect 174637 220961 174671 220989
rect 174699 220961 183485 220989
rect 183513 220961 183547 220989
rect 183575 220961 183609 220989
rect 183637 220961 183671 220989
rect 183699 220961 192485 220989
rect 192513 220961 192547 220989
rect 192575 220961 192609 220989
rect 192637 220961 192671 220989
rect 192699 220961 201485 220989
rect 201513 220961 201547 220989
rect 201575 220961 201609 220989
rect 201637 220961 201671 220989
rect 201699 220961 210485 220989
rect 210513 220961 210547 220989
rect 210575 220961 210609 220989
rect 210637 220961 210671 220989
rect 210699 220961 219485 220989
rect 219513 220961 219547 220989
rect 219575 220961 219609 220989
rect 219637 220961 219671 220989
rect 219699 220961 228485 220989
rect 228513 220961 228547 220989
rect 228575 220961 228609 220989
rect 228637 220961 228671 220989
rect 228699 220961 237485 220989
rect 237513 220961 237547 220989
rect 237575 220961 237609 220989
rect 237637 220961 237671 220989
rect 237699 220961 246485 220989
rect 246513 220961 246547 220989
rect 246575 220961 246609 220989
rect 246637 220961 246671 220989
rect 246699 220961 255485 220989
rect 255513 220961 255547 220989
rect 255575 220961 255609 220989
rect 255637 220961 255671 220989
rect 255699 220961 264485 220989
rect 264513 220961 264547 220989
rect 264575 220961 264609 220989
rect 264637 220961 264671 220989
rect 264699 220961 273485 220989
rect 273513 220961 273547 220989
rect 273575 220961 273609 220989
rect 273637 220961 273671 220989
rect 273699 220961 282485 220989
rect 282513 220961 282547 220989
rect 282575 220961 282609 220989
rect 282637 220961 282671 220989
rect 282699 220961 291485 220989
rect 291513 220961 291547 220989
rect 291575 220961 291609 220989
rect 291637 220961 291671 220989
rect 291699 220961 298728 220989
rect 298756 220961 298790 220989
rect 298818 220961 298852 220989
rect 298880 220961 298914 220989
rect 298942 220961 298990 220989
rect -958 220913 298990 220961
rect -958 218175 298990 218223
rect -958 218147 -430 218175
rect -402 218147 -368 218175
rect -340 218147 -306 218175
rect -278 218147 -244 218175
rect -216 218147 1625 218175
rect 1653 218147 1687 218175
rect 1715 218147 1749 218175
rect 1777 218147 1811 218175
rect 1839 218147 10625 218175
rect 10653 218147 10687 218175
rect 10715 218147 10749 218175
rect 10777 218147 10811 218175
rect 10839 218147 19625 218175
rect 19653 218147 19687 218175
rect 19715 218147 19749 218175
rect 19777 218147 19811 218175
rect 19839 218147 28625 218175
rect 28653 218147 28687 218175
rect 28715 218147 28749 218175
rect 28777 218147 28811 218175
rect 28839 218147 37625 218175
rect 37653 218147 37687 218175
rect 37715 218147 37749 218175
rect 37777 218147 37811 218175
rect 37839 218147 46625 218175
rect 46653 218147 46687 218175
rect 46715 218147 46749 218175
rect 46777 218147 46811 218175
rect 46839 218147 52259 218175
rect 52287 218147 52321 218175
rect 52349 218147 67619 218175
rect 67647 218147 67681 218175
rect 67709 218147 82979 218175
rect 83007 218147 83041 218175
rect 83069 218147 98339 218175
rect 98367 218147 98401 218175
rect 98429 218147 113699 218175
rect 113727 218147 113761 218175
rect 113789 218147 129059 218175
rect 129087 218147 129121 218175
rect 129149 218147 144419 218175
rect 144447 218147 144481 218175
rect 144509 218147 154625 218175
rect 154653 218147 154687 218175
rect 154715 218147 154749 218175
rect 154777 218147 154811 218175
rect 154839 218147 163625 218175
rect 163653 218147 163687 218175
rect 163715 218147 163749 218175
rect 163777 218147 163811 218175
rect 163839 218147 172625 218175
rect 172653 218147 172687 218175
rect 172715 218147 172749 218175
rect 172777 218147 172811 218175
rect 172839 218147 181625 218175
rect 181653 218147 181687 218175
rect 181715 218147 181749 218175
rect 181777 218147 181811 218175
rect 181839 218147 190625 218175
rect 190653 218147 190687 218175
rect 190715 218147 190749 218175
rect 190777 218147 190811 218175
rect 190839 218147 199625 218175
rect 199653 218147 199687 218175
rect 199715 218147 199749 218175
rect 199777 218147 199811 218175
rect 199839 218147 208625 218175
rect 208653 218147 208687 218175
rect 208715 218147 208749 218175
rect 208777 218147 208811 218175
rect 208839 218147 217625 218175
rect 217653 218147 217687 218175
rect 217715 218147 217749 218175
rect 217777 218147 217811 218175
rect 217839 218147 226625 218175
rect 226653 218147 226687 218175
rect 226715 218147 226749 218175
rect 226777 218147 226811 218175
rect 226839 218147 235625 218175
rect 235653 218147 235687 218175
rect 235715 218147 235749 218175
rect 235777 218147 235811 218175
rect 235839 218147 244625 218175
rect 244653 218147 244687 218175
rect 244715 218147 244749 218175
rect 244777 218147 244811 218175
rect 244839 218147 253625 218175
rect 253653 218147 253687 218175
rect 253715 218147 253749 218175
rect 253777 218147 253811 218175
rect 253839 218147 262625 218175
rect 262653 218147 262687 218175
rect 262715 218147 262749 218175
rect 262777 218147 262811 218175
rect 262839 218147 271625 218175
rect 271653 218147 271687 218175
rect 271715 218147 271749 218175
rect 271777 218147 271811 218175
rect 271839 218147 280625 218175
rect 280653 218147 280687 218175
rect 280715 218147 280749 218175
rect 280777 218147 280811 218175
rect 280839 218147 289625 218175
rect 289653 218147 289687 218175
rect 289715 218147 289749 218175
rect 289777 218147 289811 218175
rect 289839 218147 298248 218175
rect 298276 218147 298310 218175
rect 298338 218147 298372 218175
rect 298400 218147 298434 218175
rect 298462 218147 298990 218175
rect -958 218113 298990 218147
rect -958 218085 -430 218113
rect -402 218085 -368 218113
rect -340 218085 -306 218113
rect -278 218085 -244 218113
rect -216 218085 1625 218113
rect 1653 218085 1687 218113
rect 1715 218085 1749 218113
rect 1777 218085 1811 218113
rect 1839 218085 10625 218113
rect 10653 218085 10687 218113
rect 10715 218085 10749 218113
rect 10777 218085 10811 218113
rect 10839 218085 19625 218113
rect 19653 218085 19687 218113
rect 19715 218085 19749 218113
rect 19777 218085 19811 218113
rect 19839 218085 28625 218113
rect 28653 218085 28687 218113
rect 28715 218085 28749 218113
rect 28777 218085 28811 218113
rect 28839 218085 37625 218113
rect 37653 218085 37687 218113
rect 37715 218085 37749 218113
rect 37777 218085 37811 218113
rect 37839 218085 46625 218113
rect 46653 218085 46687 218113
rect 46715 218085 46749 218113
rect 46777 218085 46811 218113
rect 46839 218085 52259 218113
rect 52287 218085 52321 218113
rect 52349 218085 67619 218113
rect 67647 218085 67681 218113
rect 67709 218085 82979 218113
rect 83007 218085 83041 218113
rect 83069 218085 98339 218113
rect 98367 218085 98401 218113
rect 98429 218085 113699 218113
rect 113727 218085 113761 218113
rect 113789 218085 129059 218113
rect 129087 218085 129121 218113
rect 129149 218085 144419 218113
rect 144447 218085 144481 218113
rect 144509 218085 154625 218113
rect 154653 218085 154687 218113
rect 154715 218085 154749 218113
rect 154777 218085 154811 218113
rect 154839 218085 163625 218113
rect 163653 218085 163687 218113
rect 163715 218085 163749 218113
rect 163777 218085 163811 218113
rect 163839 218085 172625 218113
rect 172653 218085 172687 218113
rect 172715 218085 172749 218113
rect 172777 218085 172811 218113
rect 172839 218085 181625 218113
rect 181653 218085 181687 218113
rect 181715 218085 181749 218113
rect 181777 218085 181811 218113
rect 181839 218085 190625 218113
rect 190653 218085 190687 218113
rect 190715 218085 190749 218113
rect 190777 218085 190811 218113
rect 190839 218085 199625 218113
rect 199653 218085 199687 218113
rect 199715 218085 199749 218113
rect 199777 218085 199811 218113
rect 199839 218085 208625 218113
rect 208653 218085 208687 218113
rect 208715 218085 208749 218113
rect 208777 218085 208811 218113
rect 208839 218085 217625 218113
rect 217653 218085 217687 218113
rect 217715 218085 217749 218113
rect 217777 218085 217811 218113
rect 217839 218085 226625 218113
rect 226653 218085 226687 218113
rect 226715 218085 226749 218113
rect 226777 218085 226811 218113
rect 226839 218085 235625 218113
rect 235653 218085 235687 218113
rect 235715 218085 235749 218113
rect 235777 218085 235811 218113
rect 235839 218085 244625 218113
rect 244653 218085 244687 218113
rect 244715 218085 244749 218113
rect 244777 218085 244811 218113
rect 244839 218085 253625 218113
rect 253653 218085 253687 218113
rect 253715 218085 253749 218113
rect 253777 218085 253811 218113
rect 253839 218085 262625 218113
rect 262653 218085 262687 218113
rect 262715 218085 262749 218113
rect 262777 218085 262811 218113
rect 262839 218085 271625 218113
rect 271653 218085 271687 218113
rect 271715 218085 271749 218113
rect 271777 218085 271811 218113
rect 271839 218085 280625 218113
rect 280653 218085 280687 218113
rect 280715 218085 280749 218113
rect 280777 218085 280811 218113
rect 280839 218085 289625 218113
rect 289653 218085 289687 218113
rect 289715 218085 289749 218113
rect 289777 218085 289811 218113
rect 289839 218085 298248 218113
rect 298276 218085 298310 218113
rect 298338 218085 298372 218113
rect 298400 218085 298434 218113
rect 298462 218085 298990 218113
rect -958 218051 298990 218085
rect -958 218023 -430 218051
rect -402 218023 -368 218051
rect -340 218023 -306 218051
rect -278 218023 -244 218051
rect -216 218023 1625 218051
rect 1653 218023 1687 218051
rect 1715 218023 1749 218051
rect 1777 218023 1811 218051
rect 1839 218023 10625 218051
rect 10653 218023 10687 218051
rect 10715 218023 10749 218051
rect 10777 218023 10811 218051
rect 10839 218023 19625 218051
rect 19653 218023 19687 218051
rect 19715 218023 19749 218051
rect 19777 218023 19811 218051
rect 19839 218023 28625 218051
rect 28653 218023 28687 218051
rect 28715 218023 28749 218051
rect 28777 218023 28811 218051
rect 28839 218023 37625 218051
rect 37653 218023 37687 218051
rect 37715 218023 37749 218051
rect 37777 218023 37811 218051
rect 37839 218023 46625 218051
rect 46653 218023 46687 218051
rect 46715 218023 46749 218051
rect 46777 218023 46811 218051
rect 46839 218023 52259 218051
rect 52287 218023 52321 218051
rect 52349 218023 67619 218051
rect 67647 218023 67681 218051
rect 67709 218023 82979 218051
rect 83007 218023 83041 218051
rect 83069 218023 98339 218051
rect 98367 218023 98401 218051
rect 98429 218023 113699 218051
rect 113727 218023 113761 218051
rect 113789 218023 129059 218051
rect 129087 218023 129121 218051
rect 129149 218023 144419 218051
rect 144447 218023 144481 218051
rect 144509 218023 154625 218051
rect 154653 218023 154687 218051
rect 154715 218023 154749 218051
rect 154777 218023 154811 218051
rect 154839 218023 163625 218051
rect 163653 218023 163687 218051
rect 163715 218023 163749 218051
rect 163777 218023 163811 218051
rect 163839 218023 172625 218051
rect 172653 218023 172687 218051
rect 172715 218023 172749 218051
rect 172777 218023 172811 218051
rect 172839 218023 181625 218051
rect 181653 218023 181687 218051
rect 181715 218023 181749 218051
rect 181777 218023 181811 218051
rect 181839 218023 190625 218051
rect 190653 218023 190687 218051
rect 190715 218023 190749 218051
rect 190777 218023 190811 218051
rect 190839 218023 199625 218051
rect 199653 218023 199687 218051
rect 199715 218023 199749 218051
rect 199777 218023 199811 218051
rect 199839 218023 208625 218051
rect 208653 218023 208687 218051
rect 208715 218023 208749 218051
rect 208777 218023 208811 218051
rect 208839 218023 217625 218051
rect 217653 218023 217687 218051
rect 217715 218023 217749 218051
rect 217777 218023 217811 218051
rect 217839 218023 226625 218051
rect 226653 218023 226687 218051
rect 226715 218023 226749 218051
rect 226777 218023 226811 218051
rect 226839 218023 235625 218051
rect 235653 218023 235687 218051
rect 235715 218023 235749 218051
rect 235777 218023 235811 218051
rect 235839 218023 244625 218051
rect 244653 218023 244687 218051
rect 244715 218023 244749 218051
rect 244777 218023 244811 218051
rect 244839 218023 253625 218051
rect 253653 218023 253687 218051
rect 253715 218023 253749 218051
rect 253777 218023 253811 218051
rect 253839 218023 262625 218051
rect 262653 218023 262687 218051
rect 262715 218023 262749 218051
rect 262777 218023 262811 218051
rect 262839 218023 271625 218051
rect 271653 218023 271687 218051
rect 271715 218023 271749 218051
rect 271777 218023 271811 218051
rect 271839 218023 280625 218051
rect 280653 218023 280687 218051
rect 280715 218023 280749 218051
rect 280777 218023 280811 218051
rect 280839 218023 289625 218051
rect 289653 218023 289687 218051
rect 289715 218023 289749 218051
rect 289777 218023 289811 218051
rect 289839 218023 298248 218051
rect 298276 218023 298310 218051
rect 298338 218023 298372 218051
rect 298400 218023 298434 218051
rect 298462 218023 298990 218051
rect -958 217989 298990 218023
rect -958 217961 -430 217989
rect -402 217961 -368 217989
rect -340 217961 -306 217989
rect -278 217961 -244 217989
rect -216 217961 1625 217989
rect 1653 217961 1687 217989
rect 1715 217961 1749 217989
rect 1777 217961 1811 217989
rect 1839 217961 10625 217989
rect 10653 217961 10687 217989
rect 10715 217961 10749 217989
rect 10777 217961 10811 217989
rect 10839 217961 19625 217989
rect 19653 217961 19687 217989
rect 19715 217961 19749 217989
rect 19777 217961 19811 217989
rect 19839 217961 28625 217989
rect 28653 217961 28687 217989
rect 28715 217961 28749 217989
rect 28777 217961 28811 217989
rect 28839 217961 37625 217989
rect 37653 217961 37687 217989
rect 37715 217961 37749 217989
rect 37777 217961 37811 217989
rect 37839 217961 46625 217989
rect 46653 217961 46687 217989
rect 46715 217961 46749 217989
rect 46777 217961 46811 217989
rect 46839 217961 52259 217989
rect 52287 217961 52321 217989
rect 52349 217961 67619 217989
rect 67647 217961 67681 217989
rect 67709 217961 82979 217989
rect 83007 217961 83041 217989
rect 83069 217961 98339 217989
rect 98367 217961 98401 217989
rect 98429 217961 113699 217989
rect 113727 217961 113761 217989
rect 113789 217961 129059 217989
rect 129087 217961 129121 217989
rect 129149 217961 144419 217989
rect 144447 217961 144481 217989
rect 144509 217961 154625 217989
rect 154653 217961 154687 217989
rect 154715 217961 154749 217989
rect 154777 217961 154811 217989
rect 154839 217961 163625 217989
rect 163653 217961 163687 217989
rect 163715 217961 163749 217989
rect 163777 217961 163811 217989
rect 163839 217961 172625 217989
rect 172653 217961 172687 217989
rect 172715 217961 172749 217989
rect 172777 217961 172811 217989
rect 172839 217961 181625 217989
rect 181653 217961 181687 217989
rect 181715 217961 181749 217989
rect 181777 217961 181811 217989
rect 181839 217961 190625 217989
rect 190653 217961 190687 217989
rect 190715 217961 190749 217989
rect 190777 217961 190811 217989
rect 190839 217961 199625 217989
rect 199653 217961 199687 217989
rect 199715 217961 199749 217989
rect 199777 217961 199811 217989
rect 199839 217961 208625 217989
rect 208653 217961 208687 217989
rect 208715 217961 208749 217989
rect 208777 217961 208811 217989
rect 208839 217961 217625 217989
rect 217653 217961 217687 217989
rect 217715 217961 217749 217989
rect 217777 217961 217811 217989
rect 217839 217961 226625 217989
rect 226653 217961 226687 217989
rect 226715 217961 226749 217989
rect 226777 217961 226811 217989
rect 226839 217961 235625 217989
rect 235653 217961 235687 217989
rect 235715 217961 235749 217989
rect 235777 217961 235811 217989
rect 235839 217961 244625 217989
rect 244653 217961 244687 217989
rect 244715 217961 244749 217989
rect 244777 217961 244811 217989
rect 244839 217961 253625 217989
rect 253653 217961 253687 217989
rect 253715 217961 253749 217989
rect 253777 217961 253811 217989
rect 253839 217961 262625 217989
rect 262653 217961 262687 217989
rect 262715 217961 262749 217989
rect 262777 217961 262811 217989
rect 262839 217961 271625 217989
rect 271653 217961 271687 217989
rect 271715 217961 271749 217989
rect 271777 217961 271811 217989
rect 271839 217961 280625 217989
rect 280653 217961 280687 217989
rect 280715 217961 280749 217989
rect 280777 217961 280811 217989
rect 280839 217961 289625 217989
rect 289653 217961 289687 217989
rect 289715 217961 289749 217989
rect 289777 217961 289811 217989
rect 289839 217961 298248 217989
rect 298276 217961 298310 217989
rect 298338 217961 298372 217989
rect 298400 217961 298434 217989
rect 298462 217961 298990 217989
rect -958 217913 298990 217961
rect -958 212175 298990 212223
rect -958 212147 -910 212175
rect -882 212147 -848 212175
rect -820 212147 -786 212175
rect -758 212147 -724 212175
rect -696 212147 3485 212175
rect 3513 212147 3547 212175
rect 3575 212147 3609 212175
rect 3637 212147 3671 212175
rect 3699 212147 12485 212175
rect 12513 212147 12547 212175
rect 12575 212147 12609 212175
rect 12637 212147 12671 212175
rect 12699 212147 21485 212175
rect 21513 212147 21547 212175
rect 21575 212147 21609 212175
rect 21637 212147 21671 212175
rect 21699 212147 30485 212175
rect 30513 212147 30547 212175
rect 30575 212147 30609 212175
rect 30637 212147 30671 212175
rect 30699 212147 39485 212175
rect 39513 212147 39547 212175
rect 39575 212147 39609 212175
rect 39637 212147 39671 212175
rect 39699 212147 48485 212175
rect 48513 212147 48547 212175
rect 48575 212147 48609 212175
rect 48637 212147 48671 212175
rect 48699 212147 59939 212175
rect 59967 212147 60001 212175
rect 60029 212147 75299 212175
rect 75327 212147 75361 212175
rect 75389 212147 90659 212175
rect 90687 212147 90721 212175
rect 90749 212147 106019 212175
rect 106047 212147 106081 212175
rect 106109 212147 121379 212175
rect 121407 212147 121441 212175
rect 121469 212147 136739 212175
rect 136767 212147 136801 212175
rect 136829 212147 156485 212175
rect 156513 212147 156547 212175
rect 156575 212147 156609 212175
rect 156637 212147 156671 212175
rect 156699 212147 165485 212175
rect 165513 212147 165547 212175
rect 165575 212147 165609 212175
rect 165637 212147 165671 212175
rect 165699 212147 174485 212175
rect 174513 212147 174547 212175
rect 174575 212147 174609 212175
rect 174637 212147 174671 212175
rect 174699 212147 183485 212175
rect 183513 212147 183547 212175
rect 183575 212147 183609 212175
rect 183637 212147 183671 212175
rect 183699 212147 192485 212175
rect 192513 212147 192547 212175
rect 192575 212147 192609 212175
rect 192637 212147 192671 212175
rect 192699 212147 201485 212175
rect 201513 212147 201547 212175
rect 201575 212147 201609 212175
rect 201637 212147 201671 212175
rect 201699 212147 210485 212175
rect 210513 212147 210547 212175
rect 210575 212147 210609 212175
rect 210637 212147 210671 212175
rect 210699 212147 219485 212175
rect 219513 212147 219547 212175
rect 219575 212147 219609 212175
rect 219637 212147 219671 212175
rect 219699 212147 228485 212175
rect 228513 212147 228547 212175
rect 228575 212147 228609 212175
rect 228637 212147 228671 212175
rect 228699 212147 237485 212175
rect 237513 212147 237547 212175
rect 237575 212147 237609 212175
rect 237637 212147 237671 212175
rect 237699 212147 246485 212175
rect 246513 212147 246547 212175
rect 246575 212147 246609 212175
rect 246637 212147 246671 212175
rect 246699 212147 255485 212175
rect 255513 212147 255547 212175
rect 255575 212147 255609 212175
rect 255637 212147 255671 212175
rect 255699 212147 264485 212175
rect 264513 212147 264547 212175
rect 264575 212147 264609 212175
rect 264637 212147 264671 212175
rect 264699 212147 273485 212175
rect 273513 212147 273547 212175
rect 273575 212147 273609 212175
rect 273637 212147 273671 212175
rect 273699 212147 282485 212175
rect 282513 212147 282547 212175
rect 282575 212147 282609 212175
rect 282637 212147 282671 212175
rect 282699 212147 291485 212175
rect 291513 212147 291547 212175
rect 291575 212147 291609 212175
rect 291637 212147 291671 212175
rect 291699 212147 298728 212175
rect 298756 212147 298790 212175
rect 298818 212147 298852 212175
rect 298880 212147 298914 212175
rect 298942 212147 298990 212175
rect -958 212113 298990 212147
rect -958 212085 -910 212113
rect -882 212085 -848 212113
rect -820 212085 -786 212113
rect -758 212085 -724 212113
rect -696 212085 3485 212113
rect 3513 212085 3547 212113
rect 3575 212085 3609 212113
rect 3637 212085 3671 212113
rect 3699 212085 12485 212113
rect 12513 212085 12547 212113
rect 12575 212085 12609 212113
rect 12637 212085 12671 212113
rect 12699 212085 21485 212113
rect 21513 212085 21547 212113
rect 21575 212085 21609 212113
rect 21637 212085 21671 212113
rect 21699 212085 30485 212113
rect 30513 212085 30547 212113
rect 30575 212085 30609 212113
rect 30637 212085 30671 212113
rect 30699 212085 39485 212113
rect 39513 212085 39547 212113
rect 39575 212085 39609 212113
rect 39637 212085 39671 212113
rect 39699 212085 48485 212113
rect 48513 212085 48547 212113
rect 48575 212085 48609 212113
rect 48637 212085 48671 212113
rect 48699 212085 59939 212113
rect 59967 212085 60001 212113
rect 60029 212085 75299 212113
rect 75327 212085 75361 212113
rect 75389 212085 90659 212113
rect 90687 212085 90721 212113
rect 90749 212085 106019 212113
rect 106047 212085 106081 212113
rect 106109 212085 121379 212113
rect 121407 212085 121441 212113
rect 121469 212085 136739 212113
rect 136767 212085 136801 212113
rect 136829 212085 156485 212113
rect 156513 212085 156547 212113
rect 156575 212085 156609 212113
rect 156637 212085 156671 212113
rect 156699 212085 165485 212113
rect 165513 212085 165547 212113
rect 165575 212085 165609 212113
rect 165637 212085 165671 212113
rect 165699 212085 174485 212113
rect 174513 212085 174547 212113
rect 174575 212085 174609 212113
rect 174637 212085 174671 212113
rect 174699 212085 183485 212113
rect 183513 212085 183547 212113
rect 183575 212085 183609 212113
rect 183637 212085 183671 212113
rect 183699 212085 192485 212113
rect 192513 212085 192547 212113
rect 192575 212085 192609 212113
rect 192637 212085 192671 212113
rect 192699 212085 201485 212113
rect 201513 212085 201547 212113
rect 201575 212085 201609 212113
rect 201637 212085 201671 212113
rect 201699 212085 210485 212113
rect 210513 212085 210547 212113
rect 210575 212085 210609 212113
rect 210637 212085 210671 212113
rect 210699 212085 219485 212113
rect 219513 212085 219547 212113
rect 219575 212085 219609 212113
rect 219637 212085 219671 212113
rect 219699 212085 228485 212113
rect 228513 212085 228547 212113
rect 228575 212085 228609 212113
rect 228637 212085 228671 212113
rect 228699 212085 237485 212113
rect 237513 212085 237547 212113
rect 237575 212085 237609 212113
rect 237637 212085 237671 212113
rect 237699 212085 246485 212113
rect 246513 212085 246547 212113
rect 246575 212085 246609 212113
rect 246637 212085 246671 212113
rect 246699 212085 255485 212113
rect 255513 212085 255547 212113
rect 255575 212085 255609 212113
rect 255637 212085 255671 212113
rect 255699 212085 264485 212113
rect 264513 212085 264547 212113
rect 264575 212085 264609 212113
rect 264637 212085 264671 212113
rect 264699 212085 273485 212113
rect 273513 212085 273547 212113
rect 273575 212085 273609 212113
rect 273637 212085 273671 212113
rect 273699 212085 282485 212113
rect 282513 212085 282547 212113
rect 282575 212085 282609 212113
rect 282637 212085 282671 212113
rect 282699 212085 291485 212113
rect 291513 212085 291547 212113
rect 291575 212085 291609 212113
rect 291637 212085 291671 212113
rect 291699 212085 298728 212113
rect 298756 212085 298790 212113
rect 298818 212085 298852 212113
rect 298880 212085 298914 212113
rect 298942 212085 298990 212113
rect -958 212051 298990 212085
rect -958 212023 -910 212051
rect -882 212023 -848 212051
rect -820 212023 -786 212051
rect -758 212023 -724 212051
rect -696 212023 3485 212051
rect 3513 212023 3547 212051
rect 3575 212023 3609 212051
rect 3637 212023 3671 212051
rect 3699 212023 12485 212051
rect 12513 212023 12547 212051
rect 12575 212023 12609 212051
rect 12637 212023 12671 212051
rect 12699 212023 21485 212051
rect 21513 212023 21547 212051
rect 21575 212023 21609 212051
rect 21637 212023 21671 212051
rect 21699 212023 30485 212051
rect 30513 212023 30547 212051
rect 30575 212023 30609 212051
rect 30637 212023 30671 212051
rect 30699 212023 39485 212051
rect 39513 212023 39547 212051
rect 39575 212023 39609 212051
rect 39637 212023 39671 212051
rect 39699 212023 48485 212051
rect 48513 212023 48547 212051
rect 48575 212023 48609 212051
rect 48637 212023 48671 212051
rect 48699 212023 59939 212051
rect 59967 212023 60001 212051
rect 60029 212023 75299 212051
rect 75327 212023 75361 212051
rect 75389 212023 90659 212051
rect 90687 212023 90721 212051
rect 90749 212023 106019 212051
rect 106047 212023 106081 212051
rect 106109 212023 121379 212051
rect 121407 212023 121441 212051
rect 121469 212023 136739 212051
rect 136767 212023 136801 212051
rect 136829 212023 156485 212051
rect 156513 212023 156547 212051
rect 156575 212023 156609 212051
rect 156637 212023 156671 212051
rect 156699 212023 165485 212051
rect 165513 212023 165547 212051
rect 165575 212023 165609 212051
rect 165637 212023 165671 212051
rect 165699 212023 174485 212051
rect 174513 212023 174547 212051
rect 174575 212023 174609 212051
rect 174637 212023 174671 212051
rect 174699 212023 183485 212051
rect 183513 212023 183547 212051
rect 183575 212023 183609 212051
rect 183637 212023 183671 212051
rect 183699 212023 192485 212051
rect 192513 212023 192547 212051
rect 192575 212023 192609 212051
rect 192637 212023 192671 212051
rect 192699 212023 201485 212051
rect 201513 212023 201547 212051
rect 201575 212023 201609 212051
rect 201637 212023 201671 212051
rect 201699 212023 210485 212051
rect 210513 212023 210547 212051
rect 210575 212023 210609 212051
rect 210637 212023 210671 212051
rect 210699 212023 219485 212051
rect 219513 212023 219547 212051
rect 219575 212023 219609 212051
rect 219637 212023 219671 212051
rect 219699 212023 228485 212051
rect 228513 212023 228547 212051
rect 228575 212023 228609 212051
rect 228637 212023 228671 212051
rect 228699 212023 237485 212051
rect 237513 212023 237547 212051
rect 237575 212023 237609 212051
rect 237637 212023 237671 212051
rect 237699 212023 246485 212051
rect 246513 212023 246547 212051
rect 246575 212023 246609 212051
rect 246637 212023 246671 212051
rect 246699 212023 255485 212051
rect 255513 212023 255547 212051
rect 255575 212023 255609 212051
rect 255637 212023 255671 212051
rect 255699 212023 264485 212051
rect 264513 212023 264547 212051
rect 264575 212023 264609 212051
rect 264637 212023 264671 212051
rect 264699 212023 273485 212051
rect 273513 212023 273547 212051
rect 273575 212023 273609 212051
rect 273637 212023 273671 212051
rect 273699 212023 282485 212051
rect 282513 212023 282547 212051
rect 282575 212023 282609 212051
rect 282637 212023 282671 212051
rect 282699 212023 291485 212051
rect 291513 212023 291547 212051
rect 291575 212023 291609 212051
rect 291637 212023 291671 212051
rect 291699 212023 298728 212051
rect 298756 212023 298790 212051
rect 298818 212023 298852 212051
rect 298880 212023 298914 212051
rect 298942 212023 298990 212051
rect -958 211989 298990 212023
rect -958 211961 -910 211989
rect -882 211961 -848 211989
rect -820 211961 -786 211989
rect -758 211961 -724 211989
rect -696 211961 3485 211989
rect 3513 211961 3547 211989
rect 3575 211961 3609 211989
rect 3637 211961 3671 211989
rect 3699 211961 12485 211989
rect 12513 211961 12547 211989
rect 12575 211961 12609 211989
rect 12637 211961 12671 211989
rect 12699 211961 21485 211989
rect 21513 211961 21547 211989
rect 21575 211961 21609 211989
rect 21637 211961 21671 211989
rect 21699 211961 30485 211989
rect 30513 211961 30547 211989
rect 30575 211961 30609 211989
rect 30637 211961 30671 211989
rect 30699 211961 39485 211989
rect 39513 211961 39547 211989
rect 39575 211961 39609 211989
rect 39637 211961 39671 211989
rect 39699 211961 48485 211989
rect 48513 211961 48547 211989
rect 48575 211961 48609 211989
rect 48637 211961 48671 211989
rect 48699 211961 59939 211989
rect 59967 211961 60001 211989
rect 60029 211961 75299 211989
rect 75327 211961 75361 211989
rect 75389 211961 90659 211989
rect 90687 211961 90721 211989
rect 90749 211961 106019 211989
rect 106047 211961 106081 211989
rect 106109 211961 121379 211989
rect 121407 211961 121441 211989
rect 121469 211961 136739 211989
rect 136767 211961 136801 211989
rect 136829 211961 156485 211989
rect 156513 211961 156547 211989
rect 156575 211961 156609 211989
rect 156637 211961 156671 211989
rect 156699 211961 165485 211989
rect 165513 211961 165547 211989
rect 165575 211961 165609 211989
rect 165637 211961 165671 211989
rect 165699 211961 174485 211989
rect 174513 211961 174547 211989
rect 174575 211961 174609 211989
rect 174637 211961 174671 211989
rect 174699 211961 183485 211989
rect 183513 211961 183547 211989
rect 183575 211961 183609 211989
rect 183637 211961 183671 211989
rect 183699 211961 192485 211989
rect 192513 211961 192547 211989
rect 192575 211961 192609 211989
rect 192637 211961 192671 211989
rect 192699 211961 201485 211989
rect 201513 211961 201547 211989
rect 201575 211961 201609 211989
rect 201637 211961 201671 211989
rect 201699 211961 210485 211989
rect 210513 211961 210547 211989
rect 210575 211961 210609 211989
rect 210637 211961 210671 211989
rect 210699 211961 219485 211989
rect 219513 211961 219547 211989
rect 219575 211961 219609 211989
rect 219637 211961 219671 211989
rect 219699 211961 228485 211989
rect 228513 211961 228547 211989
rect 228575 211961 228609 211989
rect 228637 211961 228671 211989
rect 228699 211961 237485 211989
rect 237513 211961 237547 211989
rect 237575 211961 237609 211989
rect 237637 211961 237671 211989
rect 237699 211961 246485 211989
rect 246513 211961 246547 211989
rect 246575 211961 246609 211989
rect 246637 211961 246671 211989
rect 246699 211961 255485 211989
rect 255513 211961 255547 211989
rect 255575 211961 255609 211989
rect 255637 211961 255671 211989
rect 255699 211961 264485 211989
rect 264513 211961 264547 211989
rect 264575 211961 264609 211989
rect 264637 211961 264671 211989
rect 264699 211961 273485 211989
rect 273513 211961 273547 211989
rect 273575 211961 273609 211989
rect 273637 211961 273671 211989
rect 273699 211961 282485 211989
rect 282513 211961 282547 211989
rect 282575 211961 282609 211989
rect 282637 211961 282671 211989
rect 282699 211961 291485 211989
rect 291513 211961 291547 211989
rect 291575 211961 291609 211989
rect 291637 211961 291671 211989
rect 291699 211961 298728 211989
rect 298756 211961 298790 211989
rect 298818 211961 298852 211989
rect 298880 211961 298914 211989
rect 298942 211961 298990 211989
rect -958 211913 298990 211961
rect -958 209175 298990 209223
rect -958 209147 -430 209175
rect -402 209147 -368 209175
rect -340 209147 -306 209175
rect -278 209147 -244 209175
rect -216 209147 1625 209175
rect 1653 209147 1687 209175
rect 1715 209147 1749 209175
rect 1777 209147 1811 209175
rect 1839 209147 10625 209175
rect 10653 209147 10687 209175
rect 10715 209147 10749 209175
rect 10777 209147 10811 209175
rect 10839 209147 19625 209175
rect 19653 209147 19687 209175
rect 19715 209147 19749 209175
rect 19777 209147 19811 209175
rect 19839 209147 28625 209175
rect 28653 209147 28687 209175
rect 28715 209147 28749 209175
rect 28777 209147 28811 209175
rect 28839 209147 37625 209175
rect 37653 209147 37687 209175
rect 37715 209147 37749 209175
rect 37777 209147 37811 209175
rect 37839 209147 46625 209175
rect 46653 209147 46687 209175
rect 46715 209147 46749 209175
rect 46777 209147 46811 209175
rect 46839 209147 52259 209175
rect 52287 209147 52321 209175
rect 52349 209147 67619 209175
rect 67647 209147 67681 209175
rect 67709 209147 82979 209175
rect 83007 209147 83041 209175
rect 83069 209147 98339 209175
rect 98367 209147 98401 209175
rect 98429 209147 113699 209175
rect 113727 209147 113761 209175
rect 113789 209147 129059 209175
rect 129087 209147 129121 209175
rect 129149 209147 144419 209175
rect 144447 209147 144481 209175
rect 144509 209147 154625 209175
rect 154653 209147 154687 209175
rect 154715 209147 154749 209175
rect 154777 209147 154811 209175
rect 154839 209147 163625 209175
rect 163653 209147 163687 209175
rect 163715 209147 163749 209175
rect 163777 209147 163811 209175
rect 163839 209147 172625 209175
rect 172653 209147 172687 209175
rect 172715 209147 172749 209175
rect 172777 209147 172811 209175
rect 172839 209147 181625 209175
rect 181653 209147 181687 209175
rect 181715 209147 181749 209175
rect 181777 209147 181811 209175
rect 181839 209147 190625 209175
rect 190653 209147 190687 209175
rect 190715 209147 190749 209175
rect 190777 209147 190811 209175
rect 190839 209147 199625 209175
rect 199653 209147 199687 209175
rect 199715 209147 199749 209175
rect 199777 209147 199811 209175
rect 199839 209147 208625 209175
rect 208653 209147 208687 209175
rect 208715 209147 208749 209175
rect 208777 209147 208811 209175
rect 208839 209147 217625 209175
rect 217653 209147 217687 209175
rect 217715 209147 217749 209175
rect 217777 209147 217811 209175
rect 217839 209147 226625 209175
rect 226653 209147 226687 209175
rect 226715 209147 226749 209175
rect 226777 209147 226811 209175
rect 226839 209147 235625 209175
rect 235653 209147 235687 209175
rect 235715 209147 235749 209175
rect 235777 209147 235811 209175
rect 235839 209147 244625 209175
rect 244653 209147 244687 209175
rect 244715 209147 244749 209175
rect 244777 209147 244811 209175
rect 244839 209147 253625 209175
rect 253653 209147 253687 209175
rect 253715 209147 253749 209175
rect 253777 209147 253811 209175
rect 253839 209147 262625 209175
rect 262653 209147 262687 209175
rect 262715 209147 262749 209175
rect 262777 209147 262811 209175
rect 262839 209147 271625 209175
rect 271653 209147 271687 209175
rect 271715 209147 271749 209175
rect 271777 209147 271811 209175
rect 271839 209147 280625 209175
rect 280653 209147 280687 209175
rect 280715 209147 280749 209175
rect 280777 209147 280811 209175
rect 280839 209147 289625 209175
rect 289653 209147 289687 209175
rect 289715 209147 289749 209175
rect 289777 209147 289811 209175
rect 289839 209147 298248 209175
rect 298276 209147 298310 209175
rect 298338 209147 298372 209175
rect 298400 209147 298434 209175
rect 298462 209147 298990 209175
rect -958 209113 298990 209147
rect -958 209085 -430 209113
rect -402 209085 -368 209113
rect -340 209085 -306 209113
rect -278 209085 -244 209113
rect -216 209085 1625 209113
rect 1653 209085 1687 209113
rect 1715 209085 1749 209113
rect 1777 209085 1811 209113
rect 1839 209085 10625 209113
rect 10653 209085 10687 209113
rect 10715 209085 10749 209113
rect 10777 209085 10811 209113
rect 10839 209085 19625 209113
rect 19653 209085 19687 209113
rect 19715 209085 19749 209113
rect 19777 209085 19811 209113
rect 19839 209085 28625 209113
rect 28653 209085 28687 209113
rect 28715 209085 28749 209113
rect 28777 209085 28811 209113
rect 28839 209085 37625 209113
rect 37653 209085 37687 209113
rect 37715 209085 37749 209113
rect 37777 209085 37811 209113
rect 37839 209085 46625 209113
rect 46653 209085 46687 209113
rect 46715 209085 46749 209113
rect 46777 209085 46811 209113
rect 46839 209085 52259 209113
rect 52287 209085 52321 209113
rect 52349 209085 67619 209113
rect 67647 209085 67681 209113
rect 67709 209085 82979 209113
rect 83007 209085 83041 209113
rect 83069 209085 98339 209113
rect 98367 209085 98401 209113
rect 98429 209085 113699 209113
rect 113727 209085 113761 209113
rect 113789 209085 129059 209113
rect 129087 209085 129121 209113
rect 129149 209085 144419 209113
rect 144447 209085 144481 209113
rect 144509 209085 154625 209113
rect 154653 209085 154687 209113
rect 154715 209085 154749 209113
rect 154777 209085 154811 209113
rect 154839 209085 163625 209113
rect 163653 209085 163687 209113
rect 163715 209085 163749 209113
rect 163777 209085 163811 209113
rect 163839 209085 172625 209113
rect 172653 209085 172687 209113
rect 172715 209085 172749 209113
rect 172777 209085 172811 209113
rect 172839 209085 181625 209113
rect 181653 209085 181687 209113
rect 181715 209085 181749 209113
rect 181777 209085 181811 209113
rect 181839 209085 190625 209113
rect 190653 209085 190687 209113
rect 190715 209085 190749 209113
rect 190777 209085 190811 209113
rect 190839 209085 199625 209113
rect 199653 209085 199687 209113
rect 199715 209085 199749 209113
rect 199777 209085 199811 209113
rect 199839 209085 208625 209113
rect 208653 209085 208687 209113
rect 208715 209085 208749 209113
rect 208777 209085 208811 209113
rect 208839 209085 217625 209113
rect 217653 209085 217687 209113
rect 217715 209085 217749 209113
rect 217777 209085 217811 209113
rect 217839 209085 226625 209113
rect 226653 209085 226687 209113
rect 226715 209085 226749 209113
rect 226777 209085 226811 209113
rect 226839 209085 235625 209113
rect 235653 209085 235687 209113
rect 235715 209085 235749 209113
rect 235777 209085 235811 209113
rect 235839 209085 244625 209113
rect 244653 209085 244687 209113
rect 244715 209085 244749 209113
rect 244777 209085 244811 209113
rect 244839 209085 253625 209113
rect 253653 209085 253687 209113
rect 253715 209085 253749 209113
rect 253777 209085 253811 209113
rect 253839 209085 262625 209113
rect 262653 209085 262687 209113
rect 262715 209085 262749 209113
rect 262777 209085 262811 209113
rect 262839 209085 271625 209113
rect 271653 209085 271687 209113
rect 271715 209085 271749 209113
rect 271777 209085 271811 209113
rect 271839 209085 280625 209113
rect 280653 209085 280687 209113
rect 280715 209085 280749 209113
rect 280777 209085 280811 209113
rect 280839 209085 289625 209113
rect 289653 209085 289687 209113
rect 289715 209085 289749 209113
rect 289777 209085 289811 209113
rect 289839 209085 298248 209113
rect 298276 209085 298310 209113
rect 298338 209085 298372 209113
rect 298400 209085 298434 209113
rect 298462 209085 298990 209113
rect -958 209051 298990 209085
rect -958 209023 -430 209051
rect -402 209023 -368 209051
rect -340 209023 -306 209051
rect -278 209023 -244 209051
rect -216 209023 1625 209051
rect 1653 209023 1687 209051
rect 1715 209023 1749 209051
rect 1777 209023 1811 209051
rect 1839 209023 10625 209051
rect 10653 209023 10687 209051
rect 10715 209023 10749 209051
rect 10777 209023 10811 209051
rect 10839 209023 19625 209051
rect 19653 209023 19687 209051
rect 19715 209023 19749 209051
rect 19777 209023 19811 209051
rect 19839 209023 28625 209051
rect 28653 209023 28687 209051
rect 28715 209023 28749 209051
rect 28777 209023 28811 209051
rect 28839 209023 37625 209051
rect 37653 209023 37687 209051
rect 37715 209023 37749 209051
rect 37777 209023 37811 209051
rect 37839 209023 46625 209051
rect 46653 209023 46687 209051
rect 46715 209023 46749 209051
rect 46777 209023 46811 209051
rect 46839 209023 52259 209051
rect 52287 209023 52321 209051
rect 52349 209023 67619 209051
rect 67647 209023 67681 209051
rect 67709 209023 82979 209051
rect 83007 209023 83041 209051
rect 83069 209023 98339 209051
rect 98367 209023 98401 209051
rect 98429 209023 113699 209051
rect 113727 209023 113761 209051
rect 113789 209023 129059 209051
rect 129087 209023 129121 209051
rect 129149 209023 144419 209051
rect 144447 209023 144481 209051
rect 144509 209023 154625 209051
rect 154653 209023 154687 209051
rect 154715 209023 154749 209051
rect 154777 209023 154811 209051
rect 154839 209023 163625 209051
rect 163653 209023 163687 209051
rect 163715 209023 163749 209051
rect 163777 209023 163811 209051
rect 163839 209023 172625 209051
rect 172653 209023 172687 209051
rect 172715 209023 172749 209051
rect 172777 209023 172811 209051
rect 172839 209023 181625 209051
rect 181653 209023 181687 209051
rect 181715 209023 181749 209051
rect 181777 209023 181811 209051
rect 181839 209023 190625 209051
rect 190653 209023 190687 209051
rect 190715 209023 190749 209051
rect 190777 209023 190811 209051
rect 190839 209023 199625 209051
rect 199653 209023 199687 209051
rect 199715 209023 199749 209051
rect 199777 209023 199811 209051
rect 199839 209023 208625 209051
rect 208653 209023 208687 209051
rect 208715 209023 208749 209051
rect 208777 209023 208811 209051
rect 208839 209023 217625 209051
rect 217653 209023 217687 209051
rect 217715 209023 217749 209051
rect 217777 209023 217811 209051
rect 217839 209023 226625 209051
rect 226653 209023 226687 209051
rect 226715 209023 226749 209051
rect 226777 209023 226811 209051
rect 226839 209023 235625 209051
rect 235653 209023 235687 209051
rect 235715 209023 235749 209051
rect 235777 209023 235811 209051
rect 235839 209023 244625 209051
rect 244653 209023 244687 209051
rect 244715 209023 244749 209051
rect 244777 209023 244811 209051
rect 244839 209023 253625 209051
rect 253653 209023 253687 209051
rect 253715 209023 253749 209051
rect 253777 209023 253811 209051
rect 253839 209023 262625 209051
rect 262653 209023 262687 209051
rect 262715 209023 262749 209051
rect 262777 209023 262811 209051
rect 262839 209023 271625 209051
rect 271653 209023 271687 209051
rect 271715 209023 271749 209051
rect 271777 209023 271811 209051
rect 271839 209023 280625 209051
rect 280653 209023 280687 209051
rect 280715 209023 280749 209051
rect 280777 209023 280811 209051
rect 280839 209023 289625 209051
rect 289653 209023 289687 209051
rect 289715 209023 289749 209051
rect 289777 209023 289811 209051
rect 289839 209023 298248 209051
rect 298276 209023 298310 209051
rect 298338 209023 298372 209051
rect 298400 209023 298434 209051
rect 298462 209023 298990 209051
rect -958 208989 298990 209023
rect -958 208961 -430 208989
rect -402 208961 -368 208989
rect -340 208961 -306 208989
rect -278 208961 -244 208989
rect -216 208961 1625 208989
rect 1653 208961 1687 208989
rect 1715 208961 1749 208989
rect 1777 208961 1811 208989
rect 1839 208961 10625 208989
rect 10653 208961 10687 208989
rect 10715 208961 10749 208989
rect 10777 208961 10811 208989
rect 10839 208961 19625 208989
rect 19653 208961 19687 208989
rect 19715 208961 19749 208989
rect 19777 208961 19811 208989
rect 19839 208961 28625 208989
rect 28653 208961 28687 208989
rect 28715 208961 28749 208989
rect 28777 208961 28811 208989
rect 28839 208961 37625 208989
rect 37653 208961 37687 208989
rect 37715 208961 37749 208989
rect 37777 208961 37811 208989
rect 37839 208961 46625 208989
rect 46653 208961 46687 208989
rect 46715 208961 46749 208989
rect 46777 208961 46811 208989
rect 46839 208961 52259 208989
rect 52287 208961 52321 208989
rect 52349 208961 67619 208989
rect 67647 208961 67681 208989
rect 67709 208961 82979 208989
rect 83007 208961 83041 208989
rect 83069 208961 98339 208989
rect 98367 208961 98401 208989
rect 98429 208961 113699 208989
rect 113727 208961 113761 208989
rect 113789 208961 129059 208989
rect 129087 208961 129121 208989
rect 129149 208961 144419 208989
rect 144447 208961 144481 208989
rect 144509 208961 154625 208989
rect 154653 208961 154687 208989
rect 154715 208961 154749 208989
rect 154777 208961 154811 208989
rect 154839 208961 163625 208989
rect 163653 208961 163687 208989
rect 163715 208961 163749 208989
rect 163777 208961 163811 208989
rect 163839 208961 172625 208989
rect 172653 208961 172687 208989
rect 172715 208961 172749 208989
rect 172777 208961 172811 208989
rect 172839 208961 181625 208989
rect 181653 208961 181687 208989
rect 181715 208961 181749 208989
rect 181777 208961 181811 208989
rect 181839 208961 190625 208989
rect 190653 208961 190687 208989
rect 190715 208961 190749 208989
rect 190777 208961 190811 208989
rect 190839 208961 199625 208989
rect 199653 208961 199687 208989
rect 199715 208961 199749 208989
rect 199777 208961 199811 208989
rect 199839 208961 208625 208989
rect 208653 208961 208687 208989
rect 208715 208961 208749 208989
rect 208777 208961 208811 208989
rect 208839 208961 217625 208989
rect 217653 208961 217687 208989
rect 217715 208961 217749 208989
rect 217777 208961 217811 208989
rect 217839 208961 226625 208989
rect 226653 208961 226687 208989
rect 226715 208961 226749 208989
rect 226777 208961 226811 208989
rect 226839 208961 235625 208989
rect 235653 208961 235687 208989
rect 235715 208961 235749 208989
rect 235777 208961 235811 208989
rect 235839 208961 244625 208989
rect 244653 208961 244687 208989
rect 244715 208961 244749 208989
rect 244777 208961 244811 208989
rect 244839 208961 253625 208989
rect 253653 208961 253687 208989
rect 253715 208961 253749 208989
rect 253777 208961 253811 208989
rect 253839 208961 262625 208989
rect 262653 208961 262687 208989
rect 262715 208961 262749 208989
rect 262777 208961 262811 208989
rect 262839 208961 271625 208989
rect 271653 208961 271687 208989
rect 271715 208961 271749 208989
rect 271777 208961 271811 208989
rect 271839 208961 280625 208989
rect 280653 208961 280687 208989
rect 280715 208961 280749 208989
rect 280777 208961 280811 208989
rect 280839 208961 289625 208989
rect 289653 208961 289687 208989
rect 289715 208961 289749 208989
rect 289777 208961 289811 208989
rect 289839 208961 298248 208989
rect 298276 208961 298310 208989
rect 298338 208961 298372 208989
rect 298400 208961 298434 208989
rect 298462 208961 298990 208989
rect -958 208913 298990 208961
rect -958 203175 298990 203223
rect -958 203147 -910 203175
rect -882 203147 -848 203175
rect -820 203147 -786 203175
rect -758 203147 -724 203175
rect -696 203147 3485 203175
rect 3513 203147 3547 203175
rect 3575 203147 3609 203175
rect 3637 203147 3671 203175
rect 3699 203147 12485 203175
rect 12513 203147 12547 203175
rect 12575 203147 12609 203175
rect 12637 203147 12671 203175
rect 12699 203147 21485 203175
rect 21513 203147 21547 203175
rect 21575 203147 21609 203175
rect 21637 203147 21671 203175
rect 21699 203147 30485 203175
rect 30513 203147 30547 203175
rect 30575 203147 30609 203175
rect 30637 203147 30671 203175
rect 30699 203147 39485 203175
rect 39513 203147 39547 203175
rect 39575 203147 39609 203175
rect 39637 203147 39671 203175
rect 39699 203147 48485 203175
rect 48513 203147 48547 203175
rect 48575 203147 48609 203175
rect 48637 203147 48671 203175
rect 48699 203147 59939 203175
rect 59967 203147 60001 203175
rect 60029 203147 75299 203175
rect 75327 203147 75361 203175
rect 75389 203147 90659 203175
rect 90687 203147 90721 203175
rect 90749 203147 106019 203175
rect 106047 203147 106081 203175
rect 106109 203147 121379 203175
rect 121407 203147 121441 203175
rect 121469 203147 136739 203175
rect 136767 203147 136801 203175
rect 136829 203147 156485 203175
rect 156513 203147 156547 203175
rect 156575 203147 156609 203175
rect 156637 203147 156671 203175
rect 156699 203147 165485 203175
rect 165513 203147 165547 203175
rect 165575 203147 165609 203175
rect 165637 203147 165671 203175
rect 165699 203147 174485 203175
rect 174513 203147 174547 203175
rect 174575 203147 174609 203175
rect 174637 203147 174671 203175
rect 174699 203147 183485 203175
rect 183513 203147 183547 203175
rect 183575 203147 183609 203175
rect 183637 203147 183671 203175
rect 183699 203147 192485 203175
rect 192513 203147 192547 203175
rect 192575 203147 192609 203175
rect 192637 203147 192671 203175
rect 192699 203147 201485 203175
rect 201513 203147 201547 203175
rect 201575 203147 201609 203175
rect 201637 203147 201671 203175
rect 201699 203147 210485 203175
rect 210513 203147 210547 203175
rect 210575 203147 210609 203175
rect 210637 203147 210671 203175
rect 210699 203147 219485 203175
rect 219513 203147 219547 203175
rect 219575 203147 219609 203175
rect 219637 203147 219671 203175
rect 219699 203147 228485 203175
rect 228513 203147 228547 203175
rect 228575 203147 228609 203175
rect 228637 203147 228671 203175
rect 228699 203147 237485 203175
rect 237513 203147 237547 203175
rect 237575 203147 237609 203175
rect 237637 203147 237671 203175
rect 237699 203147 246485 203175
rect 246513 203147 246547 203175
rect 246575 203147 246609 203175
rect 246637 203147 246671 203175
rect 246699 203147 255485 203175
rect 255513 203147 255547 203175
rect 255575 203147 255609 203175
rect 255637 203147 255671 203175
rect 255699 203147 264485 203175
rect 264513 203147 264547 203175
rect 264575 203147 264609 203175
rect 264637 203147 264671 203175
rect 264699 203147 273485 203175
rect 273513 203147 273547 203175
rect 273575 203147 273609 203175
rect 273637 203147 273671 203175
rect 273699 203147 282485 203175
rect 282513 203147 282547 203175
rect 282575 203147 282609 203175
rect 282637 203147 282671 203175
rect 282699 203147 291485 203175
rect 291513 203147 291547 203175
rect 291575 203147 291609 203175
rect 291637 203147 291671 203175
rect 291699 203147 298728 203175
rect 298756 203147 298790 203175
rect 298818 203147 298852 203175
rect 298880 203147 298914 203175
rect 298942 203147 298990 203175
rect -958 203113 298990 203147
rect -958 203085 -910 203113
rect -882 203085 -848 203113
rect -820 203085 -786 203113
rect -758 203085 -724 203113
rect -696 203085 3485 203113
rect 3513 203085 3547 203113
rect 3575 203085 3609 203113
rect 3637 203085 3671 203113
rect 3699 203085 12485 203113
rect 12513 203085 12547 203113
rect 12575 203085 12609 203113
rect 12637 203085 12671 203113
rect 12699 203085 21485 203113
rect 21513 203085 21547 203113
rect 21575 203085 21609 203113
rect 21637 203085 21671 203113
rect 21699 203085 30485 203113
rect 30513 203085 30547 203113
rect 30575 203085 30609 203113
rect 30637 203085 30671 203113
rect 30699 203085 39485 203113
rect 39513 203085 39547 203113
rect 39575 203085 39609 203113
rect 39637 203085 39671 203113
rect 39699 203085 48485 203113
rect 48513 203085 48547 203113
rect 48575 203085 48609 203113
rect 48637 203085 48671 203113
rect 48699 203085 59939 203113
rect 59967 203085 60001 203113
rect 60029 203085 75299 203113
rect 75327 203085 75361 203113
rect 75389 203085 90659 203113
rect 90687 203085 90721 203113
rect 90749 203085 106019 203113
rect 106047 203085 106081 203113
rect 106109 203085 121379 203113
rect 121407 203085 121441 203113
rect 121469 203085 136739 203113
rect 136767 203085 136801 203113
rect 136829 203085 156485 203113
rect 156513 203085 156547 203113
rect 156575 203085 156609 203113
rect 156637 203085 156671 203113
rect 156699 203085 165485 203113
rect 165513 203085 165547 203113
rect 165575 203085 165609 203113
rect 165637 203085 165671 203113
rect 165699 203085 174485 203113
rect 174513 203085 174547 203113
rect 174575 203085 174609 203113
rect 174637 203085 174671 203113
rect 174699 203085 183485 203113
rect 183513 203085 183547 203113
rect 183575 203085 183609 203113
rect 183637 203085 183671 203113
rect 183699 203085 192485 203113
rect 192513 203085 192547 203113
rect 192575 203085 192609 203113
rect 192637 203085 192671 203113
rect 192699 203085 201485 203113
rect 201513 203085 201547 203113
rect 201575 203085 201609 203113
rect 201637 203085 201671 203113
rect 201699 203085 210485 203113
rect 210513 203085 210547 203113
rect 210575 203085 210609 203113
rect 210637 203085 210671 203113
rect 210699 203085 219485 203113
rect 219513 203085 219547 203113
rect 219575 203085 219609 203113
rect 219637 203085 219671 203113
rect 219699 203085 228485 203113
rect 228513 203085 228547 203113
rect 228575 203085 228609 203113
rect 228637 203085 228671 203113
rect 228699 203085 237485 203113
rect 237513 203085 237547 203113
rect 237575 203085 237609 203113
rect 237637 203085 237671 203113
rect 237699 203085 246485 203113
rect 246513 203085 246547 203113
rect 246575 203085 246609 203113
rect 246637 203085 246671 203113
rect 246699 203085 255485 203113
rect 255513 203085 255547 203113
rect 255575 203085 255609 203113
rect 255637 203085 255671 203113
rect 255699 203085 264485 203113
rect 264513 203085 264547 203113
rect 264575 203085 264609 203113
rect 264637 203085 264671 203113
rect 264699 203085 273485 203113
rect 273513 203085 273547 203113
rect 273575 203085 273609 203113
rect 273637 203085 273671 203113
rect 273699 203085 282485 203113
rect 282513 203085 282547 203113
rect 282575 203085 282609 203113
rect 282637 203085 282671 203113
rect 282699 203085 291485 203113
rect 291513 203085 291547 203113
rect 291575 203085 291609 203113
rect 291637 203085 291671 203113
rect 291699 203085 298728 203113
rect 298756 203085 298790 203113
rect 298818 203085 298852 203113
rect 298880 203085 298914 203113
rect 298942 203085 298990 203113
rect -958 203051 298990 203085
rect -958 203023 -910 203051
rect -882 203023 -848 203051
rect -820 203023 -786 203051
rect -758 203023 -724 203051
rect -696 203023 3485 203051
rect 3513 203023 3547 203051
rect 3575 203023 3609 203051
rect 3637 203023 3671 203051
rect 3699 203023 12485 203051
rect 12513 203023 12547 203051
rect 12575 203023 12609 203051
rect 12637 203023 12671 203051
rect 12699 203023 21485 203051
rect 21513 203023 21547 203051
rect 21575 203023 21609 203051
rect 21637 203023 21671 203051
rect 21699 203023 30485 203051
rect 30513 203023 30547 203051
rect 30575 203023 30609 203051
rect 30637 203023 30671 203051
rect 30699 203023 39485 203051
rect 39513 203023 39547 203051
rect 39575 203023 39609 203051
rect 39637 203023 39671 203051
rect 39699 203023 48485 203051
rect 48513 203023 48547 203051
rect 48575 203023 48609 203051
rect 48637 203023 48671 203051
rect 48699 203023 59939 203051
rect 59967 203023 60001 203051
rect 60029 203023 75299 203051
rect 75327 203023 75361 203051
rect 75389 203023 90659 203051
rect 90687 203023 90721 203051
rect 90749 203023 106019 203051
rect 106047 203023 106081 203051
rect 106109 203023 121379 203051
rect 121407 203023 121441 203051
rect 121469 203023 136739 203051
rect 136767 203023 136801 203051
rect 136829 203023 156485 203051
rect 156513 203023 156547 203051
rect 156575 203023 156609 203051
rect 156637 203023 156671 203051
rect 156699 203023 165485 203051
rect 165513 203023 165547 203051
rect 165575 203023 165609 203051
rect 165637 203023 165671 203051
rect 165699 203023 174485 203051
rect 174513 203023 174547 203051
rect 174575 203023 174609 203051
rect 174637 203023 174671 203051
rect 174699 203023 183485 203051
rect 183513 203023 183547 203051
rect 183575 203023 183609 203051
rect 183637 203023 183671 203051
rect 183699 203023 192485 203051
rect 192513 203023 192547 203051
rect 192575 203023 192609 203051
rect 192637 203023 192671 203051
rect 192699 203023 201485 203051
rect 201513 203023 201547 203051
rect 201575 203023 201609 203051
rect 201637 203023 201671 203051
rect 201699 203023 210485 203051
rect 210513 203023 210547 203051
rect 210575 203023 210609 203051
rect 210637 203023 210671 203051
rect 210699 203023 219485 203051
rect 219513 203023 219547 203051
rect 219575 203023 219609 203051
rect 219637 203023 219671 203051
rect 219699 203023 228485 203051
rect 228513 203023 228547 203051
rect 228575 203023 228609 203051
rect 228637 203023 228671 203051
rect 228699 203023 237485 203051
rect 237513 203023 237547 203051
rect 237575 203023 237609 203051
rect 237637 203023 237671 203051
rect 237699 203023 246485 203051
rect 246513 203023 246547 203051
rect 246575 203023 246609 203051
rect 246637 203023 246671 203051
rect 246699 203023 255485 203051
rect 255513 203023 255547 203051
rect 255575 203023 255609 203051
rect 255637 203023 255671 203051
rect 255699 203023 264485 203051
rect 264513 203023 264547 203051
rect 264575 203023 264609 203051
rect 264637 203023 264671 203051
rect 264699 203023 273485 203051
rect 273513 203023 273547 203051
rect 273575 203023 273609 203051
rect 273637 203023 273671 203051
rect 273699 203023 282485 203051
rect 282513 203023 282547 203051
rect 282575 203023 282609 203051
rect 282637 203023 282671 203051
rect 282699 203023 291485 203051
rect 291513 203023 291547 203051
rect 291575 203023 291609 203051
rect 291637 203023 291671 203051
rect 291699 203023 298728 203051
rect 298756 203023 298790 203051
rect 298818 203023 298852 203051
rect 298880 203023 298914 203051
rect 298942 203023 298990 203051
rect -958 202989 298990 203023
rect -958 202961 -910 202989
rect -882 202961 -848 202989
rect -820 202961 -786 202989
rect -758 202961 -724 202989
rect -696 202961 3485 202989
rect 3513 202961 3547 202989
rect 3575 202961 3609 202989
rect 3637 202961 3671 202989
rect 3699 202961 12485 202989
rect 12513 202961 12547 202989
rect 12575 202961 12609 202989
rect 12637 202961 12671 202989
rect 12699 202961 21485 202989
rect 21513 202961 21547 202989
rect 21575 202961 21609 202989
rect 21637 202961 21671 202989
rect 21699 202961 30485 202989
rect 30513 202961 30547 202989
rect 30575 202961 30609 202989
rect 30637 202961 30671 202989
rect 30699 202961 39485 202989
rect 39513 202961 39547 202989
rect 39575 202961 39609 202989
rect 39637 202961 39671 202989
rect 39699 202961 48485 202989
rect 48513 202961 48547 202989
rect 48575 202961 48609 202989
rect 48637 202961 48671 202989
rect 48699 202961 59939 202989
rect 59967 202961 60001 202989
rect 60029 202961 75299 202989
rect 75327 202961 75361 202989
rect 75389 202961 90659 202989
rect 90687 202961 90721 202989
rect 90749 202961 106019 202989
rect 106047 202961 106081 202989
rect 106109 202961 121379 202989
rect 121407 202961 121441 202989
rect 121469 202961 136739 202989
rect 136767 202961 136801 202989
rect 136829 202961 156485 202989
rect 156513 202961 156547 202989
rect 156575 202961 156609 202989
rect 156637 202961 156671 202989
rect 156699 202961 165485 202989
rect 165513 202961 165547 202989
rect 165575 202961 165609 202989
rect 165637 202961 165671 202989
rect 165699 202961 174485 202989
rect 174513 202961 174547 202989
rect 174575 202961 174609 202989
rect 174637 202961 174671 202989
rect 174699 202961 183485 202989
rect 183513 202961 183547 202989
rect 183575 202961 183609 202989
rect 183637 202961 183671 202989
rect 183699 202961 192485 202989
rect 192513 202961 192547 202989
rect 192575 202961 192609 202989
rect 192637 202961 192671 202989
rect 192699 202961 201485 202989
rect 201513 202961 201547 202989
rect 201575 202961 201609 202989
rect 201637 202961 201671 202989
rect 201699 202961 210485 202989
rect 210513 202961 210547 202989
rect 210575 202961 210609 202989
rect 210637 202961 210671 202989
rect 210699 202961 219485 202989
rect 219513 202961 219547 202989
rect 219575 202961 219609 202989
rect 219637 202961 219671 202989
rect 219699 202961 228485 202989
rect 228513 202961 228547 202989
rect 228575 202961 228609 202989
rect 228637 202961 228671 202989
rect 228699 202961 237485 202989
rect 237513 202961 237547 202989
rect 237575 202961 237609 202989
rect 237637 202961 237671 202989
rect 237699 202961 246485 202989
rect 246513 202961 246547 202989
rect 246575 202961 246609 202989
rect 246637 202961 246671 202989
rect 246699 202961 255485 202989
rect 255513 202961 255547 202989
rect 255575 202961 255609 202989
rect 255637 202961 255671 202989
rect 255699 202961 264485 202989
rect 264513 202961 264547 202989
rect 264575 202961 264609 202989
rect 264637 202961 264671 202989
rect 264699 202961 273485 202989
rect 273513 202961 273547 202989
rect 273575 202961 273609 202989
rect 273637 202961 273671 202989
rect 273699 202961 282485 202989
rect 282513 202961 282547 202989
rect 282575 202961 282609 202989
rect 282637 202961 282671 202989
rect 282699 202961 291485 202989
rect 291513 202961 291547 202989
rect 291575 202961 291609 202989
rect 291637 202961 291671 202989
rect 291699 202961 298728 202989
rect 298756 202961 298790 202989
rect 298818 202961 298852 202989
rect 298880 202961 298914 202989
rect 298942 202961 298990 202989
rect -958 202913 298990 202961
rect -958 200175 298990 200223
rect -958 200147 -430 200175
rect -402 200147 -368 200175
rect -340 200147 -306 200175
rect -278 200147 -244 200175
rect -216 200147 1625 200175
rect 1653 200147 1687 200175
rect 1715 200147 1749 200175
rect 1777 200147 1811 200175
rect 1839 200147 10625 200175
rect 10653 200147 10687 200175
rect 10715 200147 10749 200175
rect 10777 200147 10811 200175
rect 10839 200147 19625 200175
rect 19653 200147 19687 200175
rect 19715 200147 19749 200175
rect 19777 200147 19811 200175
rect 19839 200147 28625 200175
rect 28653 200147 28687 200175
rect 28715 200147 28749 200175
rect 28777 200147 28811 200175
rect 28839 200147 37625 200175
rect 37653 200147 37687 200175
rect 37715 200147 37749 200175
rect 37777 200147 37811 200175
rect 37839 200147 46625 200175
rect 46653 200147 46687 200175
rect 46715 200147 46749 200175
rect 46777 200147 46811 200175
rect 46839 200147 154625 200175
rect 154653 200147 154687 200175
rect 154715 200147 154749 200175
rect 154777 200147 154811 200175
rect 154839 200147 163625 200175
rect 163653 200147 163687 200175
rect 163715 200147 163749 200175
rect 163777 200147 163811 200175
rect 163839 200147 172625 200175
rect 172653 200147 172687 200175
rect 172715 200147 172749 200175
rect 172777 200147 172811 200175
rect 172839 200147 181625 200175
rect 181653 200147 181687 200175
rect 181715 200147 181749 200175
rect 181777 200147 181811 200175
rect 181839 200147 190625 200175
rect 190653 200147 190687 200175
rect 190715 200147 190749 200175
rect 190777 200147 190811 200175
rect 190839 200147 199625 200175
rect 199653 200147 199687 200175
rect 199715 200147 199749 200175
rect 199777 200147 199811 200175
rect 199839 200147 208625 200175
rect 208653 200147 208687 200175
rect 208715 200147 208749 200175
rect 208777 200147 208811 200175
rect 208839 200147 217625 200175
rect 217653 200147 217687 200175
rect 217715 200147 217749 200175
rect 217777 200147 217811 200175
rect 217839 200147 226625 200175
rect 226653 200147 226687 200175
rect 226715 200147 226749 200175
rect 226777 200147 226811 200175
rect 226839 200147 235625 200175
rect 235653 200147 235687 200175
rect 235715 200147 235749 200175
rect 235777 200147 235811 200175
rect 235839 200147 244625 200175
rect 244653 200147 244687 200175
rect 244715 200147 244749 200175
rect 244777 200147 244811 200175
rect 244839 200147 253625 200175
rect 253653 200147 253687 200175
rect 253715 200147 253749 200175
rect 253777 200147 253811 200175
rect 253839 200147 262625 200175
rect 262653 200147 262687 200175
rect 262715 200147 262749 200175
rect 262777 200147 262811 200175
rect 262839 200147 271625 200175
rect 271653 200147 271687 200175
rect 271715 200147 271749 200175
rect 271777 200147 271811 200175
rect 271839 200147 280625 200175
rect 280653 200147 280687 200175
rect 280715 200147 280749 200175
rect 280777 200147 280811 200175
rect 280839 200147 289625 200175
rect 289653 200147 289687 200175
rect 289715 200147 289749 200175
rect 289777 200147 289811 200175
rect 289839 200147 298248 200175
rect 298276 200147 298310 200175
rect 298338 200147 298372 200175
rect 298400 200147 298434 200175
rect 298462 200147 298990 200175
rect -958 200113 298990 200147
rect -958 200085 -430 200113
rect -402 200085 -368 200113
rect -340 200085 -306 200113
rect -278 200085 -244 200113
rect -216 200085 1625 200113
rect 1653 200085 1687 200113
rect 1715 200085 1749 200113
rect 1777 200085 1811 200113
rect 1839 200085 10625 200113
rect 10653 200085 10687 200113
rect 10715 200085 10749 200113
rect 10777 200085 10811 200113
rect 10839 200085 19625 200113
rect 19653 200085 19687 200113
rect 19715 200085 19749 200113
rect 19777 200085 19811 200113
rect 19839 200085 28625 200113
rect 28653 200085 28687 200113
rect 28715 200085 28749 200113
rect 28777 200085 28811 200113
rect 28839 200085 37625 200113
rect 37653 200085 37687 200113
rect 37715 200085 37749 200113
rect 37777 200085 37811 200113
rect 37839 200085 46625 200113
rect 46653 200085 46687 200113
rect 46715 200085 46749 200113
rect 46777 200085 46811 200113
rect 46839 200085 154625 200113
rect 154653 200085 154687 200113
rect 154715 200085 154749 200113
rect 154777 200085 154811 200113
rect 154839 200085 163625 200113
rect 163653 200085 163687 200113
rect 163715 200085 163749 200113
rect 163777 200085 163811 200113
rect 163839 200085 172625 200113
rect 172653 200085 172687 200113
rect 172715 200085 172749 200113
rect 172777 200085 172811 200113
rect 172839 200085 181625 200113
rect 181653 200085 181687 200113
rect 181715 200085 181749 200113
rect 181777 200085 181811 200113
rect 181839 200085 190625 200113
rect 190653 200085 190687 200113
rect 190715 200085 190749 200113
rect 190777 200085 190811 200113
rect 190839 200085 199625 200113
rect 199653 200085 199687 200113
rect 199715 200085 199749 200113
rect 199777 200085 199811 200113
rect 199839 200085 208625 200113
rect 208653 200085 208687 200113
rect 208715 200085 208749 200113
rect 208777 200085 208811 200113
rect 208839 200085 217625 200113
rect 217653 200085 217687 200113
rect 217715 200085 217749 200113
rect 217777 200085 217811 200113
rect 217839 200085 226625 200113
rect 226653 200085 226687 200113
rect 226715 200085 226749 200113
rect 226777 200085 226811 200113
rect 226839 200085 235625 200113
rect 235653 200085 235687 200113
rect 235715 200085 235749 200113
rect 235777 200085 235811 200113
rect 235839 200085 244625 200113
rect 244653 200085 244687 200113
rect 244715 200085 244749 200113
rect 244777 200085 244811 200113
rect 244839 200085 253625 200113
rect 253653 200085 253687 200113
rect 253715 200085 253749 200113
rect 253777 200085 253811 200113
rect 253839 200085 262625 200113
rect 262653 200085 262687 200113
rect 262715 200085 262749 200113
rect 262777 200085 262811 200113
rect 262839 200085 271625 200113
rect 271653 200085 271687 200113
rect 271715 200085 271749 200113
rect 271777 200085 271811 200113
rect 271839 200085 280625 200113
rect 280653 200085 280687 200113
rect 280715 200085 280749 200113
rect 280777 200085 280811 200113
rect 280839 200085 289625 200113
rect 289653 200085 289687 200113
rect 289715 200085 289749 200113
rect 289777 200085 289811 200113
rect 289839 200085 298248 200113
rect 298276 200085 298310 200113
rect 298338 200085 298372 200113
rect 298400 200085 298434 200113
rect 298462 200085 298990 200113
rect -958 200051 298990 200085
rect -958 200023 -430 200051
rect -402 200023 -368 200051
rect -340 200023 -306 200051
rect -278 200023 -244 200051
rect -216 200023 1625 200051
rect 1653 200023 1687 200051
rect 1715 200023 1749 200051
rect 1777 200023 1811 200051
rect 1839 200023 10625 200051
rect 10653 200023 10687 200051
rect 10715 200023 10749 200051
rect 10777 200023 10811 200051
rect 10839 200023 19625 200051
rect 19653 200023 19687 200051
rect 19715 200023 19749 200051
rect 19777 200023 19811 200051
rect 19839 200023 28625 200051
rect 28653 200023 28687 200051
rect 28715 200023 28749 200051
rect 28777 200023 28811 200051
rect 28839 200023 37625 200051
rect 37653 200023 37687 200051
rect 37715 200023 37749 200051
rect 37777 200023 37811 200051
rect 37839 200023 46625 200051
rect 46653 200023 46687 200051
rect 46715 200023 46749 200051
rect 46777 200023 46811 200051
rect 46839 200023 154625 200051
rect 154653 200023 154687 200051
rect 154715 200023 154749 200051
rect 154777 200023 154811 200051
rect 154839 200023 163625 200051
rect 163653 200023 163687 200051
rect 163715 200023 163749 200051
rect 163777 200023 163811 200051
rect 163839 200023 172625 200051
rect 172653 200023 172687 200051
rect 172715 200023 172749 200051
rect 172777 200023 172811 200051
rect 172839 200023 181625 200051
rect 181653 200023 181687 200051
rect 181715 200023 181749 200051
rect 181777 200023 181811 200051
rect 181839 200023 190625 200051
rect 190653 200023 190687 200051
rect 190715 200023 190749 200051
rect 190777 200023 190811 200051
rect 190839 200023 199625 200051
rect 199653 200023 199687 200051
rect 199715 200023 199749 200051
rect 199777 200023 199811 200051
rect 199839 200023 208625 200051
rect 208653 200023 208687 200051
rect 208715 200023 208749 200051
rect 208777 200023 208811 200051
rect 208839 200023 217625 200051
rect 217653 200023 217687 200051
rect 217715 200023 217749 200051
rect 217777 200023 217811 200051
rect 217839 200023 226625 200051
rect 226653 200023 226687 200051
rect 226715 200023 226749 200051
rect 226777 200023 226811 200051
rect 226839 200023 235625 200051
rect 235653 200023 235687 200051
rect 235715 200023 235749 200051
rect 235777 200023 235811 200051
rect 235839 200023 244625 200051
rect 244653 200023 244687 200051
rect 244715 200023 244749 200051
rect 244777 200023 244811 200051
rect 244839 200023 253625 200051
rect 253653 200023 253687 200051
rect 253715 200023 253749 200051
rect 253777 200023 253811 200051
rect 253839 200023 262625 200051
rect 262653 200023 262687 200051
rect 262715 200023 262749 200051
rect 262777 200023 262811 200051
rect 262839 200023 271625 200051
rect 271653 200023 271687 200051
rect 271715 200023 271749 200051
rect 271777 200023 271811 200051
rect 271839 200023 280625 200051
rect 280653 200023 280687 200051
rect 280715 200023 280749 200051
rect 280777 200023 280811 200051
rect 280839 200023 289625 200051
rect 289653 200023 289687 200051
rect 289715 200023 289749 200051
rect 289777 200023 289811 200051
rect 289839 200023 298248 200051
rect 298276 200023 298310 200051
rect 298338 200023 298372 200051
rect 298400 200023 298434 200051
rect 298462 200023 298990 200051
rect -958 199989 298990 200023
rect -958 199961 -430 199989
rect -402 199961 -368 199989
rect -340 199961 -306 199989
rect -278 199961 -244 199989
rect -216 199961 1625 199989
rect 1653 199961 1687 199989
rect 1715 199961 1749 199989
rect 1777 199961 1811 199989
rect 1839 199961 10625 199989
rect 10653 199961 10687 199989
rect 10715 199961 10749 199989
rect 10777 199961 10811 199989
rect 10839 199961 19625 199989
rect 19653 199961 19687 199989
rect 19715 199961 19749 199989
rect 19777 199961 19811 199989
rect 19839 199961 28625 199989
rect 28653 199961 28687 199989
rect 28715 199961 28749 199989
rect 28777 199961 28811 199989
rect 28839 199961 37625 199989
rect 37653 199961 37687 199989
rect 37715 199961 37749 199989
rect 37777 199961 37811 199989
rect 37839 199961 46625 199989
rect 46653 199961 46687 199989
rect 46715 199961 46749 199989
rect 46777 199961 46811 199989
rect 46839 199961 154625 199989
rect 154653 199961 154687 199989
rect 154715 199961 154749 199989
rect 154777 199961 154811 199989
rect 154839 199961 163625 199989
rect 163653 199961 163687 199989
rect 163715 199961 163749 199989
rect 163777 199961 163811 199989
rect 163839 199961 172625 199989
rect 172653 199961 172687 199989
rect 172715 199961 172749 199989
rect 172777 199961 172811 199989
rect 172839 199961 181625 199989
rect 181653 199961 181687 199989
rect 181715 199961 181749 199989
rect 181777 199961 181811 199989
rect 181839 199961 190625 199989
rect 190653 199961 190687 199989
rect 190715 199961 190749 199989
rect 190777 199961 190811 199989
rect 190839 199961 199625 199989
rect 199653 199961 199687 199989
rect 199715 199961 199749 199989
rect 199777 199961 199811 199989
rect 199839 199961 208625 199989
rect 208653 199961 208687 199989
rect 208715 199961 208749 199989
rect 208777 199961 208811 199989
rect 208839 199961 217625 199989
rect 217653 199961 217687 199989
rect 217715 199961 217749 199989
rect 217777 199961 217811 199989
rect 217839 199961 226625 199989
rect 226653 199961 226687 199989
rect 226715 199961 226749 199989
rect 226777 199961 226811 199989
rect 226839 199961 235625 199989
rect 235653 199961 235687 199989
rect 235715 199961 235749 199989
rect 235777 199961 235811 199989
rect 235839 199961 244625 199989
rect 244653 199961 244687 199989
rect 244715 199961 244749 199989
rect 244777 199961 244811 199989
rect 244839 199961 253625 199989
rect 253653 199961 253687 199989
rect 253715 199961 253749 199989
rect 253777 199961 253811 199989
rect 253839 199961 262625 199989
rect 262653 199961 262687 199989
rect 262715 199961 262749 199989
rect 262777 199961 262811 199989
rect 262839 199961 271625 199989
rect 271653 199961 271687 199989
rect 271715 199961 271749 199989
rect 271777 199961 271811 199989
rect 271839 199961 280625 199989
rect 280653 199961 280687 199989
rect 280715 199961 280749 199989
rect 280777 199961 280811 199989
rect 280839 199961 289625 199989
rect 289653 199961 289687 199989
rect 289715 199961 289749 199989
rect 289777 199961 289811 199989
rect 289839 199961 298248 199989
rect 298276 199961 298310 199989
rect 298338 199961 298372 199989
rect 298400 199961 298434 199989
rect 298462 199961 298990 199989
rect -958 199913 298990 199961
rect -958 194175 298990 194223
rect -958 194147 -910 194175
rect -882 194147 -848 194175
rect -820 194147 -786 194175
rect -758 194147 -724 194175
rect -696 194147 3485 194175
rect 3513 194147 3547 194175
rect 3575 194147 3609 194175
rect 3637 194147 3671 194175
rect 3699 194147 12485 194175
rect 12513 194147 12547 194175
rect 12575 194147 12609 194175
rect 12637 194147 12671 194175
rect 12699 194147 21485 194175
rect 21513 194147 21547 194175
rect 21575 194147 21609 194175
rect 21637 194147 21671 194175
rect 21699 194147 30485 194175
rect 30513 194147 30547 194175
rect 30575 194147 30609 194175
rect 30637 194147 30671 194175
rect 30699 194147 39485 194175
rect 39513 194147 39547 194175
rect 39575 194147 39609 194175
rect 39637 194147 39671 194175
rect 39699 194147 48485 194175
rect 48513 194147 48547 194175
rect 48575 194147 48609 194175
rect 48637 194147 48671 194175
rect 48699 194147 57485 194175
rect 57513 194147 57547 194175
rect 57575 194147 57609 194175
rect 57637 194147 57671 194175
rect 57699 194147 66485 194175
rect 66513 194147 66547 194175
rect 66575 194147 66609 194175
rect 66637 194147 66671 194175
rect 66699 194147 75485 194175
rect 75513 194147 75547 194175
rect 75575 194147 75609 194175
rect 75637 194147 75671 194175
rect 75699 194147 84485 194175
rect 84513 194147 84547 194175
rect 84575 194147 84609 194175
rect 84637 194147 84671 194175
rect 84699 194147 93485 194175
rect 93513 194147 93547 194175
rect 93575 194147 93609 194175
rect 93637 194147 93671 194175
rect 93699 194147 102485 194175
rect 102513 194147 102547 194175
rect 102575 194147 102609 194175
rect 102637 194147 102671 194175
rect 102699 194147 111485 194175
rect 111513 194147 111547 194175
rect 111575 194147 111609 194175
rect 111637 194147 111671 194175
rect 111699 194147 120485 194175
rect 120513 194147 120547 194175
rect 120575 194147 120609 194175
rect 120637 194147 120671 194175
rect 120699 194147 129485 194175
rect 129513 194147 129547 194175
rect 129575 194147 129609 194175
rect 129637 194147 129671 194175
rect 129699 194147 138485 194175
rect 138513 194147 138547 194175
rect 138575 194147 138609 194175
rect 138637 194147 138671 194175
rect 138699 194147 147485 194175
rect 147513 194147 147547 194175
rect 147575 194147 147609 194175
rect 147637 194147 147671 194175
rect 147699 194147 156485 194175
rect 156513 194147 156547 194175
rect 156575 194147 156609 194175
rect 156637 194147 156671 194175
rect 156699 194147 165485 194175
rect 165513 194147 165547 194175
rect 165575 194147 165609 194175
rect 165637 194147 165671 194175
rect 165699 194147 174485 194175
rect 174513 194147 174547 194175
rect 174575 194147 174609 194175
rect 174637 194147 174671 194175
rect 174699 194147 183485 194175
rect 183513 194147 183547 194175
rect 183575 194147 183609 194175
rect 183637 194147 183671 194175
rect 183699 194147 192485 194175
rect 192513 194147 192547 194175
rect 192575 194147 192609 194175
rect 192637 194147 192671 194175
rect 192699 194147 201485 194175
rect 201513 194147 201547 194175
rect 201575 194147 201609 194175
rect 201637 194147 201671 194175
rect 201699 194147 210485 194175
rect 210513 194147 210547 194175
rect 210575 194147 210609 194175
rect 210637 194147 210671 194175
rect 210699 194147 219485 194175
rect 219513 194147 219547 194175
rect 219575 194147 219609 194175
rect 219637 194147 219671 194175
rect 219699 194147 228485 194175
rect 228513 194147 228547 194175
rect 228575 194147 228609 194175
rect 228637 194147 228671 194175
rect 228699 194147 237485 194175
rect 237513 194147 237547 194175
rect 237575 194147 237609 194175
rect 237637 194147 237671 194175
rect 237699 194147 246485 194175
rect 246513 194147 246547 194175
rect 246575 194147 246609 194175
rect 246637 194147 246671 194175
rect 246699 194147 255485 194175
rect 255513 194147 255547 194175
rect 255575 194147 255609 194175
rect 255637 194147 255671 194175
rect 255699 194147 264485 194175
rect 264513 194147 264547 194175
rect 264575 194147 264609 194175
rect 264637 194147 264671 194175
rect 264699 194147 273485 194175
rect 273513 194147 273547 194175
rect 273575 194147 273609 194175
rect 273637 194147 273671 194175
rect 273699 194147 282485 194175
rect 282513 194147 282547 194175
rect 282575 194147 282609 194175
rect 282637 194147 282671 194175
rect 282699 194147 291485 194175
rect 291513 194147 291547 194175
rect 291575 194147 291609 194175
rect 291637 194147 291671 194175
rect 291699 194147 298728 194175
rect 298756 194147 298790 194175
rect 298818 194147 298852 194175
rect 298880 194147 298914 194175
rect 298942 194147 298990 194175
rect -958 194113 298990 194147
rect -958 194085 -910 194113
rect -882 194085 -848 194113
rect -820 194085 -786 194113
rect -758 194085 -724 194113
rect -696 194085 3485 194113
rect 3513 194085 3547 194113
rect 3575 194085 3609 194113
rect 3637 194085 3671 194113
rect 3699 194085 12485 194113
rect 12513 194085 12547 194113
rect 12575 194085 12609 194113
rect 12637 194085 12671 194113
rect 12699 194085 21485 194113
rect 21513 194085 21547 194113
rect 21575 194085 21609 194113
rect 21637 194085 21671 194113
rect 21699 194085 30485 194113
rect 30513 194085 30547 194113
rect 30575 194085 30609 194113
rect 30637 194085 30671 194113
rect 30699 194085 39485 194113
rect 39513 194085 39547 194113
rect 39575 194085 39609 194113
rect 39637 194085 39671 194113
rect 39699 194085 48485 194113
rect 48513 194085 48547 194113
rect 48575 194085 48609 194113
rect 48637 194085 48671 194113
rect 48699 194085 57485 194113
rect 57513 194085 57547 194113
rect 57575 194085 57609 194113
rect 57637 194085 57671 194113
rect 57699 194085 66485 194113
rect 66513 194085 66547 194113
rect 66575 194085 66609 194113
rect 66637 194085 66671 194113
rect 66699 194085 75485 194113
rect 75513 194085 75547 194113
rect 75575 194085 75609 194113
rect 75637 194085 75671 194113
rect 75699 194085 84485 194113
rect 84513 194085 84547 194113
rect 84575 194085 84609 194113
rect 84637 194085 84671 194113
rect 84699 194085 93485 194113
rect 93513 194085 93547 194113
rect 93575 194085 93609 194113
rect 93637 194085 93671 194113
rect 93699 194085 102485 194113
rect 102513 194085 102547 194113
rect 102575 194085 102609 194113
rect 102637 194085 102671 194113
rect 102699 194085 111485 194113
rect 111513 194085 111547 194113
rect 111575 194085 111609 194113
rect 111637 194085 111671 194113
rect 111699 194085 120485 194113
rect 120513 194085 120547 194113
rect 120575 194085 120609 194113
rect 120637 194085 120671 194113
rect 120699 194085 129485 194113
rect 129513 194085 129547 194113
rect 129575 194085 129609 194113
rect 129637 194085 129671 194113
rect 129699 194085 138485 194113
rect 138513 194085 138547 194113
rect 138575 194085 138609 194113
rect 138637 194085 138671 194113
rect 138699 194085 147485 194113
rect 147513 194085 147547 194113
rect 147575 194085 147609 194113
rect 147637 194085 147671 194113
rect 147699 194085 156485 194113
rect 156513 194085 156547 194113
rect 156575 194085 156609 194113
rect 156637 194085 156671 194113
rect 156699 194085 165485 194113
rect 165513 194085 165547 194113
rect 165575 194085 165609 194113
rect 165637 194085 165671 194113
rect 165699 194085 174485 194113
rect 174513 194085 174547 194113
rect 174575 194085 174609 194113
rect 174637 194085 174671 194113
rect 174699 194085 183485 194113
rect 183513 194085 183547 194113
rect 183575 194085 183609 194113
rect 183637 194085 183671 194113
rect 183699 194085 192485 194113
rect 192513 194085 192547 194113
rect 192575 194085 192609 194113
rect 192637 194085 192671 194113
rect 192699 194085 201485 194113
rect 201513 194085 201547 194113
rect 201575 194085 201609 194113
rect 201637 194085 201671 194113
rect 201699 194085 210485 194113
rect 210513 194085 210547 194113
rect 210575 194085 210609 194113
rect 210637 194085 210671 194113
rect 210699 194085 219485 194113
rect 219513 194085 219547 194113
rect 219575 194085 219609 194113
rect 219637 194085 219671 194113
rect 219699 194085 228485 194113
rect 228513 194085 228547 194113
rect 228575 194085 228609 194113
rect 228637 194085 228671 194113
rect 228699 194085 237485 194113
rect 237513 194085 237547 194113
rect 237575 194085 237609 194113
rect 237637 194085 237671 194113
rect 237699 194085 246485 194113
rect 246513 194085 246547 194113
rect 246575 194085 246609 194113
rect 246637 194085 246671 194113
rect 246699 194085 255485 194113
rect 255513 194085 255547 194113
rect 255575 194085 255609 194113
rect 255637 194085 255671 194113
rect 255699 194085 264485 194113
rect 264513 194085 264547 194113
rect 264575 194085 264609 194113
rect 264637 194085 264671 194113
rect 264699 194085 273485 194113
rect 273513 194085 273547 194113
rect 273575 194085 273609 194113
rect 273637 194085 273671 194113
rect 273699 194085 282485 194113
rect 282513 194085 282547 194113
rect 282575 194085 282609 194113
rect 282637 194085 282671 194113
rect 282699 194085 291485 194113
rect 291513 194085 291547 194113
rect 291575 194085 291609 194113
rect 291637 194085 291671 194113
rect 291699 194085 298728 194113
rect 298756 194085 298790 194113
rect 298818 194085 298852 194113
rect 298880 194085 298914 194113
rect 298942 194085 298990 194113
rect -958 194051 298990 194085
rect -958 194023 -910 194051
rect -882 194023 -848 194051
rect -820 194023 -786 194051
rect -758 194023 -724 194051
rect -696 194023 3485 194051
rect 3513 194023 3547 194051
rect 3575 194023 3609 194051
rect 3637 194023 3671 194051
rect 3699 194023 12485 194051
rect 12513 194023 12547 194051
rect 12575 194023 12609 194051
rect 12637 194023 12671 194051
rect 12699 194023 21485 194051
rect 21513 194023 21547 194051
rect 21575 194023 21609 194051
rect 21637 194023 21671 194051
rect 21699 194023 30485 194051
rect 30513 194023 30547 194051
rect 30575 194023 30609 194051
rect 30637 194023 30671 194051
rect 30699 194023 39485 194051
rect 39513 194023 39547 194051
rect 39575 194023 39609 194051
rect 39637 194023 39671 194051
rect 39699 194023 48485 194051
rect 48513 194023 48547 194051
rect 48575 194023 48609 194051
rect 48637 194023 48671 194051
rect 48699 194023 57485 194051
rect 57513 194023 57547 194051
rect 57575 194023 57609 194051
rect 57637 194023 57671 194051
rect 57699 194023 66485 194051
rect 66513 194023 66547 194051
rect 66575 194023 66609 194051
rect 66637 194023 66671 194051
rect 66699 194023 75485 194051
rect 75513 194023 75547 194051
rect 75575 194023 75609 194051
rect 75637 194023 75671 194051
rect 75699 194023 84485 194051
rect 84513 194023 84547 194051
rect 84575 194023 84609 194051
rect 84637 194023 84671 194051
rect 84699 194023 93485 194051
rect 93513 194023 93547 194051
rect 93575 194023 93609 194051
rect 93637 194023 93671 194051
rect 93699 194023 102485 194051
rect 102513 194023 102547 194051
rect 102575 194023 102609 194051
rect 102637 194023 102671 194051
rect 102699 194023 111485 194051
rect 111513 194023 111547 194051
rect 111575 194023 111609 194051
rect 111637 194023 111671 194051
rect 111699 194023 120485 194051
rect 120513 194023 120547 194051
rect 120575 194023 120609 194051
rect 120637 194023 120671 194051
rect 120699 194023 129485 194051
rect 129513 194023 129547 194051
rect 129575 194023 129609 194051
rect 129637 194023 129671 194051
rect 129699 194023 138485 194051
rect 138513 194023 138547 194051
rect 138575 194023 138609 194051
rect 138637 194023 138671 194051
rect 138699 194023 147485 194051
rect 147513 194023 147547 194051
rect 147575 194023 147609 194051
rect 147637 194023 147671 194051
rect 147699 194023 156485 194051
rect 156513 194023 156547 194051
rect 156575 194023 156609 194051
rect 156637 194023 156671 194051
rect 156699 194023 165485 194051
rect 165513 194023 165547 194051
rect 165575 194023 165609 194051
rect 165637 194023 165671 194051
rect 165699 194023 174485 194051
rect 174513 194023 174547 194051
rect 174575 194023 174609 194051
rect 174637 194023 174671 194051
rect 174699 194023 183485 194051
rect 183513 194023 183547 194051
rect 183575 194023 183609 194051
rect 183637 194023 183671 194051
rect 183699 194023 192485 194051
rect 192513 194023 192547 194051
rect 192575 194023 192609 194051
rect 192637 194023 192671 194051
rect 192699 194023 201485 194051
rect 201513 194023 201547 194051
rect 201575 194023 201609 194051
rect 201637 194023 201671 194051
rect 201699 194023 210485 194051
rect 210513 194023 210547 194051
rect 210575 194023 210609 194051
rect 210637 194023 210671 194051
rect 210699 194023 219485 194051
rect 219513 194023 219547 194051
rect 219575 194023 219609 194051
rect 219637 194023 219671 194051
rect 219699 194023 228485 194051
rect 228513 194023 228547 194051
rect 228575 194023 228609 194051
rect 228637 194023 228671 194051
rect 228699 194023 237485 194051
rect 237513 194023 237547 194051
rect 237575 194023 237609 194051
rect 237637 194023 237671 194051
rect 237699 194023 246485 194051
rect 246513 194023 246547 194051
rect 246575 194023 246609 194051
rect 246637 194023 246671 194051
rect 246699 194023 255485 194051
rect 255513 194023 255547 194051
rect 255575 194023 255609 194051
rect 255637 194023 255671 194051
rect 255699 194023 264485 194051
rect 264513 194023 264547 194051
rect 264575 194023 264609 194051
rect 264637 194023 264671 194051
rect 264699 194023 273485 194051
rect 273513 194023 273547 194051
rect 273575 194023 273609 194051
rect 273637 194023 273671 194051
rect 273699 194023 282485 194051
rect 282513 194023 282547 194051
rect 282575 194023 282609 194051
rect 282637 194023 282671 194051
rect 282699 194023 291485 194051
rect 291513 194023 291547 194051
rect 291575 194023 291609 194051
rect 291637 194023 291671 194051
rect 291699 194023 298728 194051
rect 298756 194023 298790 194051
rect 298818 194023 298852 194051
rect 298880 194023 298914 194051
rect 298942 194023 298990 194051
rect -958 193989 298990 194023
rect -958 193961 -910 193989
rect -882 193961 -848 193989
rect -820 193961 -786 193989
rect -758 193961 -724 193989
rect -696 193961 3485 193989
rect 3513 193961 3547 193989
rect 3575 193961 3609 193989
rect 3637 193961 3671 193989
rect 3699 193961 12485 193989
rect 12513 193961 12547 193989
rect 12575 193961 12609 193989
rect 12637 193961 12671 193989
rect 12699 193961 21485 193989
rect 21513 193961 21547 193989
rect 21575 193961 21609 193989
rect 21637 193961 21671 193989
rect 21699 193961 30485 193989
rect 30513 193961 30547 193989
rect 30575 193961 30609 193989
rect 30637 193961 30671 193989
rect 30699 193961 39485 193989
rect 39513 193961 39547 193989
rect 39575 193961 39609 193989
rect 39637 193961 39671 193989
rect 39699 193961 48485 193989
rect 48513 193961 48547 193989
rect 48575 193961 48609 193989
rect 48637 193961 48671 193989
rect 48699 193961 57485 193989
rect 57513 193961 57547 193989
rect 57575 193961 57609 193989
rect 57637 193961 57671 193989
rect 57699 193961 66485 193989
rect 66513 193961 66547 193989
rect 66575 193961 66609 193989
rect 66637 193961 66671 193989
rect 66699 193961 75485 193989
rect 75513 193961 75547 193989
rect 75575 193961 75609 193989
rect 75637 193961 75671 193989
rect 75699 193961 84485 193989
rect 84513 193961 84547 193989
rect 84575 193961 84609 193989
rect 84637 193961 84671 193989
rect 84699 193961 93485 193989
rect 93513 193961 93547 193989
rect 93575 193961 93609 193989
rect 93637 193961 93671 193989
rect 93699 193961 102485 193989
rect 102513 193961 102547 193989
rect 102575 193961 102609 193989
rect 102637 193961 102671 193989
rect 102699 193961 111485 193989
rect 111513 193961 111547 193989
rect 111575 193961 111609 193989
rect 111637 193961 111671 193989
rect 111699 193961 120485 193989
rect 120513 193961 120547 193989
rect 120575 193961 120609 193989
rect 120637 193961 120671 193989
rect 120699 193961 129485 193989
rect 129513 193961 129547 193989
rect 129575 193961 129609 193989
rect 129637 193961 129671 193989
rect 129699 193961 138485 193989
rect 138513 193961 138547 193989
rect 138575 193961 138609 193989
rect 138637 193961 138671 193989
rect 138699 193961 147485 193989
rect 147513 193961 147547 193989
rect 147575 193961 147609 193989
rect 147637 193961 147671 193989
rect 147699 193961 156485 193989
rect 156513 193961 156547 193989
rect 156575 193961 156609 193989
rect 156637 193961 156671 193989
rect 156699 193961 165485 193989
rect 165513 193961 165547 193989
rect 165575 193961 165609 193989
rect 165637 193961 165671 193989
rect 165699 193961 174485 193989
rect 174513 193961 174547 193989
rect 174575 193961 174609 193989
rect 174637 193961 174671 193989
rect 174699 193961 183485 193989
rect 183513 193961 183547 193989
rect 183575 193961 183609 193989
rect 183637 193961 183671 193989
rect 183699 193961 192485 193989
rect 192513 193961 192547 193989
rect 192575 193961 192609 193989
rect 192637 193961 192671 193989
rect 192699 193961 201485 193989
rect 201513 193961 201547 193989
rect 201575 193961 201609 193989
rect 201637 193961 201671 193989
rect 201699 193961 210485 193989
rect 210513 193961 210547 193989
rect 210575 193961 210609 193989
rect 210637 193961 210671 193989
rect 210699 193961 219485 193989
rect 219513 193961 219547 193989
rect 219575 193961 219609 193989
rect 219637 193961 219671 193989
rect 219699 193961 228485 193989
rect 228513 193961 228547 193989
rect 228575 193961 228609 193989
rect 228637 193961 228671 193989
rect 228699 193961 237485 193989
rect 237513 193961 237547 193989
rect 237575 193961 237609 193989
rect 237637 193961 237671 193989
rect 237699 193961 246485 193989
rect 246513 193961 246547 193989
rect 246575 193961 246609 193989
rect 246637 193961 246671 193989
rect 246699 193961 255485 193989
rect 255513 193961 255547 193989
rect 255575 193961 255609 193989
rect 255637 193961 255671 193989
rect 255699 193961 264485 193989
rect 264513 193961 264547 193989
rect 264575 193961 264609 193989
rect 264637 193961 264671 193989
rect 264699 193961 273485 193989
rect 273513 193961 273547 193989
rect 273575 193961 273609 193989
rect 273637 193961 273671 193989
rect 273699 193961 282485 193989
rect 282513 193961 282547 193989
rect 282575 193961 282609 193989
rect 282637 193961 282671 193989
rect 282699 193961 291485 193989
rect 291513 193961 291547 193989
rect 291575 193961 291609 193989
rect 291637 193961 291671 193989
rect 291699 193961 298728 193989
rect 298756 193961 298790 193989
rect 298818 193961 298852 193989
rect 298880 193961 298914 193989
rect 298942 193961 298990 193989
rect -958 193913 298990 193961
rect -958 191175 298990 191223
rect -958 191147 -430 191175
rect -402 191147 -368 191175
rect -340 191147 -306 191175
rect -278 191147 -244 191175
rect -216 191147 1625 191175
rect 1653 191147 1687 191175
rect 1715 191147 1749 191175
rect 1777 191147 1811 191175
rect 1839 191147 10625 191175
rect 10653 191147 10687 191175
rect 10715 191147 10749 191175
rect 10777 191147 10811 191175
rect 10839 191147 19625 191175
rect 19653 191147 19687 191175
rect 19715 191147 19749 191175
rect 19777 191147 19811 191175
rect 19839 191147 28625 191175
rect 28653 191147 28687 191175
rect 28715 191147 28749 191175
rect 28777 191147 28811 191175
rect 28839 191147 37625 191175
rect 37653 191147 37687 191175
rect 37715 191147 37749 191175
rect 37777 191147 37811 191175
rect 37839 191147 46625 191175
rect 46653 191147 46687 191175
rect 46715 191147 46749 191175
rect 46777 191147 46811 191175
rect 46839 191147 154625 191175
rect 154653 191147 154687 191175
rect 154715 191147 154749 191175
rect 154777 191147 154811 191175
rect 154839 191147 163625 191175
rect 163653 191147 163687 191175
rect 163715 191147 163749 191175
rect 163777 191147 163811 191175
rect 163839 191147 172625 191175
rect 172653 191147 172687 191175
rect 172715 191147 172749 191175
rect 172777 191147 172811 191175
rect 172839 191147 181625 191175
rect 181653 191147 181687 191175
rect 181715 191147 181749 191175
rect 181777 191147 181811 191175
rect 181839 191147 190625 191175
rect 190653 191147 190687 191175
rect 190715 191147 190749 191175
rect 190777 191147 190811 191175
rect 190839 191147 199625 191175
rect 199653 191147 199687 191175
rect 199715 191147 199749 191175
rect 199777 191147 199811 191175
rect 199839 191147 208625 191175
rect 208653 191147 208687 191175
rect 208715 191147 208749 191175
rect 208777 191147 208811 191175
rect 208839 191147 217625 191175
rect 217653 191147 217687 191175
rect 217715 191147 217749 191175
rect 217777 191147 217811 191175
rect 217839 191147 226625 191175
rect 226653 191147 226687 191175
rect 226715 191147 226749 191175
rect 226777 191147 226811 191175
rect 226839 191147 235625 191175
rect 235653 191147 235687 191175
rect 235715 191147 235749 191175
rect 235777 191147 235811 191175
rect 235839 191147 244625 191175
rect 244653 191147 244687 191175
rect 244715 191147 244749 191175
rect 244777 191147 244811 191175
rect 244839 191147 253625 191175
rect 253653 191147 253687 191175
rect 253715 191147 253749 191175
rect 253777 191147 253811 191175
rect 253839 191147 262625 191175
rect 262653 191147 262687 191175
rect 262715 191147 262749 191175
rect 262777 191147 262811 191175
rect 262839 191147 271625 191175
rect 271653 191147 271687 191175
rect 271715 191147 271749 191175
rect 271777 191147 271811 191175
rect 271839 191147 280625 191175
rect 280653 191147 280687 191175
rect 280715 191147 280749 191175
rect 280777 191147 280811 191175
rect 280839 191147 289625 191175
rect 289653 191147 289687 191175
rect 289715 191147 289749 191175
rect 289777 191147 289811 191175
rect 289839 191147 298248 191175
rect 298276 191147 298310 191175
rect 298338 191147 298372 191175
rect 298400 191147 298434 191175
rect 298462 191147 298990 191175
rect -958 191113 298990 191147
rect -958 191085 -430 191113
rect -402 191085 -368 191113
rect -340 191085 -306 191113
rect -278 191085 -244 191113
rect -216 191085 1625 191113
rect 1653 191085 1687 191113
rect 1715 191085 1749 191113
rect 1777 191085 1811 191113
rect 1839 191085 10625 191113
rect 10653 191085 10687 191113
rect 10715 191085 10749 191113
rect 10777 191085 10811 191113
rect 10839 191085 19625 191113
rect 19653 191085 19687 191113
rect 19715 191085 19749 191113
rect 19777 191085 19811 191113
rect 19839 191085 28625 191113
rect 28653 191085 28687 191113
rect 28715 191085 28749 191113
rect 28777 191085 28811 191113
rect 28839 191085 37625 191113
rect 37653 191085 37687 191113
rect 37715 191085 37749 191113
rect 37777 191085 37811 191113
rect 37839 191085 46625 191113
rect 46653 191085 46687 191113
rect 46715 191085 46749 191113
rect 46777 191085 46811 191113
rect 46839 191085 154625 191113
rect 154653 191085 154687 191113
rect 154715 191085 154749 191113
rect 154777 191085 154811 191113
rect 154839 191085 163625 191113
rect 163653 191085 163687 191113
rect 163715 191085 163749 191113
rect 163777 191085 163811 191113
rect 163839 191085 172625 191113
rect 172653 191085 172687 191113
rect 172715 191085 172749 191113
rect 172777 191085 172811 191113
rect 172839 191085 181625 191113
rect 181653 191085 181687 191113
rect 181715 191085 181749 191113
rect 181777 191085 181811 191113
rect 181839 191085 190625 191113
rect 190653 191085 190687 191113
rect 190715 191085 190749 191113
rect 190777 191085 190811 191113
rect 190839 191085 199625 191113
rect 199653 191085 199687 191113
rect 199715 191085 199749 191113
rect 199777 191085 199811 191113
rect 199839 191085 208625 191113
rect 208653 191085 208687 191113
rect 208715 191085 208749 191113
rect 208777 191085 208811 191113
rect 208839 191085 217625 191113
rect 217653 191085 217687 191113
rect 217715 191085 217749 191113
rect 217777 191085 217811 191113
rect 217839 191085 226625 191113
rect 226653 191085 226687 191113
rect 226715 191085 226749 191113
rect 226777 191085 226811 191113
rect 226839 191085 235625 191113
rect 235653 191085 235687 191113
rect 235715 191085 235749 191113
rect 235777 191085 235811 191113
rect 235839 191085 244625 191113
rect 244653 191085 244687 191113
rect 244715 191085 244749 191113
rect 244777 191085 244811 191113
rect 244839 191085 253625 191113
rect 253653 191085 253687 191113
rect 253715 191085 253749 191113
rect 253777 191085 253811 191113
rect 253839 191085 262625 191113
rect 262653 191085 262687 191113
rect 262715 191085 262749 191113
rect 262777 191085 262811 191113
rect 262839 191085 271625 191113
rect 271653 191085 271687 191113
rect 271715 191085 271749 191113
rect 271777 191085 271811 191113
rect 271839 191085 280625 191113
rect 280653 191085 280687 191113
rect 280715 191085 280749 191113
rect 280777 191085 280811 191113
rect 280839 191085 289625 191113
rect 289653 191085 289687 191113
rect 289715 191085 289749 191113
rect 289777 191085 289811 191113
rect 289839 191085 298248 191113
rect 298276 191085 298310 191113
rect 298338 191085 298372 191113
rect 298400 191085 298434 191113
rect 298462 191085 298990 191113
rect -958 191051 298990 191085
rect -958 191023 -430 191051
rect -402 191023 -368 191051
rect -340 191023 -306 191051
rect -278 191023 -244 191051
rect -216 191023 1625 191051
rect 1653 191023 1687 191051
rect 1715 191023 1749 191051
rect 1777 191023 1811 191051
rect 1839 191023 10625 191051
rect 10653 191023 10687 191051
rect 10715 191023 10749 191051
rect 10777 191023 10811 191051
rect 10839 191023 19625 191051
rect 19653 191023 19687 191051
rect 19715 191023 19749 191051
rect 19777 191023 19811 191051
rect 19839 191023 28625 191051
rect 28653 191023 28687 191051
rect 28715 191023 28749 191051
rect 28777 191023 28811 191051
rect 28839 191023 37625 191051
rect 37653 191023 37687 191051
rect 37715 191023 37749 191051
rect 37777 191023 37811 191051
rect 37839 191023 46625 191051
rect 46653 191023 46687 191051
rect 46715 191023 46749 191051
rect 46777 191023 46811 191051
rect 46839 191023 154625 191051
rect 154653 191023 154687 191051
rect 154715 191023 154749 191051
rect 154777 191023 154811 191051
rect 154839 191023 163625 191051
rect 163653 191023 163687 191051
rect 163715 191023 163749 191051
rect 163777 191023 163811 191051
rect 163839 191023 172625 191051
rect 172653 191023 172687 191051
rect 172715 191023 172749 191051
rect 172777 191023 172811 191051
rect 172839 191023 181625 191051
rect 181653 191023 181687 191051
rect 181715 191023 181749 191051
rect 181777 191023 181811 191051
rect 181839 191023 190625 191051
rect 190653 191023 190687 191051
rect 190715 191023 190749 191051
rect 190777 191023 190811 191051
rect 190839 191023 199625 191051
rect 199653 191023 199687 191051
rect 199715 191023 199749 191051
rect 199777 191023 199811 191051
rect 199839 191023 208625 191051
rect 208653 191023 208687 191051
rect 208715 191023 208749 191051
rect 208777 191023 208811 191051
rect 208839 191023 217625 191051
rect 217653 191023 217687 191051
rect 217715 191023 217749 191051
rect 217777 191023 217811 191051
rect 217839 191023 226625 191051
rect 226653 191023 226687 191051
rect 226715 191023 226749 191051
rect 226777 191023 226811 191051
rect 226839 191023 235625 191051
rect 235653 191023 235687 191051
rect 235715 191023 235749 191051
rect 235777 191023 235811 191051
rect 235839 191023 244625 191051
rect 244653 191023 244687 191051
rect 244715 191023 244749 191051
rect 244777 191023 244811 191051
rect 244839 191023 253625 191051
rect 253653 191023 253687 191051
rect 253715 191023 253749 191051
rect 253777 191023 253811 191051
rect 253839 191023 262625 191051
rect 262653 191023 262687 191051
rect 262715 191023 262749 191051
rect 262777 191023 262811 191051
rect 262839 191023 271625 191051
rect 271653 191023 271687 191051
rect 271715 191023 271749 191051
rect 271777 191023 271811 191051
rect 271839 191023 280625 191051
rect 280653 191023 280687 191051
rect 280715 191023 280749 191051
rect 280777 191023 280811 191051
rect 280839 191023 289625 191051
rect 289653 191023 289687 191051
rect 289715 191023 289749 191051
rect 289777 191023 289811 191051
rect 289839 191023 298248 191051
rect 298276 191023 298310 191051
rect 298338 191023 298372 191051
rect 298400 191023 298434 191051
rect 298462 191023 298990 191051
rect -958 190989 298990 191023
rect -958 190961 -430 190989
rect -402 190961 -368 190989
rect -340 190961 -306 190989
rect -278 190961 -244 190989
rect -216 190961 1625 190989
rect 1653 190961 1687 190989
rect 1715 190961 1749 190989
rect 1777 190961 1811 190989
rect 1839 190961 10625 190989
rect 10653 190961 10687 190989
rect 10715 190961 10749 190989
rect 10777 190961 10811 190989
rect 10839 190961 19625 190989
rect 19653 190961 19687 190989
rect 19715 190961 19749 190989
rect 19777 190961 19811 190989
rect 19839 190961 28625 190989
rect 28653 190961 28687 190989
rect 28715 190961 28749 190989
rect 28777 190961 28811 190989
rect 28839 190961 37625 190989
rect 37653 190961 37687 190989
rect 37715 190961 37749 190989
rect 37777 190961 37811 190989
rect 37839 190961 46625 190989
rect 46653 190961 46687 190989
rect 46715 190961 46749 190989
rect 46777 190961 46811 190989
rect 46839 190961 154625 190989
rect 154653 190961 154687 190989
rect 154715 190961 154749 190989
rect 154777 190961 154811 190989
rect 154839 190961 163625 190989
rect 163653 190961 163687 190989
rect 163715 190961 163749 190989
rect 163777 190961 163811 190989
rect 163839 190961 172625 190989
rect 172653 190961 172687 190989
rect 172715 190961 172749 190989
rect 172777 190961 172811 190989
rect 172839 190961 181625 190989
rect 181653 190961 181687 190989
rect 181715 190961 181749 190989
rect 181777 190961 181811 190989
rect 181839 190961 190625 190989
rect 190653 190961 190687 190989
rect 190715 190961 190749 190989
rect 190777 190961 190811 190989
rect 190839 190961 199625 190989
rect 199653 190961 199687 190989
rect 199715 190961 199749 190989
rect 199777 190961 199811 190989
rect 199839 190961 208625 190989
rect 208653 190961 208687 190989
rect 208715 190961 208749 190989
rect 208777 190961 208811 190989
rect 208839 190961 217625 190989
rect 217653 190961 217687 190989
rect 217715 190961 217749 190989
rect 217777 190961 217811 190989
rect 217839 190961 226625 190989
rect 226653 190961 226687 190989
rect 226715 190961 226749 190989
rect 226777 190961 226811 190989
rect 226839 190961 235625 190989
rect 235653 190961 235687 190989
rect 235715 190961 235749 190989
rect 235777 190961 235811 190989
rect 235839 190961 244625 190989
rect 244653 190961 244687 190989
rect 244715 190961 244749 190989
rect 244777 190961 244811 190989
rect 244839 190961 253625 190989
rect 253653 190961 253687 190989
rect 253715 190961 253749 190989
rect 253777 190961 253811 190989
rect 253839 190961 262625 190989
rect 262653 190961 262687 190989
rect 262715 190961 262749 190989
rect 262777 190961 262811 190989
rect 262839 190961 271625 190989
rect 271653 190961 271687 190989
rect 271715 190961 271749 190989
rect 271777 190961 271811 190989
rect 271839 190961 280625 190989
rect 280653 190961 280687 190989
rect 280715 190961 280749 190989
rect 280777 190961 280811 190989
rect 280839 190961 289625 190989
rect 289653 190961 289687 190989
rect 289715 190961 289749 190989
rect 289777 190961 289811 190989
rect 289839 190961 298248 190989
rect 298276 190961 298310 190989
rect 298338 190961 298372 190989
rect 298400 190961 298434 190989
rect 298462 190961 298990 190989
rect -958 190913 298990 190961
rect -958 185175 298990 185223
rect -958 185147 -910 185175
rect -882 185147 -848 185175
rect -820 185147 -786 185175
rect -758 185147 -724 185175
rect -696 185147 3485 185175
rect 3513 185147 3547 185175
rect 3575 185147 3609 185175
rect 3637 185147 3671 185175
rect 3699 185147 12485 185175
rect 12513 185147 12547 185175
rect 12575 185147 12609 185175
rect 12637 185147 12671 185175
rect 12699 185147 21485 185175
rect 21513 185147 21547 185175
rect 21575 185147 21609 185175
rect 21637 185147 21671 185175
rect 21699 185147 30485 185175
rect 30513 185147 30547 185175
rect 30575 185147 30609 185175
rect 30637 185147 30671 185175
rect 30699 185147 39485 185175
rect 39513 185147 39547 185175
rect 39575 185147 39609 185175
rect 39637 185147 39671 185175
rect 39699 185147 48485 185175
rect 48513 185147 48547 185175
rect 48575 185147 48609 185175
rect 48637 185147 48671 185175
rect 48699 185147 57485 185175
rect 57513 185147 57547 185175
rect 57575 185147 57609 185175
rect 57637 185147 57671 185175
rect 57699 185147 66485 185175
rect 66513 185147 66547 185175
rect 66575 185147 66609 185175
rect 66637 185147 66671 185175
rect 66699 185147 75485 185175
rect 75513 185147 75547 185175
rect 75575 185147 75609 185175
rect 75637 185147 75671 185175
rect 75699 185147 84485 185175
rect 84513 185147 84547 185175
rect 84575 185147 84609 185175
rect 84637 185147 84671 185175
rect 84699 185147 93485 185175
rect 93513 185147 93547 185175
rect 93575 185147 93609 185175
rect 93637 185147 93671 185175
rect 93699 185147 102485 185175
rect 102513 185147 102547 185175
rect 102575 185147 102609 185175
rect 102637 185147 102671 185175
rect 102699 185147 111485 185175
rect 111513 185147 111547 185175
rect 111575 185147 111609 185175
rect 111637 185147 111671 185175
rect 111699 185147 120485 185175
rect 120513 185147 120547 185175
rect 120575 185147 120609 185175
rect 120637 185147 120671 185175
rect 120699 185147 129485 185175
rect 129513 185147 129547 185175
rect 129575 185147 129609 185175
rect 129637 185147 129671 185175
rect 129699 185147 138485 185175
rect 138513 185147 138547 185175
rect 138575 185147 138609 185175
rect 138637 185147 138671 185175
rect 138699 185147 147485 185175
rect 147513 185147 147547 185175
rect 147575 185147 147609 185175
rect 147637 185147 147671 185175
rect 147699 185147 156485 185175
rect 156513 185147 156547 185175
rect 156575 185147 156609 185175
rect 156637 185147 156671 185175
rect 156699 185147 165485 185175
rect 165513 185147 165547 185175
rect 165575 185147 165609 185175
rect 165637 185147 165671 185175
rect 165699 185147 174485 185175
rect 174513 185147 174547 185175
rect 174575 185147 174609 185175
rect 174637 185147 174671 185175
rect 174699 185147 183485 185175
rect 183513 185147 183547 185175
rect 183575 185147 183609 185175
rect 183637 185147 183671 185175
rect 183699 185147 192485 185175
rect 192513 185147 192547 185175
rect 192575 185147 192609 185175
rect 192637 185147 192671 185175
rect 192699 185147 201485 185175
rect 201513 185147 201547 185175
rect 201575 185147 201609 185175
rect 201637 185147 201671 185175
rect 201699 185147 210485 185175
rect 210513 185147 210547 185175
rect 210575 185147 210609 185175
rect 210637 185147 210671 185175
rect 210699 185147 219485 185175
rect 219513 185147 219547 185175
rect 219575 185147 219609 185175
rect 219637 185147 219671 185175
rect 219699 185147 228485 185175
rect 228513 185147 228547 185175
rect 228575 185147 228609 185175
rect 228637 185147 228671 185175
rect 228699 185147 237485 185175
rect 237513 185147 237547 185175
rect 237575 185147 237609 185175
rect 237637 185147 237671 185175
rect 237699 185147 246485 185175
rect 246513 185147 246547 185175
rect 246575 185147 246609 185175
rect 246637 185147 246671 185175
rect 246699 185147 255485 185175
rect 255513 185147 255547 185175
rect 255575 185147 255609 185175
rect 255637 185147 255671 185175
rect 255699 185147 264485 185175
rect 264513 185147 264547 185175
rect 264575 185147 264609 185175
rect 264637 185147 264671 185175
rect 264699 185147 273485 185175
rect 273513 185147 273547 185175
rect 273575 185147 273609 185175
rect 273637 185147 273671 185175
rect 273699 185147 282485 185175
rect 282513 185147 282547 185175
rect 282575 185147 282609 185175
rect 282637 185147 282671 185175
rect 282699 185147 291485 185175
rect 291513 185147 291547 185175
rect 291575 185147 291609 185175
rect 291637 185147 291671 185175
rect 291699 185147 298728 185175
rect 298756 185147 298790 185175
rect 298818 185147 298852 185175
rect 298880 185147 298914 185175
rect 298942 185147 298990 185175
rect -958 185113 298990 185147
rect -958 185085 -910 185113
rect -882 185085 -848 185113
rect -820 185085 -786 185113
rect -758 185085 -724 185113
rect -696 185085 3485 185113
rect 3513 185085 3547 185113
rect 3575 185085 3609 185113
rect 3637 185085 3671 185113
rect 3699 185085 12485 185113
rect 12513 185085 12547 185113
rect 12575 185085 12609 185113
rect 12637 185085 12671 185113
rect 12699 185085 21485 185113
rect 21513 185085 21547 185113
rect 21575 185085 21609 185113
rect 21637 185085 21671 185113
rect 21699 185085 30485 185113
rect 30513 185085 30547 185113
rect 30575 185085 30609 185113
rect 30637 185085 30671 185113
rect 30699 185085 39485 185113
rect 39513 185085 39547 185113
rect 39575 185085 39609 185113
rect 39637 185085 39671 185113
rect 39699 185085 48485 185113
rect 48513 185085 48547 185113
rect 48575 185085 48609 185113
rect 48637 185085 48671 185113
rect 48699 185085 57485 185113
rect 57513 185085 57547 185113
rect 57575 185085 57609 185113
rect 57637 185085 57671 185113
rect 57699 185085 66485 185113
rect 66513 185085 66547 185113
rect 66575 185085 66609 185113
rect 66637 185085 66671 185113
rect 66699 185085 75485 185113
rect 75513 185085 75547 185113
rect 75575 185085 75609 185113
rect 75637 185085 75671 185113
rect 75699 185085 84485 185113
rect 84513 185085 84547 185113
rect 84575 185085 84609 185113
rect 84637 185085 84671 185113
rect 84699 185085 93485 185113
rect 93513 185085 93547 185113
rect 93575 185085 93609 185113
rect 93637 185085 93671 185113
rect 93699 185085 102485 185113
rect 102513 185085 102547 185113
rect 102575 185085 102609 185113
rect 102637 185085 102671 185113
rect 102699 185085 111485 185113
rect 111513 185085 111547 185113
rect 111575 185085 111609 185113
rect 111637 185085 111671 185113
rect 111699 185085 120485 185113
rect 120513 185085 120547 185113
rect 120575 185085 120609 185113
rect 120637 185085 120671 185113
rect 120699 185085 129485 185113
rect 129513 185085 129547 185113
rect 129575 185085 129609 185113
rect 129637 185085 129671 185113
rect 129699 185085 138485 185113
rect 138513 185085 138547 185113
rect 138575 185085 138609 185113
rect 138637 185085 138671 185113
rect 138699 185085 147485 185113
rect 147513 185085 147547 185113
rect 147575 185085 147609 185113
rect 147637 185085 147671 185113
rect 147699 185085 156485 185113
rect 156513 185085 156547 185113
rect 156575 185085 156609 185113
rect 156637 185085 156671 185113
rect 156699 185085 165485 185113
rect 165513 185085 165547 185113
rect 165575 185085 165609 185113
rect 165637 185085 165671 185113
rect 165699 185085 174485 185113
rect 174513 185085 174547 185113
rect 174575 185085 174609 185113
rect 174637 185085 174671 185113
rect 174699 185085 183485 185113
rect 183513 185085 183547 185113
rect 183575 185085 183609 185113
rect 183637 185085 183671 185113
rect 183699 185085 192485 185113
rect 192513 185085 192547 185113
rect 192575 185085 192609 185113
rect 192637 185085 192671 185113
rect 192699 185085 201485 185113
rect 201513 185085 201547 185113
rect 201575 185085 201609 185113
rect 201637 185085 201671 185113
rect 201699 185085 210485 185113
rect 210513 185085 210547 185113
rect 210575 185085 210609 185113
rect 210637 185085 210671 185113
rect 210699 185085 219485 185113
rect 219513 185085 219547 185113
rect 219575 185085 219609 185113
rect 219637 185085 219671 185113
rect 219699 185085 228485 185113
rect 228513 185085 228547 185113
rect 228575 185085 228609 185113
rect 228637 185085 228671 185113
rect 228699 185085 237485 185113
rect 237513 185085 237547 185113
rect 237575 185085 237609 185113
rect 237637 185085 237671 185113
rect 237699 185085 246485 185113
rect 246513 185085 246547 185113
rect 246575 185085 246609 185113
rect 246637 185085 246671 185113
rect 246699 185085 255485 185113
rect 255513 185085 255547 185113
rect 255575 185085 255609 185113
rect 255637 185085 255671 185113
rect 255699 185085 264485 185113
rect 264513 185085 264547 185113
rect 264575 185085 264609 185113
rect 264637 185085 264671 185113
rect 264699 185085 273485 185113
rect 273513 185085 273547 185113
rect 273575 185085 273609 185113
rect 273637 185085 273671 185113
rect 273699 185085 282485 185113
rect 282513 185085 282547 185113
rect 282575 185085 282609 185113
rect 282637 185085 282671 185113
rect 282699 185085 291485 185113
rect 291513 185085 291547 185113
rect 291575 185085 291609 185113
rect 291637 185085 291671 185113
rect 291699 185085 298728 185113
rect 298756 185085 298790 185113
rect 298818 185085 298852 185113
rect 298880 185085 298914 185113
rect 298942 185085 298990 185113
rect -958 185051 298990 185085
rect -958 185023 -910 185051
rect -882 185023 -848 185051
rect -820 185023 -786 185051
rect -758 185023 -724 185051
rect -696 185023 3485 185051
rect 3513 185023 3547 185051
rect 3575 185023 3609 185051
rect 3637 185023 3671 185051
rect 3699 185023 12485 185051
rect 12513 185023 12547 185051
rect 12575 185023 12609 185051
rect 12637 185023 12671 185051
rect 12699 185023 21485 185051
rect 21513 185023 21547 185051
rect 21575 185023 21609 185051
rect 21637 185023 21671 185051
rect 21699 185023 30485 185051
rect 30513 185023 30547 185051
rect 30575 185023 30609 185051
rect 30637 185023 30671 185051
rect 30699 185023 39485 185051
rect 39513 185023 39547 185051
rect 39575 185023 39609 185051
rect 39637 185023 39671 185051
rect 39699 185023 48485 185051
rect 48513 185023 48547 185051
rect 48575 185023 48609 185051
rect 48637 185023 48671 185051
rect 48699 185023 57485 185051
rect 57513 185023 57547 185051
rect 57575 185023 57609 185051
rect 57637 185023 57671 185051
rect 57699 185023 66485 185051
rect 66513 185023 66547 185051
rect 66575 185023 66609 185051
rect 66637 185023 66671 185051
rect 66699 185023 75485 185051
rect 75513 185023 75547 185051
rect 75575 185023 75609 185051
rect 75637 185023 75671 185051
rect 75699 185023 84485 185051
rect 84513 185023 84547 185051
rect 84575 185023 84609 185051
rect 84637 185023 84671 185051
rect 84699 185023 93485 185051
rect 93513 185023 93547 185051
rect 93575 185023 93609 185051
rect 93637 185023 93671 185051
rect 93699 185023 102485 185051
rect 102513 185023 102547 185051
rect 102575 185023 102609 185051
rect 102637 185023 102671 185051
rect 102699 185023 111485 185051
rect 111513 185023 111547 185051
rect 111575 185023 111609 185051
rect 111637 185023 111671 185051
rect 111699 185023 120485 185051
rect 120513 185023 120547 185051
rect 120575 185023 120609 185051
rect 120637 185023 120671 185051
rect 120699 185023 129485 185051
rect 129513 185023 129547 185051
rect 129575 185023 129609 185051
rect 129637 185023 129671 185051
rect 129699 185023 138485 185051
rect 138513 185023 138547 185051
rect 138575 185023 138609 185051
rect 138637 185023 138671 185051
rect 138699 185023 147485 185051
rect 147513 185023 147547 185051
rect 147575 185023 147609 185051
rect 147637 185023 147671 185051
rect 147699 185023 156485 185051
rect 156513 185023 156547 185051
rect 156575 185023 156609 185051
rect 156637 185023 156671 185051
rect 156699 185023 165485 185051
rect 165513 185023 165547 185051
rect 165575 185023 165609 185051
rect 165637 185023 165671 185051
rect 165699 185023 174485 185051
rect 174513 185023 174547 185051
rect 174575 185023 174609 185051
rect 174637 185023 174671 185051
rect 174699 185023 183485 185051
rect 183513 185023 183547 185051
rect 183575 185023 183609 185051
rect 183637 185023 183671 185051
rect 183699 185023 192485 185051
rect 192513 185023 192547 185051
rect 192575 185023 192609 185051
rect 192637 185023 192671 185051
rect 192699 185023 201485 185051
rect 201513 185023 201547 185051
rect 201575 185023 201609 185051
rect 201637 185023 201671 185051
rect 201699 185023 210485 185051
rect 210513 185023 210547 185051
rect 210575 185023 210609 185051
rect 210637 185023 210671 185051
rect 210699 185023 219485 185051
rect 219513 185023 219547 185051
rect 219575 185023 219609 185051
rect 219637 185023 219671 185051
rect 219699 185023 228485 185051
rect 228513 185023 228547 185051
rect 228575 185023 228609 185051
rect 228637 185023 228671 185051
rect 228699 185023 237485 185051
rect 237513 185023 237547 185051
rect 237575 185023 237609 185051
rect 237637 185023 237671 185051
rect 237699 185023 246485 185051
rect 246513 185023 246547 185051
rect 246575 185023 246609 185051
rect 246637 185023 246671 185051
rect 246699 185023 255485 185051
rect 255513 185023 255547 185051
rect 255575 185023 255609 185051
rect 255637 185023 255671 185051
rect 255699 185023 264485 185051
rect 264513 185023 264547 185051
rect 264575 185023 264609 185051
rect 264637 185023 264671 185051
rect 264699 185023 273485 185051
rect 273513 185023 273547 185051
rect 273575 185023 273609 185051
rect 273637 185023 273671 185051
rect 273699 185023 282485 185051
rect 282513 185023 282547 185051
rect 282575 185023 282609 185051
rect 282637 185023 282671 185051
rect 282699 185023 291485 185051
rect 291513 185023 291547 185051
rect 291575 185023 291609 185051
rect 291637 185023 291671 185051
rect 291699 185023 298728 185051
rect 298756 185023 298790 185051
rect 298818 185023 298852 185051
rect 298880 185023 298914 185051
rect 298942 185023 298990 185051
rect -958 184989 298990 185023
rect -958 184961 -910 184989
rect -882 184961 -848 184989
rect -820 184961 -786 184989
rect -758 184961 -724 184989
rect -696 184961 3485 184989
rect 3513 184961 3547 184989
rect 3575 184961 3609 184989
rect 3637 184961 3671 184989
rect 3699 184961 12485 184989
rect 12513 184961 12547 184989
rect 12575 184961 12609 184989
rect 12637 184961 12671 184989
rect 12699 184961 21485 184989
rect 21513 184961 21547 184989
rect 21575 184961 21609 184989
rect 21637 184961 21671 184989
rect 21699 184961 30485 184989
rect 30513 184961 30547 184989
rect 30575 184961 30609 184989
rect 30637 184961 30671 184989
rect 30699 184961 39485 184989
rect 39513 184961 39547 184989
rect 39575 184961 39609 184989
rect 39637 184961 39671 184989
rect 39699 184961 48485 184989
rect 48513 184961 48547 184989
rect 48575 184961 48609 184989
rect 48637 184961 48671 184989
rect 48699 184961 57485 184989
rect 57513 184961 57547 184989
rect 57575 184961 57609 184989
rect 57637 184961 57671 184989
rect 57699 184961 66485 184989
rect 66513 184961 66547 184989
rect 66575 184961 66609 184989
rect 66637 184961 66671 184989
rect 66699 184961 75485 184989
rect 75513 184961 75547 184989
rect 75575 184961 75609 184989
rect 75637 184961 75671 184989
rect 75699 184961 84485 184989
rect 84513 184961 84547 184989
rect 84575 184961 84609 184989
rect 84637 184961 84671 184989
rect 84699 184961 93485 184989
rect 93513 184961 93547 184989
rect 93575 184961 93609 184989
rect 93637 184961 93671 184989
rect 93699 184961 102485 184989
rect 102513 184961 102547 184989
rect 102575 184961 102609 184989
rect 102637 184961 102671 184989
rect 102699 184961 111485 184989
rect 111513 184961 111547 184989
rect 111575 184961 111609 184989
rect 111637 184961 111671 184989
rect 111699 184961 120485 184989
rect 120513 184961 120547 184989
rect 120575 184961 120609 184989
rect 120637 184961 120671 184989
rect 120699 184961 129485 184989
rect 129513 184961 129547 184989
rect 129575 184961 129609 184989
rect 129637 184961 129671 184989
rect 129699 184961 138485 184989
rect 138513 184961 138547 184989
rect 138575 184961 138609 184989
rect 138637 184961 138671 184989
rect 138699 184961 147485 184989
rect 147513 184961 147547 184989
rect 147575 184961 147609 184989
rect 147637 184961 147671 184989
rect 147699 184961 156485 184989
rect 156513 184961 156547 184989
rect 156575 184961 156609 184989
rect 156637 184961 156671 184989
rect 156699 184961 165485 184989
rect 165513 184961 165547 184989
rect 165575 184961 165609 184989
rect 165637 184961 165671 184989
rect 165699 184961 174485 184989
rect 174513 184961 174547 184989
rect 174575 184961 174609 184989
rect 174637 184961 174671 184989
rect 174699 184961 183485 184989
rect 183513 184961 183547 184989
rect 183575 184961 183609 184989
rect 183637 184961 183671 184989
rect 183699 184961 192485 184989
rect 192513 184961 192547 184989
rect 192575 184961 192609 184989
rect 192637 184961 192671 184989
rect 192699 184961 201485 184989
rect 201513 184961 201547 184989
rect 201575 184961 201609 184989
rect 201637 184961 201671 184989
rect 201699 184961 210485 184989
rect 210513 184961 210547 184989
rect 210575 184961 210609 184989
rect 210637 184961 210671 184989
rect 210699 184961 219485 184989
rect 219513 184961 219547 184989
rect 219575 184961 219609 184989
rect 219637 184961 219671 184989
rect 219699 184961 228485 184989
rect 228513 184961 228547 184989
rect 228575 184961 228609 184989
rect 228637 184961 228671 184989
rect 228699 184961 237485 184989
rect 237513 184961 237547 184989
rect 237575 184961 237609 184989
rect 237637 184961 237671 184989
rect 237699 184961 246485 184989
rect 246513 184961 246547 184989
rect 246575 184961 246609 184989
rect 246637 184961 246671 184989
rect 246699 184961 255485 184989
rect 255513 184961 255547 184989
rect 255575 184961 255609 184989
rect 255637 184961 255671 184989
rect 255699 184961 264485 184989
rect 264513 184961 264547 184989
rect 264575 184961 264609 184989
rect 264637 184961 264671 184989
rect 264699 184961 273485 184989
rect 273513 184961 273547 184989
rect 273575 184961 273609 184989
rect 273637 184961 273671 184989
rect 273699 184961 282485 184989
rect 282513 184961 282547 184989
rect 282575 184961 282609 184989
rect 282637 184961 282671 184989
rect 282699 184961 291485 184989
rect 291513 184961 291547 184989
rect 291575 184961 291609 184989
rect 291637 184961 291671 184989
rect 291699 184961 298728 184989
rect 298756 184961 298790 184989
rect 298818 184961 298852 184989
rect 298880 184961 298914 184989
rect 298942 184961 298990 184989
rect -958 184913 298990 184961
rect -958 182175 298990 182223
rect -958 182147 -430 182175
rect -402 182147 -368 182175
rect -340 182147 -306 182175
rect -278 182147 -244 182175
rect -216 182147 1625 182175
rect 1653 182147 1687 182175
rect 1715 182147 1749 182175
rect 1777 182147 1811 182175
rect 1839 182147 10625 182175
rect 10653 182147 10687 182175
rect 10715 182147 10749 182175
rect 10777 182147 10811 182175
rect 10839 182147 19625 182175
rect 19653 182147 19687 182175
rect 19715 182147 19749 182175
rect 19777 182147 19811 182175
rect 19839 182147 28625 182175
rect 28653 182147 28687 182175
rect 28715 182147 28749 182175
rect 28777 182147 28811 182175
rect 28839 182147 37625 182175
rect 37653 182147 37687 182175
rect 37715 182147 37749 182175
rect 37777 182147 37811 182175
rect 37839 182147 46625 182175
rect 46653 182147 46687 182175
rect 46715 182147 46749 182175
rect 46777 182147 46811 182175
rect 46839 182147 52259 182175
rect 52287 182147 52321 182175
rect 52349 182147 67619 182175
rect 67647 182147 67681 182175
rect 67709 182147 82979 182175
rect 83007 182147 83041 182175
rect 83069 182147 98339 182175
rect 98367 182147 98401 182175
rect 98429 182147 113699 182175
rect 113727 182147 113761 182175
rect 113789 182147 129059 182175
rect 129087 182147 129121 182175
rect 129149 182147 144419 182175
rect 144447 182147 144481 182175
rect 144509 182147 154625 182175
rect 154653 182147 154687 182175
rect 154715 182147 154749 182175
rect 154777 182147 154811 182175
rect 154839 182147 163625 182175
rect 163653 182147 163687 182175
rect 163715 182147 163749 182175
rect 163777 182147 163811 182175
rect 163839 182147 172625 182175
rect 172653 182147 172687 182175
rect 172715 182147 172749 182175
rect 172777 182147 172811 182175
rect 172839 182147 181625 182175
rect 181653 182147 181687 182175
rect 181715 182147 181749 182175
rect 181777 182147 181811 182175
rect 181839 182147 190625 182175
rect 190653 182147 190687 182175
rect 190715 182147 190749 182175
rect 190777 182147 190811 182175
rect 190839 182147 199625 182175
rect 199653 182147 199687 182175
rect 199715 182147 199749 182175
rect 199777 182147 199811 182175
rect 199839 182147 208625 182175
rect 208653 182147 208687 182175
rect 208715 182147 208749 182175
rect 208777 182147 208811 182175
rect 208839 182147 217625 182175
rect 217653 182147 217687 182175
rect 217715 182147 217749 182175
rect 217777 182147 217811 182175
rect 217839 182147 226625 182175
rect 226653 182147 226687 182175
rect 226715 182147 226749 182175
rect 226777 182147 226811 182175
rect 226839 182147 235625 182175
rect 235653 182147 235687 182175
rect 235715 182147 235749 182175
rect 235777 182147 235811 182175
rect 235839 182147 244625 182175
rect 244653 182147 244687 182175
rect 244715 182147 244749 182175
rect 244777 182147 244811 182175
rect 244839 182147 253625 182175
rect 253653 182147 253687 182175
rect 253715 182147 253749 182175
rect 253777 182147 253811 182175
rect 253839 182147 262625 182175
rect 262653 182147 262687 182175
rect 262715 182147 262749 182175
rect 262777 182147 262811 182175
rect 262839 182147 271625 182175
rect 271653 182147 271687 182175
rect 271715 182147 271749 182175
rect 271777 182147 271811 182175
rect 271839 182147 280625 182175
rect 280653 182147 280687 182175
rect 280715 182147 280749 182175
rect 280777 182147 280811 182175
rect 280839 182147 289625 182175
rect 289653 182147 289687 182175
rect 289715 182147 289749 182175
rect 289777 182147 289811 182175
rect 289839 182147 298248 182175
rect 298276 182147 298310 182175
rect 298338 182147 298372 182175
rect 298400 182147 298434 182175
rect 298462 182147 298990 182175
rect -958 182113 298990 182147
rect -958 182085 -430 182113
rect -402 182085 -368 182113
rect -340 182085 -306 182113
rect -278 182085 -244 182113
rect -216 182085 1625 182113
rect 1653 182085 1687 182113
rect 1715 182085 1749 182113
rect 1777 182085 1811 182113
rect 1839 182085 10625 182113
rect 10653 182085 10687 182113
rect 10715 182085 10749 182113
rect 10777 182085 10811 182113
rect 10839 182085 19625 182113
rect 19653 182085 19687 182113
rect 19715 182085 19749 182113
rect 19777 182085 19811 182113
rect 19839 182085 28625 182113
rect 28653 182085 28687 182113
rect 28715 182085 28749 182113
rect 28777 182085 28811 182113
rect 28839 182085 37625 182113
rect 37653 182085 37687 182113
rect 37715 182085 37749 182113
rect 37777 182085 37811 182113
rect 37839 182085 46625 182113
rect 46653 182085 46687 182113
rect 46715 182085 46749 182113
rect 46777 182085 46811 182113
rect 46839 182085 52259 182113
rect 52287 182085 52321 182113
rect 52349 182085 67619 182113
rect 67647 182085 67681 182113
rect 67709 182085 82979 182113
rect 83007 182085 83041 182113
rect 83069 182085 98339 182113
rect 98367 182085 98401 182113
rect 98429 182085 113699 182113
rect 113727 182085 113761 182113
rect 113789 182085 129059 182113
rect 129087 182085 129121 182113
rect 129149 182085 144419 182113
rect 144447 182085 144481 182113
rect 144509 182085 154625 182113
rect 154653 182085 154687 182113
rect 154715 182085 154749 182113
rect 154777 182085 154811 182113
rect 154839 182085 163625 182113
rect 163653 182085 163687 182113
rect 163715 182085 163749 182113
rect 163777 182085 163811 182113
rect 163839 182085 172625 182113
rect 172653 182085 172687 182113
rect 172715 182085 172749 182113
rect 172777 182085 172811 182113
rect 172839 182085 181625 182113
rect 181653 182085 181687 182113
rect 181715 182085 181749 182113
rect 181777 182085 181811 182113
rect 181839 182085 190625 182113
rect 190653 182085 190687 182113
rect 190715 182085 190749 182113
rect 190777 182085 190811 182113
rect 190839 182085 199625 182113
rect 199653 182085 199687 182113
rect 199715 182085 199749 182113
rect 199777 182085 199811 182113
rect 199839 182085 208625 182113
rect 208653 182085 208687 182113
rect 208715 182085 208749 182113
rect 208777 182085 208811 182113
rect 208839 182085 217625 182113
rect 217653 182085 217687 182113
rect 217715 182085 217749 182113
rect 217777 182085 217811 182113
rect 217839 182085 226625 182113
rect 226653 182085 226687 182113
rect 226715 182085 226749 182113
rect 226777 182085 226811 182113
rect 226839 182085 235625 182113
rect 235653 182085 235687 182113
rect 235715 182085 235749 182113
rect 235777 182085 235811 182113
rect 235839 182085 244625 182113
rect 244653 182085 244687 182113
rect 244715 182085 244749 182113
rect 244777 182085 244811 182113
rect 244839 182085 253625 182113
rect 253653 182085 253687 182113
rect 253715 182085 253749 182113
rect 253777 182085 253811 182113
rect 253839 182085 262625 182113
rect 262653 182085 262687 182113
rect 262715 182085 262749 182113
rect 262777 182085 262811 182113
rect 262839 182085 271625 182113
rect 271653 182085 271687 182113
rect 271715 182085 271749 182113
rect 271777 182085 271811 182113
rect 271839 182085 280625 182113
rect 280653 182085 280687 182113
rect 280715 182085 280749 182113
rect 280777 182085 280811 182113
rect 280839 182085 289625 182113
rect 289653 182085 289687 182113
rect 289715 182085 289749 182113
rect 289777 182085 289811 182113
rect 289839 182085 298248 182113
rect 298276 182085 298310 182113
rect 298338 182085 298372 182113
rect 298400 182085 298434 182113
rect 298462 182085 298990 182113
rect -958 182051 298990 182085
rect -958 182023 -430 182051
rect -402 182023 -368 182051
rect -340 182023 -306 182051
rect -278 182023 -244 182051
rect -216 182023 1625 182051
rect 1653 182023 1687 182051
rect 1715 182023 1749 182051
rect 1777 182023 1811 182051
rect 1839 182023 10625 182051
rect 10653 182023 10687 182051
rect 10715 182023 10749 182051
rect 10777 182023 10811 182051
rect 10839 182023 19625 182051
rect 19653 182023 19687 182051
rect 19715 182023 19749 182051
rect 19777 182023 19811 182051
rect 19839 182023 28625 182051
rect 28653 182023 28687 182051
rect 28715 182023 28749 182051
rect 28777 182023 28811 182051
rect 28839 182023 37625 182051
rect 37653 182023 37687 182051
rect 37715 182023 37749 182051
rect 37777 182023 37811 182051
rect 37839 182023 46625 182051
rect 46653 182023 46687 182051
rect 46715 182023 46749 182051
rect 46777 182023 46811 182051
rect 46839 182023 52259 182051
rect 52287 182023 52321 182051
rect 52349 182023 67619 182051
rect 67647 182023 67681 182051
rect 67709 182023 82979 182051
rect 83007 182023 83041 182051
rect 83069 182023 98339 182051
rect 98367 182023 98401 182051
rect 98429 182023 113699 182051
rect 113727 182023 113761 182051
rect 113789 182023 129059 182051
rect 129087 182023 129121 182051
rect 129149 182023 144419 182051
rect 144447 182023 144481 182051
rect 144509 182023 154625 182051
rect 154653 182023 154687 182051
rect 154715 182023 154749 182051
rect 154777 182023 154811 182051
rect 154839 182023 163625 182051
rect 163653 182023 163687 182051
rect 163715 182023 163749 182051
rect 163777 182023 163811 182051
rect 163839 182023 172625 182051
rect 172653 182023 172687 182051
rect 172715 182023 172749 182051
rect 172777 182023 172811 182051
rect 172839 182023 181625 182051
rect 181653 182023 181687 182051
rect 181715 182023 181749 182051
rect 181777 182023 181811 182051
rect 181839 182023 190625 182051
rect 190653 182023 190687 182051
rect 190715 182023 190749 182051
rect 190777 182023 190811 182051
rect 190839 182023 199625 182051
rect 199653 182023 199687 182051
rect 199715 182023 199749 182051
rect 199777 182023 199811 182051
rect 199839 182023 208625 182051
rect 208653 182023 208687 182051
rect 208715 182023 208749 182051
rect 208777 182023 208811 182051
rect 208839 182023 217625 182051
rect 217653 182023 217687 182051
rect 217715 182023 217749 182051
rect 217777 182023 217811 182051
rect 217839 182023 226625 182051
rect 226653 182023 226687 182051
rect 226715 182023 226749 182051
rect 226777 182023 226811 182051
rect 226839 182023 235625 182051
rect 235653 182023 235687 182051
rect 235715 182023 235749 182051
rect 235777 182023 235811 182051
rect 235839 182023 244625 182051
rect 244653 182023 244687 182051
rect 244715 182023 244749 182051
rect 244777 182023 244811 182051
rect 244839 182023 253625 182051
rect 253653 182023 253687 182051
rect 253715 182023 253749 182051
rect 253777 182023 253811 182051
rect 253839 182023 262625 182051
rect 262653 182023 262687 182051
rect 262715 182023 262749 182051
rect 262777 182023 262811 182051
rect 262839 182023 271625 182051
rect 271653 182023 271687 182051
rect 271715 182023 271749 182051
rect 271777 182023 271811 182051
rect 271839 182023 280625 182051
rect 280653 182023 280687 182051
rect 280715 182023 280749 182051
rect 280777 182023 280811 182051
rect 280839 182023 289625 182051
rect 289653 182023 289687 182051
rect 289715 182023 289749 182051
rect 289777 182023 289811 182051
rect 289839 182023 298248 182051
rect 298276 182023 298310 182051
rect 298338 182023 298372 182051
rect 298400 182023 298434 182051
rect 298462 182023 298990 182051
rect -958 181989 298990 182023
rect -958 181961 -430 181989
rect -402 181961 -368 181989
rect -340 181961 -306 181989
rect -278 181961 -244 181989
rect -216 181961 1625 181989
rect 1653 181961 1687 181989
rect 1715 181961 1749 181989
rect 1777 181961 1811 181989
rect 1839 181961 10625 181989
rect 10653 181961 10687 181989
rect 10715 181961 10749 181989
rect 10777 181961 10811 181989
rect 10839 181961 19625 181989
rect 19653 181961 19687 181989
rect 19715 181961 19749 181989
rect 19777 181961 19811 181989
rect 19839 181961 28625 181989
rect 28653 181961 28687 181989
rect 28715 181961 28749 181989
rect 28777 181961 28811 181989
rect 28839 181961 37625 181989
rect 37653 181961 37687 181989
rect 37715 181961 37749 181989
rect 37777 181961 37811 181989
rect 37839 181961 46625 181989
rect 46653 181961 46687 181989
rect 46715 181961 46749 181989
rect 46777 181961 46811 181989
rect 46839 181961 52259 181989
rect 52287 181961 52321 181989
rect 52349 181961 67619 181989
rect 67647 181961 67681 181989
rect 67709 181961 82979 181989
rect 83007 181961 83041 181989
rect 83069 181961 98339 181989
rect 98367 181961 98401 181989
rect 98429 181961 113699 181989
rect 113727 181961 113761 181989
rect 113789 181961 129059 181989
rect 129087 181961 129121 181989
rect 129149 181961 144419 181989
rect 144447 181961 144481 181989
rect 144509 181961 154625 181989
rect 154653 181961 154687 181989
rect 154715 181961 154749 181989
rect 154777 181961 154811 181989
rect 154839 181961 163625 181989
rect 163653 181961 163687 181989
rect 163715 181961 163749 181989
rect 163777 181961 163811 181989
rect 163839 181961 172625 181989
rect 172653 181961 172687 181989
rect 172715 181961 172749 181989
rect 172777 181961 172811 181989
rect 172839 181961 181625 181989
rect 181653 181961 181687 181989
rect 181715 181961 181749 181989
rect 181777 181961 181811 181989
rect 181839 181961 190625 181989
rect 190653 181961 190687 181989
rect 190715 181961 190749 181989
rect 190777 181961 190811 181989
rect 190839 181961 199625 181989
rect 199653 181961 199687 181989
rect 199715 181961 199749 181989
rect 199777 181961 199811 181989
rect 199839 181961 208625 181989
rect 208653 181961 208687 181989
rect 208715 181961 208749 181989
rect 208777 181961 208811 181989
rect 208839 181961 217625 181989
rect 217653 181961 217687 181989
rect 217715 181961 217749 181989
rect 217777 181961 217811 181989
rect 217839 181961 226625 181989
rect 226653 181961 226687 181989
rect 226715 181961 226749 181989
rect 226777 181961 226811 181989
rect 226839 181961 235625 181989
rect 235653 181961 235687 181989
rect 235715 181961 235749 181989
rect 235777 181961 235811 181989
rect 235839 181961 244625 181989
rect 244653 181961 244687 181989
rect 244715 181961 244749 181989
rect 244777 181961 244811 181989
rect 244839 181961 253625 181989
rect 253653 181961 253687 181989
rect 253715 181961 253749 181989
rect 253777 181961 253811 181989
rect 253839 181961 262625 181989
rect 262653 181961 262687 181989
rect 262715 181961 262749 181989
rect 262777 181961 262811 181989
rect 262839 181961 271625 181989
rect 271653 181961 271687 181989
rect 271715 181961 271749 181989
rect 271777 181961 271811 181989
rect 271839 181961 280625 181989
rect 280653 181961 280687 181989
rect 280715 181961 280749 181989
rect 280777 181961 280811 181989
rect 280839 181961 289625 181989
rect 289653 181961 289687 181989
rect 289715 181961 289749 181989
rect 289777 181961 289811 181989
rect 289839 181961 298248 181989
rect 298276 181961 298310 181989
rect 298338 181961 298372 181989
rect 298400 181961 298434 181989
rect 298462 181961 298990 181989
rect -958 181913 298990 181961
rect -958 176175 298990 176223
rect -958 176147 -910 176175
rect -882 176147 -848 176175
rect -820 176147 -786 176175
rect -758 176147 -724 176175
rect -696 176147 3485 176175
rect 3513 176147 3547 176175
rect 3575 176147 3609 176175
rect 3637 176147 3671 176175
rect 3699 176147 12485 176175
rect 12513 176147 12547 176175
rect 12575 176147 12609 176175
rect 12637 176147 12671 176175
rect 12699 176147 21485 176175
rect 21513 176147 21547 176175
rect 21575 176147 21609 176175
rect 21637 176147 21671 176175
rect 21699 176147 30485 176175
rect 30513 176147 30547 176175
rect 30575 176147 30609 176175
rect 30637 176147 30671 176175
rect 30699 176147 39485 176175
rect 39513 176147 39547 176175
rect 39575 176147 39609 176175
rect 39637 176147 39671 176175
rect 39699 176147 48485 176175
rect 48513 176147 48547 176175
rect 48575 176147 48609 176175
rect 48637 176147 48671 176175
rect 48699 176147 59939 176175
rect 59967 176147 60001 176175
rect 60029 176147 75299 176175
rect 75327 176147 75361 176175
rect 75389 176147 90659 176175
rect 90687 176147 90721 176175
rect 90749 176147 106019 176175
rect 106047 176147 106081 176175
rect 106109 176147 121379 176175
rect 121407 176147 121441 176175
rect 121469 176147 136739 176175
rect 136767 176147 136801 176175
rect 136829 176147 156485 176175
rect 156513 176147 156547 176175
rect 156575 176147 156609 176175
rect 156637 176147 156671 176175
rect 156699 176147 165485 176175
rect 165513 176147 165547 176175
rect 165575 176147 165609 176175
rect 165637 176147 165671 176175
rect 165699 176147 174485 176175
rect 174513 176147 174547 176175
rect 174575 176147 174609 176175
rect 174637 176147 174671 176175
rect 174699 176147 183485 176175
rect 183513 176147 183547 176175
rect 183575 176147 183609 176175
rect 183637 176147 183671 176175
rect 183699 176147 192485 176175
rect 192513 176147 192547 176175
rect 192575 176147 192609 176175
rect 192637 176147 192671 176175
rect 192699 176147 201485 176175
rect 201513 176147 201547 176175
rect 201575 176147 201609 176175
rect 201637 176147 201671 176175
rect 201699 176147 210485 176175
rect 210513 176147 210547 176175
rect 210575 176147 210609 176175
rect 210637 176147 210671 176175
rect 210699 176147 219485 176175
rect 219513 176147 219547 176175
rect 219575 176147 219609 176175
rect 219637 176147 219671 176175
rect 219699 176147 228485 176175
rect 228513 176147 228547 176175
rect 228575 176147 228609 176175
rect 228637 176147 228671 176175
rect 228699 176147 237485 176175
rect 237513 176147 237547 176175
rect 237575 176147 237609 176175
rect 237637 176147 237671 176175
rect 237699 176147 246485 176175
rect 246513 176147 246547 176175
rect 246575 176147 246609 176175
rect 246637 176147 246671 176175
rect 246699 176147 255485 176175
rect 255513 176147 255547 176175
rect 255575 176147 255609 176175
rect 255637 176147 255671 176175
rect 255699 176147 264485 176175
rect 264513 176147 264547 176175
rect 264575 176147 264609 176175
rect 264637 176147 264671 176175
rect 264699 176147 273485 176175
rect 273513 176147 273547 176175
rect 273575 176147 273609 176175
rect 273637 176147 273671 176175
rect 273699 176147 282485 176175
rect 282513 176147 282547 176175
rect 282575 176147 282609 176175
rect 282637 176147 282671 176175
rect 282699 176147 291485 176175
rect 291513 176147 291547 176175
rect 291575 176147 291609 176175
rect 291637 176147 291671 176175
rect 291699 176147 298728 176175
rect 298756 176147 298790 176175
rect 298818 176147 298852 176175
rect 298880 176147 298914 176175
rect 298942 176147 298990 176175
rect -958 176113 298990 176147
rect -958 176085 -910 176113
rect -882 176085 -848 176113
rect -820 176085 -786 176113
rect -758 176085 -724 176113
rect -696 176085 3485 176113
rect 3513 176085 3547 176113
rect 3575 176085 3609 176113
rect 3637 176085 3671 176113
rect 3699 176085 12485 176113
rect 12513 176085 12547 176113
rect 12575 176085 12609 176113
rect 12637 176085 12671 176113
rect 12699 176085 21485 176113
rect 21513 176085 21547 176113
rect 21575 176085 21609 176113
rect 21637 176085 21671 176113
rect 21699 176085 30485 176113
rect 30513 176085 30547 176113
rect 30575 176085 30609 176113
rect 30637 176085 30671 176113
rect 30699 176085 39485 176113
rect 39513 176085 39547 176113
rect 39575 176085 39609 176113
rect 39637 176085 39671 176113
rect 39699 176085 48485 176113
rect 48513 176085 48547 176113
rect 48575 176085 48609 176113
rect 48637 176085 48671 176113
rect 48699 176085 59939 176113
rect 59967 176085 60001 176113
rect 60029 176085 75299 176113
rect 75327 176085 75361 176113
rect 75389 176085 90659 176113
rect 90687 176085 90721 176113
rect 90749 176085 106019 176113
rect 106047 176085 106081 176113
rect 106109 176085 121379 176113
rect 121407 176085 121441 176113
rect 121469 176085 136739 176113
rect 136767 176085 136801 176113
rect 136829 176085 156485 176113
rect 156513 176085 156547 176113
rect 156575 176085 156609 176113
rect 156637 176085 156671 176113
rect 156699 176085 165485 176113
rect 165513 176085 165547 176113
rect 165575 176085 165609 176113
rect 165637 176085 165671 176113
rect 165699 176085 174485 176113
rect 174513 176085 174547 176113
rect 174575 176085 174609 176113
rect 174637 176085 174671 176113
rect 174699 176085 183485 176113
rect 183513 176085 183547 176113
rect 183575 176085 183609 176113
rect 183637 176085 183671 176113
rect 183699 176085 192485 176113
rect 192513 176085 192547 176113
rect 192575 176085 192609 176113
rect 192637 176085 192671 176113
rect 192699 176085 201485 176113
rect 201513 176085 201547 176113
rect 201575 176085 201609 176113
rect 201637 176085 201671 176113
rect 201699 176085 210485 176113
rect 210513 176085 210547 176113
rect 210575 176085 210609 176113
rect 210637 176085 210671 176113
rect 210699 176085 219485 176113
rect 219513 176085 219547 176113
rect 219575 176085 219609 176113
rect 219637 176085 219671 176113
rect 219699 176085 228485 176113
rect 228513 176085 228547 176113
rect 228575 176085 228609 176113
rect 228637 176085 228671 176113
rect 228699 176085 237485 176113
rect 237513 176085 237547 176113
rect 237575 176085 237609 176113
rect 237637 176085 237671 176113
rect 237699 176085 246485 176113
rect 246513 176085 246547 176113
rect 246575 176085 246609 176113
rect 246637 176085 246671 176113
rect 246699 176085 255485 176113
rect 255513 176085 255547 176113
rect 255575 176085 255609 176113
rect 255637 176085 255671 176113
rect 255699 176085 264485 176113
rect 264513 176085 264547 176113
rect 264575 176085 264609 176113
rect 264637 176085 264671 176113
rect 264699 176085 273485 176113
rect 273513 176085 273547 176113
rect 273575 176085 273609 176113
rect 273637 176085 273671 176113
rect 273699 176085 282485 176113
rect 282513 176085 282547 176113
rect 282575 176085 282609 176113
rect 282637 176085 282671 176113
rect 282699 176085 291485 176113
rect 291513 176085 291547 176113
rect 291575 176085 291609 176113
rect 291637 176085 291671 176113
rect 291699 176085 298728 176113
rect 298756 176085 298790 176113
rect 298818 176085 298852 176113
rect 298880 176085 298914 176113
rect 298942 176085 298990 176113
rect -958 176051 298990 176085
rect -958 176023 -910 176051
rect -882 176023 -848 176051
rect -820 176023 -786 176051
rect -758 176023 -724 176051
rect -696 176023 3485 176051
rect 3513 176023 3547 176051
rect 3575 176023 3609 176051
rect 3637 176023 3671 176051
rect 3699 176023 12485 176051
rect 12513 176023 12547 176051
rect 12575 176023 12609 176051
rect 12637 176023 12671 176051
rect 12699 176023 21485 176051
rect 21513 176023 21547 176051
rect 21575 176023 21609 176051
rect 21637 176023 21671 176051
rect 21699 176023 30485 176051
rect 30513 176023 30547 176051
rect 30575 176023 30609 176051
rect 30637 176023 30671 176051
rect 30699 176023 39485 176051
rect 39513 176023 39547 176051
rect 39575 176023 39609 176051
rect 39637 176023 39671 176051
rect 39699 176023 48485 176051
rect 48513 176023 48547 176051
rect 48575 176023 48609 176051
rect 48637 176023 48671 176051
rect 48699 176023 59939 176051
rect 59967 176023 60001 176051
rect 60029 176023 75299 176051
rect 75327 176023 75361 176051
rect 75389 176023 90659 176051
rect 90687 176023 90721 176051
rect 90749 176023 106019 176051
rect 106047 176023 106081 176051
rect 106109 176023 121379 176051
rect 121407 176023 121441 176051
rect 121469 176023 136739 176051
rect 136767 176023 136801 176051
rect 136829 176023 156485 176051
rect 156513 176023 156547 176051
rect 156575 176023 156609 176051
rect 156637 176023 156671 176051
rect 156699 176023 165485 176051
rect 165513 176023 165547 176051
rect 165575 176023 165609 176051
rect 165637 176023 165671 176051
rect 165699 176023 174485 176051
rect 174513 176023 174547 176051
rect 174575 176023 174609 176051
rect 174637 176023 174671 176051
rect 174699 176023 183485 176051
rect 183513 176023 183547 176051
rect 183575 176023 183609 176051
rect 183637 176023 183671 176051
rect 183699 176023 192485 176051
rect 192513 176023 192547 176051
rect 192575 176023 192609 176051
rect 192637 176023 192671 176051
rect 192699 176023 201485 176051
rect 201513 176023 201547 176051
rect 201575 176023 201609 176051
rect 201637 176023 201671 176051
rect 201699 176023 210485 176051
rect 210513 176023 210547 176051
rect 210575 176023 210609 176051
rect 210637 176023 210671 176051
rect 210699 176023 219485 176051
rect 219513 176023 219547 176051
rect 219575 176023 219609 176051
rect 219637 176023 219671 176051
rect 219699 176023 228485 176051
rect 228513 176023 228547 176051
rect 228575 176023 228609 176051
rect 228637 176023 228671 176051
rect 228699 176023 237485 176051
rect 237513 176023 237547 176051
rect 237575 176023 237609 176051
rect 237637 176023 237671 176051
rect 237699 176023 246485 176051
rect 246513 176023 246547 176051
rect 246575 176023 246609 176051
rect 246637 176023 246671 176051
rect 246699 176023 255485 176051
rect 255513 176023 255547 176051
rect 255575 176023 255609 176051
rect 255637 176023 255671 176051
rect 255699 176023 264485 176051
rect 264513 176023 264547 176051
rect 264575 176023 264609 176051
rect 264637 176023 264671 176051
rect 264699 176023 273485 176051
rect 273513 176023 273547 176051
rect 273575 176023 273609 176051
rect 273637 176023 273671 176051
rect 273699 176023 282485 176051
rect 282513 176023 282547 176051
rect 282575 176023 282609 176051
rect 282637 176023 282671 176051
rect 282699 176023 291485 176051
rect 291513 176023 291547 176051
rect 291575 176023 291609 176051
rect 291637 176023 291671 176051
rect 291699 176023 298728 176051
rect 298756 176023 298790 176051
rect 298818 176023 298852 176051
rect 298880 176023 298914 176051
rect 298942 176023 298990 176051
rect -958 175989 298990 176023
rect -958 175961 -910 175989
rect -882 175961 -848 175989
rect -820 175961 -786 175989
rect -758 175961 -724 175989
rect -696 175961 3485 175989
rect 3513 175961 3547 175989
rect 3575 175961 3609 175989
rect 3637 175961 3671 175989
rect 3699 175961 12485 175989
rect 12513 175961 12547 175989
rect 12575 175961 12609 175989
rect 12637 175961 12671 175989
rect 12699 175961 21485 175989
rect 21513 175961 21547 175989
rect 21575 175961 21609 175989
rect 21637 175961 21671 175989
rect 21699 175961 30485 175989
rect 30513 175961 30547 175989
rect 30575 175961 30609 175989
rect 30637 175961 30671 175989
rect 30699 175961 39485 175989
rect 39513 175961 39547 175989
rect 39575 175961 39609 175989
rect 39637 175961 39671 175989
rect 39699 175961 48485 175989
rect 48513 175961 48547 175989
rect 48575 175961 48609 175989
rect 48637 175961 48671 175989
rect 48699 175961 59939 175989
rect 59967 175961 60001 175989
rect 60029 175961 75299 175989
rect 75327 175961 75361 175989
rect 75389 175961 90659 175989
rect 90687 175961 90721 175989
rect 90749 175961 106019 175989
rect 106047 175961 106081 175989
rect 106109 175961 121379 175989
rect 121407 175961 121441 175989
rect 121469 175961 136739 175989
rect 136767 175961 136801 175989
rect 136829 175961 156485 175989
rect 156513 175961 156547 175989
rect 156575 175961 156609 175989
rect 156637 175961 156671 175989
rect 156699 175961 165485 175989
rect 165513 175961 165547 175989
rect 165575 175961 165609 175989
rect 165637 175961 165671 175989
rect 165699 175961 174485 175989
rect 174513 175961 174547 175989
rect 174575 175961 174609 175989
rect 174637 175961 174671 175989
rect 174699 175961 183485 175989
rect 183513 175961 183547 175989
rect 183575 175961 183609 175989
rect 183637 175961 183671 175989
rect 183699 175961 192485 175989
rect 192513 175961 192547 175989
rect 192575 175961 192609 175989
rect 192637 175961 192671 175989
rect 192699 175961 201485 175989
rect 201513 175961 201547 175989
rect 201575 175961 201609 175989
rect 201637 175961 201671 175989
rect 201699 175961 210485 175989
rect 210513 175961 210547 175989
rect 210575 175961 210609 175989
rect 210637 175961 210671 175989
rect 210699 175961 219485 175989
rect 219513 175961 219547 175989
rect 219575 175961 219609 175989
rect 219637 175961 219671 175989
rect 219699 175961 228485 175989
rect 228513 175961 228547 175989
rect 228575 175961 228609 175989
rect 228637 175961 228671 175989
rect 228699 175961 237485 175989
rect 237513 175961 237547 175989
rect 237575 175961 237609 175989
rect 237637 175961 237671 175989
rect 237699 175961 246485 175989
rect 246513 175961 246547 175989
rect 246575 175961 246609 175989
rect 246637 175961 246671 175989
rect 246699 175961 255485 175989
rect 255513 175961 255547 175989
rect 255575 175961 255609 175989
rect 255637 175961 255671 175989
rect 255699 175961 264485 175989
rect 264513 175961 264547 175989
rect 264575 175961 264609 175989
rect 264637 175961 264671 175989
rect 264699 175961 273485 175989
rect 273513 175961 273547 175989
rect 273575 175961 273609 175989
rect 273637 175961 273671 175989
rect 273699 175961 282485 175989
rect 282513 175961 282547 175989
rect 282575 175961 282609 175989
rect 282637 175961 282671 175989
rect 282699 175961 291485 175989
rect 291513 175961 291547 175989
rect 291575 175961 291609 175989
rect 291637 175961 291671 175989
rect 291699 175961 298728 175989
rect 298756 175961 298790 175989
rect 298818 175961 298852 175989
rect 298880 175961 298914 175989
rect 298942 175961 298990 175989
rect -958 175913 298990 175961
rect -958 173175 298990 173223
rect -958 173147 -430 173175
rect -402 173147 -368 173175
rect -340 173147 -306 173175
rect -278 173147 -244 173175
rect -216 173147 1625 173175
rect 1653 173147 1687 173175
rect 1715 173147 1749 173175
rect 1777 173147 1811 173175
rect 1839 173147 10625 173175
rect 10653 173147 10687 173175
rect 10715 173147 10749 173175
rect 10777 173147 10811 173175
rect 10839 173147 19625 173175
rect 19653 173147 19687 173175
rect 19715 173147 19749 173175
rect 19777 173147 19811 173175
rect 19839 173147 28625 173175
rect 28653 173147 28687 173175
rect 28715 173147 28749 173175
rect 28777 173147 28811 173175
rect 28839 173147 37625 173175
rect 37653 173147 37687 173175
rect 37715 173147 37749 173175
rect 37777 173147 37811 173175
rect 37839 173147 46625 173175
rect 46653 173147 46687 173175
rect 46715 173147 46749 173175
rect 46777 173147 46811 173175
rect 46839 173147 52259 173175
rect 52287 173147 52321 173175
rect 52349 173147 67619 173175
rect 67647 173147 67681 173175
rect 67709 173147 82979 173175
rect 83007 173147 83041 173175
rect 83069 173147 98339 173175
rect 98367 173147 98401 173175
rect 98429 173147 113699 173175
rect 113727 173147 113761 173175
rect 113789 173147 129059 173175
rect 129087 173147 129121 173175
rect 129149 173147 144419 173175
rect 144447 173147 144481 173175
rect 144509 173147 154625 173175
rect 154653 173147 154687 173175
rect 154715 173147 154749 173175
rect 154777 173147 154811 173175
rect 154839 173147 163625 173175
rect 163653 173147 163687 173175
rect 163715 173147 163749 173175
rect 163777 173147 163811 173175
rect 163839 173147 172625 173175
rect 172653 173147 172687 173175
rect 172715 173147 172749 173175
rect 172777 173147 172811 173175
rect 172839 173147 181625 173175
rect 181653 173147 181687 173175
rect 181715 173147 181749 173175
rect 181777 173147 181811 173175
rect 181839 173147 190625 173175
rect 190653 173147 190687 173175
rect 190715 173147 190749 173175
rect 190777 173147 190811 173175
rect 190839 173147 199625 173175
rect 199653 173147 199687 173175
rect 199715 173147 199749 173175
rect 199777 173147 199811 173175
rect 199839 173147 208625 173175
rect 208653 173147 208687 173175
rect 208715 173147 208749 173175
rect 208777 173147 208811 173175
rect 208839 173147 217625 173175
rect 217653 173147 217687 173175
rect 217715 173147 217749 173175
rect 217777 173147 217811 173175
rect 217839 173147 226625 173175
rect 226653 173147 226687 173175
rect 226715 173147 226749 173175
rect 226777 173147 226811 173175
rect 226839 173147 235625 173175
rect 235653 173147 235687 173175
rect 235715 173147 235749 173175
rect 235777 173147 235811 173175
rect 235839 173147 244625 173175
rect 244653 173147 244687 173175
rect 244715 173147 244749 173175
rect 244777 173147 244811 173175
rect 244839 173147 253625 173175
rect 253653 173147 253687 173175
rect 253715 173147 253749 173175
rect 253777 173147 253811 173175
rect 253839 173147 262625 173175
rect 262653 173147 262687 173175
rect 262715 173147 262749 173175
rect 262777 173147 262811 173175
rect 262839 173147 271625 173175
rect 271653 173147 271687 173175
rect 271715 173147 271749 173175
rect 271777 173147 271811 173175
rect 271839 173147 280625 173175
rect 280653 173147 280687 173175
rect 280715 173147 280749 173175
rect 280777 173147 280811 173175
rect 280839 173147 289625 173175
rect 289653 173147 289687 173175
rect 289715 173147 289749 173175
rect 289777 173147 289811 173175
rect 289839 173147 298248 173175
rect 298276 173147 298310 173175
rect 298338 173147 298372 173175
rect 298400 173147 298434 173175
rect 298462 173147 298990 173175
rect -958 173113 298990 173147
rect -958 173085 -430 173113
rect -402 173085 -368 173113
rect -340 173085 -306 173113
rect -278 173085 -244 173113
rect -216 173085 1625 173113
rect 1653 173085 1687 173113
rect 1715 173085 1749 173113
rect 1777 173085 1811 173113
rect 1839 173085 10625 173113
rect 10653 173085 10687 173113
rect 10715 173085 10749 173113
rect 10777 173085 10811 173113
rect 10839 173085 19625 173113
rect 19653 173085 19687 173113
rect 19715 173085 19749 173113
rect 19777 173085 19811 173113
rect 19839 173085 28625 173113
rect 28653 173085 28687 173113
rect 28715 173085 28749 173113
rect 28777 173085 28811 173113
rect 28839 173085 37625 173113
rect 37653 173085 37687 173113
rect 37715 173085 37749 173113
rect 37777 173085 37811 173113
rect 37839 173085 46625 173113
rect 46653 173085 46687 173113
rect 46715 173085 46749 173113
rect 46777 173085 46811 173113
rect 46839 173085 52259 173113
rect 52287 173085 52321 173113
rect 52349 173085 67619 173113
rect 67647 173085 67681 173113
rect 67709 173085 82979 173113
rect 83007 173085 83041 173113
rect 83069 173085 98339 173113
rect 98367 173085 98401 173113
rect 98429 173085 113699 173113
rect 113727 173085 113761 173113
rect 113789 173085 129059 173113
rect 129087 173085 129121 173113
rect 129149 173085 144419 173113
rect 144447 173085 144481 173113
rect 144509 173085 154625 173113
rect 154653 173085 154687 173113
rect 154715 173085 154749 173113
rect 154777 173085 154811 173113
rect 154839 173085 163625 173113
rect 163653 173085 163687 173113
rect 163715 173085 163749 173113
rect 163777 173085 163811 173113
rect 163839 173085 172625 173113
rect 172653 173085 172687 173113
rect 172715 173085 172749 173113
rect 172777 173085 172811 173113
rect 172839 173085 181625 173113
rect 181653 173085 181687 173113
rect 181715 173085 181749 173113
rect 181777 173085 181811 173113
rect 181839 173085 190625 173113
rect 190653 173085 190687 173113
rect 190715 173085 190749 173113
rect 190777 173085 190811 173113
rect 190839 173085 199625 173113
rect 199653 173085 199687 173113
rect 199715 173085 199749 173113
rect 199777 173085 199811 173113
rect 199839 173085 208625 173113
rect 208653 173085 208687 173113
rect 208715 173085 208749 173113
rect 208777 173085 208811 173113
rect 208839 173085 217625 173113
rect 217653 173085 217687 173113
rect 217715 173085 217749 173113
rect 217777 173085 217811 173113
rect 217839 173085 226625 173113
rect 226653 173085 226687 173113
rect 226715 173085 226749 173113
rect 226777 173085 226811 173113
rect 226839 173085 235625 173113
rect 235653 173085 235687 173113
rect 235715 173085 235749 173113
rect 235777 173085 235811 173113
rect 235839 173085 244625 173113
rect 244653 173085 244687 173113
rect 244715 173085 244749 173113
rect 244777 173085 244811 173113
rect 244839 173085 253625 173113
rect 253653 173085 253687 173113
rect 253715 173085 253749 173113
rect 253777 173085 253811 173113
rect 253839 173085 262625 173113
rect 262653 173085 262687 173113
rect 262715 173085 262749 173113
rect 262777 173085 262811 173113
rect 262839 173085 271625 173113
rect 271653 173085 271687 173113
rect 271715 173085 271749 173113
rect 271777 173085 271811 173113
rect 271839 173085 280625 173113
rect 280653 173085 280687 173113
rect 280715 173085 280749 173113
rect 280777 173085 280811 173113
rect 280839 173085 289625 173113
rect 289653 173085 289687 173113
rect 289715 173085 289749 173113
rect 289777 173085 289811 173113
rect 289839 173085 298248 173113
rect 298276 173085 298310 173113
rect 298338 173085 298372 173113
rect 298400 173085 298434 173113
rect 298462 173085 298990 173113
rect -958 173051 298990 173085
rect -958 173023 -430 173051
rect -402 173023 -368 173051
rect -340 173023 -306 173051
rect -278 173023 -244 173051
rect -216 173023 1625 173051
rect 1653 173023 1687 173051
rect 1715 173023 1749 173051
rect 1777 173023 1811 173051
rect 1839 173023 10625 173051
rect 10653 173023 10687 173051
rect 10715 173023 10749 173051
rect 10777 173023 10811 173051
rect 10839 173023 19625 173051
rect 19653 173023 19687 173051
rect 19715 173023 19749 173051
rect 19777 173023 19811 173051
rect 19839 173023 28625 173051
rect 28653 173023 28687 173051
rect 28715 173023 28749 173051
rect 28777 173023 28811 173051
rect 28839 173023 37625 173051
rect 37653 173023 37687 173051
rect 37715 173023 37749 173051
rect 37777 173023 37811 173051
rect 37839 173023 46625 173051
rect 46653 173023 46687 173051
rect 46715 173023 46749 173051
rect 46777 173023 46811 173051
rect 46839 173023 52259 173051
rect 52287 173023 52321 173051
rect 52349 173023 67619 173051
rect 67647 173023 67681 173051
rect 67709 173023 82979 173051
rect 83007 173023 83041 173051
rect 83069 173023 98339 173051
rect 98367 173023 98401 173051
rect 98429 173023 113699 173051
rect 113727 173023 113761 173051
rect 113789 173023 129059 173051
rect 129087 173023 129121 173051
rect 129149 173023 144419 173051
rect 144447 173023 144481 173051
rect 144509 173023 154625 173051
rect 154653 173023 154687 173051
rect 154715 173023 154749 173051
rect 154777 173023 154811 173051
rect 154839 173023 163625 173051
rect 163653 173023 163687 173051
rect 163715 173023 163749 173051
rect 163777 173023 163811 173051
rect 163839 173023 172625 173051
rect 172653 173023 172687 173051
rect 172715 173023 172749 173051
rect 172777 173023 172811 173051
rect 172839 173023 181625 173051
rect 181653 173023 181687 173051
rect 181715 173023 181749 173051
rect 181777 173023 181811 173051
rect 181839 173023 190625 173051
rect 190653 173023 190687 173051
rect 190715 173023 190749 173051
rect 190777 173023 190811 173051
rect 190839 173023 199625 173051
rect 199653 173023 199687 173051
rect 199715 173023 199749 173051
rect 199777 173023 199811 173051
rect 199839 173023 208625 173051
rect 208653 173023 208687 173051
rect 208715 173023 208749 173051
rect 208777 173023 208811 173051
rect 208839 173023 217625 173051
rect 217653 173023 217687 173051
rect 217715 173023 217749 173051
rect 217777 173023 217811 173051
rect 217839 173023 226625 173051
rect 226653 173023 226687 173051
rect 226715 173023 226749 173051
rect 226777 173023 226811 173051
rect 226839 173023 235625 173051
rect 235653 173023 235687 173051
rect 235715 173023 235749 173051
rect 235777 173023 235811 173051
rect 235839 173023 244625 173051
rect 244653 173023 244687 173051
rect 244715 173023 244749 173051
rect 244777 173023 244811 173051
rect 244839 173023 253625 173051
rect 253653 173023 253687 173051
rect 253715 173023 253749 173051
rect 253777 173023 253811 173051
rect 253839 173023 262625 173051
rect 262653 173023 262687 173051
rect 262715 173023 262749 173051
rect 262777 173023 262811 173051
rect 262839 173023 271625 173051
rect 271653 173023 271687 173051
rect 271715 173023 271749 173051
rect 271777 173023 271811 173051
rect 271839 173023 280625 173051
rect 280653 173023 280687 173051
rect 280715 173023 280749 173051
rect 280777 173023 280811 173051
rect 280839 173023 289625 173051
rect 289653 173023 289687 173051
rect 289715 173023 289749 173051
rect 289777 173023 289811 173051
rect 289839 173023 298248 173051
rect 298276 173023 298310 173051
rect 298338 173023 298372 173051
rect 298400 173023 298434 173051
rect 298462 173023 298990 173051
rect -958 172989 298990 173023
rect -958 172961 -430 172989
rect -402 172961 -368 172989
rect -340 172961 -306 172989
rect -278 172961 -244 172989
rect -216 172961 1625 172989
rect 1653 172961 1687 172989
rect 1715 172961 1749 172989
rect 1777 172961 1811 172989
rect 1839 172961 10625 172989
rect 10653 172961 10687 172989
rect 10715 172961 10749 172989
rect 10777 172961 10811 172989
rect 10839 172961 19625 172989
rect 19653 172961 19687 172989
rect 19715 172961 19749 172989
rect 19777 172961 19811 172989
rect 19839 172961 28625 172989
rect 28653 172961 28687 172989
rect 28715 172961 28749 172989
rect 28777 172961 28811 172989
rect 28839 172961 37625 172989
rect 37653 172961 37687 172989
rect 37715 172961 37749 172989
rect 37777 172961 37811 172989
rect 37839 172961 46625 172989
rect 46653 172961 46687 172989
rect 46715 172961 46749 172989
rect 46777 172961 46811 172989
rect 46839 172961 52259 172989
rect 52287 172961 52321 172989
rect 52349 172961 67619 172989
rect 67647 172961 67681 172989
rect 67709 172961 82979 172989
rect 83007 172961 83041 172989
rect 83069 172961 98339 172989
rect 98367 172961 98401 172989
rect 98429 172961 113699 172989
rect 113727 172961 113761 172989
rect 113789 172961 129059 172989
rect 129087 172961 129121 172989
rect 129149 172961 144419 172989
rect 144447 172961 144481 172989
rect 144509 172961 154625 172989
rect 154653 172961 154687 172989
rect 154715 172961 154749 172989
rect 154777 172961 154811 172989
rect 154839 172961 163625 172989
rect 163653 172961 163687 172989
rect 163715 172961 163749 172989
rect 163777 172961 163811 172989
rect 163839 172961 172625 172989
rect 172653 172961 172687 172989
rect 172715 172961 172749 172989
rect 172777 172961 172811 172989
rect 172839 172961 181625 172989
rect 181653 172961 181687 172989
rect 181715 172961 181749 172989
rect 181777 172961 181811 172989
rect 181839 172961 190625 172989
rect 190653 172961 190687 172989
rect 190715 172961 190749 172989
rect 190777 172961 190811 172989
rect 190839 172961 199625 172989
rect 199653 172961 199687 172989
rect 199715 172961 199749 172989
rect 199777 172961 199811 172989
rect 199839 172961 208625 172989
rect 208653 172961 208687 172989
rect 208715 172961 208749 172989
rect 208777 172961 208811 172989
rect 208839 172961 217625 172989
rect 217653 172961 217687 172989
rect 217715 172961 217749 172989
rect 217777 172961 217811 172989
rect 217839 172961 226625 172989
rect 226653 172961 226687 172989
rect 226715 172961 226749 172989
rect 226777 172961 226811 172989
rect 226839 172961 235625 172989
rect 235653 172961 235687 172989
rect 235715 172961 235749 172989
rect 235777 172961 235811 172989
rect 235839 172961 244625 172989
rect 244653 172961 244687 172989
rect 244715 172961 244749 172989
rect 244777 172961 244811 172989
rect 244839 172961 253625 172989
rect 253653 172961 253687 172989
rect 253715 172961 253749 172989
rect 253777 172961 253811 172989
rect 253839 172961 262625 172989
rect 262653 172961 262687 172989
rect 262715 172961 262749 172989
rect 262777 172961 262811 172989
rect 262839 172961 271625 172989
rect 271653 172961 271687 172989
rect 271715 172961 271749 172989
rect 271777 172961 271811 172989
rect 271839 172961 280625 172989
rect 280653 172961 280687 172989
rect 280715 172961 280749 172989
rect 280777 172961 280811 172989
rect 280839 172961 289625 172989
rect 289653 172961 289687 172989
rect 289715 172961 289749 172989
rect 289777 172961 289811 172989
rect 289839 172961 298248 172989
rect 298276 172961 298310 172989
rect 298338 172961 298372 172989
rect 298400 172961 298434 172989
rect 298462 172961 298990 172989
rect -958 172913 298990 172961
rect -958 167175 298990 167223
rect -958 167147 -910 167175
rect -882 167147 -848 167175
rect -820 167147 -786 167175
rect -758 167147 -724 167175
rect -696 167147 3485 167175
rect 3513 167147 3547 167175
rect 3575 167147 3609 167175
rect 3637 167147 3671 167175
rect 3699 167147 12485 167175
rect 12513 167147 12547 167175
rect 12575 167147 12609 167175
rect 12637 167147 12671 167175
rect 12699 167147 21485 167175
rect 21513 167147 21547 167175
rect 21575 167147 21609 167175
rect 21637 167147 21671 167175
rect 21699 167147 30485 167175
rect 30513 167147 30547 167175
rect 30575 167147 30609 167175
rect 30637 167147 30671 167175
rect 30699 167147 39485 167175
rect 39513 167147 39547 167175
rect 39575 167147 39609 167175
rect 39637 167147 39671 167175
rect 39699 167147 48485 167175
rect 48513 167147 48547 167175
rect 48575 167147 48609 167175
rect 48637 167147 48671 167175
rect 48699 167147 59939 167175
rect 59967 167147 60001 167175
rect 60029 167147 75299 167175
rect 75327 167147 75361 167175
rect 75389 167147 90659 167175
rect 90687 167147 90721 167175
rect 90749 167147 106019 167175
rect 106047 167147 106081 167175
rect 106109 167147 121379 167175
rect 121407 167147 121441 167175
rect 121469 167147 136739 167175
rect 136767 167147 136801 167175
rect 136829 167147 156485 167175
rect 156513 167147 156547 167175
rect 156575 167147 156609 167175
rect 156637 167147 156671 167175
rect 156699 167147 165485 167175
rect 165513 167147 165547 167175
rect 165575 167147 165609 167175
rect 165637 167147 165671 167175
rect 165699 167147 174485 167175
rect 174513 167147 174547 167175
rect 174575 167147 174609 167175
rect 174637 167147 174671 167175
rect 174699 167147 183485 167175
rect 183513 167147 183547 167175
rect 183575 167147 183609 167175
rect 183637 167147 183671 167175
rect 183699 167147 192485 167175
rect 192513 167147 192547 167175
rect 192575 167147 192609 167175
rect 192637 167147 192671 167175
rect 192699 167147 201485 167175
rect 201513 167147 201547 167175
rect 201575 167147 201609 167175
rect 201637 167147 201671 167175
rect 201699 167147 210485 167175
rect 210513 167147 210547 167175
rect 210575 167147 210609 167175
rect 210637 167147 210671 167175
rect 210699 167147 219485 167175
rect 219513 167147 219547 167175
rect 219575 167147 219609 167175
rect 219637 167147 219671 167175
rect 219699 167147 228485 167175
rect 228513 167147 228547 167175
rect 228575 167147 228609 167175
rect 228637 167147 228671 167175
rect 228699 167147 237485 167175
rect 237513 167147 237547 167175
rect 237575 167147 237609 167175
rect 237637 167147 237671 167175
rect 237699 167147 246485 167175
rect 246513 167147 246547 167175
rect 246575 167147 246609 167175
rect 246637 167147 246671 167175
rect 246699 167147 255485 167175
rect 255513 167147 255547 167175
rect 255575 167147 255609 167175
rect 255637 167147 255671 167175
rect 255699 167147 264485 167175
rect 264513 167147 264547 167175
rect 264575 167147 264609 167175
rect 264637 167147 264671 167175
rect 264699 167147 273485 167175
rect 273513 167147 273547 167175
rect 273575 167147 273609 167175
rect 273637 167147 273671 167175
rect 273699 167147 282485 167175
rect 282513 167147 282547 167175
rect 282575 167147 282609 167175
rect 282637 167147 282671 167175
rect 282699 167147 291485 167175
rect 291513 167147 291547 167175
rect 291575 167147 291609 167175
rect 291637 167147 291671 167175
rect 291699 167147 298728 167175
rect 298756 167147 298790 167175
rect 298818 167147 298852 167175
rect 298880 167147 298914 167175
rect 298942 167147 298990 167175
rect -958 167113 298990 167147
rect -958 167085 -910 167113
rect -882 167085 -848 167113
rect -820 167085 -786 167113
rect -758 167085 -724 167113
rect -696 167085 3485 167113
rect 3513 167085 3547 167113
rect 3575 167085 3609 167113
rect 3637 167085 3671 167113
rect 3699 167085 12485 167113
rect 12513 167085 12547 167113
rect 12575 167085 12609 167113
rect 12637 167085 12671 167113
rect 12699 167085 21485 167113
rect 21513 167085 21547 167113
rect 21575 167085 21609 167113
rect 21637 167085 21671 167113
rect 21699 167085 30485 167113
rect 30513 167085 30547 167113
rect 30575 167085 30609 167113
rect 30637 167085 30671 167113
rect 30699 167085 39485 167113
rect 39513 167085 39547 167113
rect 39575 167085 39609 167113
rect 39637 167085 39671 167113
rect 39699 167085 48485 167113
rect 48513 167085 48547 167113
rect 48575 167085 48609 167113
rect 48637 167085 48671 167113
rect 48699 167085 59939 167113
rect 59967 167085 60001 167113
rect 60029 167085 75299 167113
rect 75327 167085 75361 167113
rect 75389 167085 90659 167113
rect 90687 167085 90721 167113
rect 90749 167085 106019 167113
rect 106047 167085 106081 167113
rect 106109 167085 121379 167113
rect 121407 167085 121441 167113
rect 121469 167085 136739 167113
rect 136767 167085 136801 167113
rect 136829 167085 156485 167113
rect 156513 167085 156547 167113
rect 156575 167085 156609 167113
rect 156637 167085 156671 167113
rect 156699 167085 165485 167113
rect 165513 167085 165547 167113
rect 165575 167085 165609 167113
rect 165637 167085 165671 167113
rect 165699 167085 174485 167113
rect 174513 167085 174547 167113
rect 174575 167085 174609 167113
rect 174637 167085 174671 167113
rect 174699 167085 183485 167113
rect 183513 167085 183547 167113
rect 183575 167085 183609 167113
rect 183637 167085 183671 167113
rect 183699 167085 192485 167113
rect 192513 167085 192547 167113
rect 192575 167085 192609 167113
rect 192637 167085 192671 167113
rect 192699 167085 201485 167113
rect 201513 167085 201547 167113
rect 201575 167085 201609 167113
rect 201637 167085 201671 167113
rect 201699 167085 210485 167113
rect 210513 167085 210547 167113
rect 210575 167085 210609 167113
rect 210637 167085 210671 167113
rect 210699 167085 219485 167113
rect 219513 167085 219547 167113
rect 219575 167085 219609 167113
rect 219637 167085 219671 167113
rect 219699 167085 228485 167113
rect 228513 167085 228547 167113
rect 228575 167085 228609 167113
rect 228637 167085 228671 167113
rect 228699 167085 237485 167113
rect 237513 167085 237547 167113
rect 237575 167085 237609 167113
rect 237637 167085 237671 167113
rect 237699 167085 246485 167113
rect 246513 167085 246547 167113
rect 246575 167085 246609 167113
rect 246637 167085 246671 167113
rect 246699 167085 255485 167113
rect 255513 167085 255547 167113
rect 255575 167085 255609 167113
rect 255637 167085 255671 167113
rect 255699 167085 264485 167113
rect 264513 167085 264547 167113
rect 264575 167085 264609 167113
rect 264637 167085 264671 167113
rect 264699 167085 273485 167113
rect 273513 167085 273547 167113
rect 273575 167085 273609 167113
rect 273637 167085 273671 167113
rect 273699 167085 282485 167113
rect 282513 167085 282547 167113
rect 282575 167085 282609 167113
rect 282637 167085 282671 167113
rect 282699 167085 291485 167113
rect 291513 167085 291547 167113
rect 291575 167085 291609 167113
rect 291637 167085 291671 167113
rect 291699 167085 298728 167113
rect 298756 167085 298790 167113
rect 298818 167085 298852 167113
rect 298880 167085 298914 167113
rect 298942 167085 298990 167113
rect -958 167051 298990 167085
rect -958 167023 -910 167051
rect -882 167023 -848 167051
rect -820 167023 -786 167051
rect -758 167023 -724 167051
rect -696 167023 3485 167051
rect 3513 167023 3547 167051
rect 3575 167023 3609 167051
rect 3637 167023 3671 167051
rect 3699 167023 12485 167051
rect 12513 167023 12547 167051
rect 12575 167023 12609 167051
rect 12637 167023 12671 167051
rect 12699 167023 21485 167051
rect 21513 167023 21547 167051
rect 21575 167023 21609 167051
rect 21637 167023 21671 167051
rect 21699 167023 30485 167051
rect 30513 167023 30547 167051
rect 30575 167023 30609 167051
rect 30637 167023 30671 167051
rect 30699 167023 39485 167051
rect 39513 167023 39547 167051
rect 39575 167023 39609 167051
rect 39637 167023 39671 167051
rect 39699 167023 48485 167051
rect 48513 167023 48547 167051
rect 48575 167023 48609 167051
rect 48637 167023 48671 167051
rect 48699 167023 59939 167051
rect 59967 167023 60001 167051
rect 60029 167023 75299 167051
rect 75327 167023 75361 167051
rect 75389 167023 90659 167051
rect 90687 167023 90721 167051
rect 90749 167023 106019 167051
rect 106047 167023 106081 167051
rect 106109 167023 121379 167051
rect 121407 167023 121441 167051
rect 121469 167023 136739 167051
rect 136767 167023 136801 167051
rect 136829 167023 156485 167051
rect 156513 167023 156547 167051
rect 156575 167023 156609 167051
rect 156637 167023 156671 167051
rect 156699 167023 165485 167051
rect 165513 167023 165547 167051
rect 165575 167023 165609 167051
rect 165637 167023 165671 167051
rect 165699 167023 174485 167051
rect 174513 167023 174547 167051
rect 174575 167023 174609 167051
rect 174637 167023 174671 167051
rect 174699 167023 183485 167051
rect 183513 167023 183547 167051
rect 183575 167023 183609 167051
rect 183637 167023 183671 167051
rect 183699 167023 192485 167051
rect 192513 167023 192547 167051
rect 192575 167023 192609 167051
rect 192637 167023 192671 167051
rect 192699 167023 201485 167051
rect 201513 167023 201547 167051
rect 201575 167023 201609 167051
rect 201637 167023 201671 167051
rect 201699 167023 210485 167051
rect 210513 167023 210547 167051
rect 210575 167023 210609 167051
rect 210637 167023 210671 167051
rect 210699 167023 219485 167051
rect 219513 167023 219547 167051
rect 219575 167023 219609 167051
rect 219637 167023 219671 167051
rect 219699 167023 228485 167051
rect 228513 167023 228547 167051
rect 228575 167023 228609 167051
rect 228637 167023 228671 167051
rect 228699 167023 237485 167051
rect 237513 167023 237547 167051
rect 237575 167023 237609 167051
rect 237637 167023 237671 167051
rect 237699 167023 246485 167051
rect 246513 167023 246547 167051
rect 246575 167023 246609 167051
rect 246637 167023 246671 167051
rect 246699 167023 255485 167051
rect 255513 167023 255547 167051
rect 255575 167023 255609 167051
rect 255637 167023 255671 167051
rect 255699 167023 264485 167051
rect 264513 167023 264547 167051
rect 264575 167023 264609 167051
rect 264637 167023 264671 167051
rect 264699 167023 273485 167051
rect 273513 167023 273547 167051
rect 273575 167023 273609 167051
rect 273637 167023 273671 167051
rect 273699 167023 282485 167051
rect 282513 167023 282547 167051
rect 282575 167023 282609 167051
rect 282637 167023 282671 167051
rect 282699 167023 291485 167051
rect 291513 167023 291547 167051
rect 291575 167023 291609 167051
rect 291637 167023 291671 167051
rect 291699 167023 298728 167051
rect 298756 167023 298790 167051
rect 298818 167023 298852 167051
rect 298880 167023 298914 167051
rect 298942 167023 298990 167051
rect -958 166989 298990 167023
rect -958 166961 -910 166989
rect -882 166961 -848 166989
rect -820 166961 -786 166989
rect -758 166961 -724 166989
rect -696 166961 3485 166989
rect 3513 166961 3547 166989
rect 3575 166961 3609 166989
rect 3637 166961 3671 166989
rect 3699 166961 12485 166989
rect 12513 166961 12547 166989
rect 12575 166961 12609 166989
rect 12637 166961 12671 166989
rect 12699 166961 21485 166989
rect 21513 166961 21547 166989
rect 21575 166961 21609 166989
rect 21637 166961 21671 166989
rect 21699 166961 30485 166989
rect 30513 166961 30547 166989
rect 30575 166961 30609 166989
rect 30637 166961 30671 166989
rect 30699 166961 39485 166989
rect 39513 166961 39547 166989
rect 39575 166961 39609 166989
rect 39637 166961 39671 166989
rect 39699 166961 48485 166989
rect 48513 166961 48547 166989
rect 48575 166961 48609 166989
rect 48637 166961 48671 166989
rect 48699 166961 59939 166989
rect 59967 166961 60001 166989
rect 60029 166961 75299 166989
rect 75327 166961 75361 166989
rect 75389 166961 90659 166989
rect 90687 166961 90721 166989
rect 90749 166961 106019 166989
rect 106047 166961 106081 166989
rect 106109 166961 121379 166989
rect 121407 166961 121441 166989
rect 121469 166961 136739 166989
rect 136767 166961 136801 166989
rect 136829 166961 156485 166989
rect 156513 166961 156547 166989
rect 156575 166961 156609 166989
rect 156637 166961 156671 166989
rect 156699 166961 165485 166989
rect 165513 166961 165547 166989
rect 165575 166961 165609 166989
rect 165637 166961 165671 166989
rect 165699 166961 174485 166989
rect 174513 166961 174547 166989
rect 174575 166961 174609 166989
rect 174637 166961 174671 166989
rect 174699 166961 183485 166989
rect 183513 166961 183547 166989
rect 183575 166961 183609 166989
rect 183637 166961 183671 166989
rect 183699 166961 192485 166989
rect 192513 166961 192547 166989
rect 192575 166961 192609 166989
rect 192637 166961 192671 166989
rect 192699 166961 201485 166989
rect 201513 166961 201547 166989
rect 201575 166961 201609 166989
rect 201637 166961 201671 166989
rect 201699 166961 210485 166989
rect 210513 166961 210547 166989
rect 210575 166961 210609 166989
rect 210637 166961 210671 166989
rect 210699 166961 219485 166989
rect 219513 166961 219547 166989
rect 219575 166961 219609 166989
rect 219637 166961 219671 166989
rect 219699 166961 228485 166989
rect 228513 166961 228547 166989
rect 228575 166961 228609 166989
rect 228637 166961 228671 166989
rect 228699 166961 237485 166989
rect 237513 166961 237547 166989
rect 237575 166961 237609 166989
rect 237637 166961 237671 166989
rect 237699 166961 246485 166989
rect 246513 166961 246547 166989
rect 246575 166961 246609 166989
rect 246637 166961 246671 166989
rect 246699 166961 255485 166989
rect 255513 166961 255547 166989
rect 255575 166961 255609 166989
rect 255637 166961 255671 166989
rect 255699 166961 264485 166989
rect 264513 166961 264547 166989
rect 264575 166961 264609 166989
rect 264637 166961 264671 166989
rect 264699 166961 273485 166989
rect 273513 166961 273547 166989
rect 273575 166961 273609 166989
rect 273637 166961 273671 166989
rect 273699 166961 282485 166989
rect 282513 166961 282547 166989
rect 282575 166961 282609 166989
rect 282637 166961 282671 166989
rect 282699 166961 291485 166989
rect 291513 166961 291547 166989
rect 291575 166961 291609 166989
rect 291637 166961 291671 166989
rect 291699 166961 298728 166989
rect 298756 166961 298790 166989
rect 298818 166961 298852 166989
rect 298880 166961 298914 166989
rect 298942 166961 298990 166989
rect -958 166913 298990 166961
rect -958 164175 298990 164223
rect -958 164147 -430 164175
rect -402 164147 -368 164175
rect -340 164147 -306 164175
rect -278 164147 -244 164175
rect -216 164147 1625 164175
rect 1653 164147 1687 164175
rect 1715 164147 1749 164175
rect 1777 164147 1811 164175
rect 1839 164147 10625 164175
rect 10653 164147 10687 164175
rect 10715 164147 10749 164175
rect 10777 164147 10811 164175
rect 10839 164147 19625 164175
rect 19653 164147 19687 164175
rect 19715 164147 19749 164175
rect 19777 164147 19811 164175
rect 19839 164147 28625 164175
rect 28653 164147 28687 164175
rect 28715 164147 28749 164175
rect 28777 164147 28811 164175
rect 28839 164147 37625 164175
rect 37653 164147 37687 164175
rect 37715 164147 37749 164175
rect 37777 164147 37811 164175
rect 37839 164147 46625 164175
rect 46653 164147 46687 164175
rect 46715 164147 46749 164175
rect 46777 164147 46811 164175
rect 46839 164147 52259 164175
rect 52287 164147 52321 164175
rect 52349 164147 67619 164175
rect 67647 164147 67681 164175
rect 67709 164147 82979 164175
rect 83007 164147 83041 164175
rect 83069 164147 98339 164175
rect 98367 164147 98401 164175
rect 98429 164147 113699 164175
rect 113727 164147 113761 164175
rect 113789 164147 129059 164175
rect 129087 164147 129121 164175
rect 129149 164147 144419 164175
rect 144447 164147 144481 164175
rect 144509 164147 154625 164175
rect 154653 164147 154687 164175
rect 154715 164147 154749 164175
rect 154777 164147 154811 164175
rect 154839 164147 163625 164175
rect 163653 164147 163687 164175
rect 163715 164147 163749 164175
rect 163777 164147 163811 164175
rect 163839 164147 172625 164175
rect 172653 164147 172687 164175
rect 172715 164147 172749 164175
rect 172777 164147 172811 164175
rect 172839 164147 181625 164175
rect 181653 164147 181687 164175
rect 181715 164147 181749 164175
rect 181777 164147 181811 164175
rect 181839 164147 190625 164175
rect 190653 164147 190687 164175
rect 190715 164147 190749 164175
rect 190777 164147 190811 164175
rect 190839 164147 199625 164175
rect 199653 164147 199687 164175
rect 199715 164147 199749 164175
rect 199777 164147 199811 164175
rect 199839 164147 208625 164175
rect 208653 164147 208687 164175
rect 208715 164147 208749 164175
rect 208777 164147 208811 164175
rect 208839 164147 217625 164175
rect 217653 164147 217687 164175
rect 217715 164147 217749 164175
rect 217777 164147 217811 164175
rect 217839 164147 226625 164175
rect 226653 164147 226687 164175
rect 226715 164147 226749 164175
rect 226777 164147 226811 164175
rect 226839 164147 235625 164175
rect 235653 164147 235687 164175
rect 235715 164147 235749 164175
rect 235777 164147 235811 164175
rect 235839 164147 244625 164175
rect 244653 164147 244687 164175
rect 244715 164147 244749 164175
rect 244777 164147 244811 164175
rect 244839 164147 253625 164175
rect 253653 164147 253687 164175
rect 253715 164147 253749 164175
rect 253777 164147 253811 164175
rect 253839 164147 262625 164175
rect 262653 164147 262687 164175
rect 262715 164147 262749 164175
rect 262777 164147 262811 164175
rect 262839 164147 271625 164175
rect 271653 164147 271687 164175
rect 271715 164147 271749 164175
rect 271777 164147 271811 164175
rect 271839 164147 280625 164175
rect 280653 164147 280687 164175
rect 280715 164147 280749 164175
rect 280777 164147 280811 164175
rect 280839 164147 289625 164175
rect 289653 164147 289687 164175
rect 289715 164147 289749 164175
rect 289777 164147 289811 164175
rect 289839 164147 298248 164175
rect 298276 164147 298310 164175
rect 298338 164147 298372 164175
rect 298400 164147 298434 164175
rect 298462 164147 298990 164175
rect -958 164113 298990 164147
rect -958 164085 -430 164113
rect -402 164085 -368 164113
rect -340 164085 -306 164113
rect -278 164085 -244 164113
rect -216 164085 1625 164113
rect 1653 164085 1687 164113
rect 1715 164085 1749 164113
rect 1777 164085 1811 164113
rect 1839 164085 10625 164113
rect 10653 164085 10687 164113
rect 10715 164085 10749 164113
rect 10777 164085 10811 164113
rect 10839 164085 19625 164113
rect 19653 164085 19687 164113
rect 19715 164085 19749 164113
rect 19777 164085 19811 164113
rect 19839 164085 28625 164113
rect 28653 164085 28687 164113
rect 28715 164085 28749 164113
rect 28777 164085 28811 164113
rect 28839 164085 37625 164113
rect 37653 164085 37687 164113
rect 37715 164085 37749 164113
rect 37777 164085 37811 164113
rect 37839 164085 46625 164113
rect 46653 164085 46687 164113
rect 46715 164085 46749 164113
rect 46777 164085 46811 164113
rect 46839 164085 52259 164113
rect 52287 164085 52321 164113
rect 52349 164085 67619 164113
rect 67647 164085 67681 164113
rect 67709 164085 82979 164113
rect 83007 164085 83041 164113
rect 83069 164085 98339 164113
rect 98367 164085 98401 164113
rect 98429 164085 113699 164113
rect 113727 164085 113761 164113
rect 113789 164085 129059 164113
rect 129087 164085 129121 164113
rect 129149 164085 144419 164113
rect 144447 164085 144481 164113
rect 144509 164085 154625 164113
rect 154653 164085 154687 164113
rect 154715 164085 154749 164113
rect 154777 164085 154811 164113
rect 154839 164085 163625 164113
rect 163653 164085 163687 164113
rect 163715 164085 163749 164113
rect 163777 164085 163811 164113
rect 163839 164085 172625 164113
rect 172653 164085 172687 164113
rect 172715 164085 172749 164113
rect 172777 164085 172811 164113
rect 172839 164085 181625 164113
rect 181653 164085 181687 164113
rect 181715 164085 181749 164113
rect 181777 164085 181811 164113
rect 181839 164085 190625 164113
rect 190653 164085 190687 164113
rect 190715 164085 190749 164113
rect 190777 164085 190811 164113
rect 190839 164085 199625 164113
rect 199653 164085 199687 164113
rect 199715 164085 199749 164113
rect 199777 164085 199811 164113
rect 199839 164085 208625 164113
rect 208653 164085 208687 164113
rect 208715 164085 208749 164113
rect 208777 164085 208811 164113
rect 208839 164085 217625 164113
rect 217653 164085 217687 164113
rect 217715 164085 217749 164113
rect 217777 164085 217811 164113
rect 217839 164085 226625 164113
rect 226653 164085 226687 164113
rect 226715 164085 226749 164113
rect 226777 164085 226811 164113
rect 226839 164085 235625 164113
rect 235653 164085 235687 164113
rect 235715 164085 235749 164113
rect 235777 164085 235811 164113
rect 235839 164085 244625 164113
rect 244653 164085 244687 164113
rect 244715 164085 244749 164113
rect 244777 164085 244811 164113
rect 244839 164085 253625 164113
rect 253653 164085 253687 164113
rect 253715 164085 253749 164113
rect 253777 164085 253811 164113
rect 253839 164085 262625 164113
rect 262653 164085 262687 164113
rect 262715 164085 262749 164113
rect 262777 164085 262811 164113
rect 262839 164085 271625 164113
rect 271653 164085 271687 164113
rect 271715 164085 271749 164113
rect 271777 164085 271811 164113
rect 271839 164085 280625 164113
rect 280653 164085 280687 164113
rect 280715 164085 280749 164113
rect 280777 164085 280811 164113
rect 280839 164085 289625 164113
rect 289653 164085 289687 164113
rect 289715 164085 289749 164113
rect 289777 164085 289811 164113
rect 289839 164085 298248 164113
rect 298276 164085 298310 164113
rect 298338 164085 298372 164113
rect 298400 164085 298434 164113
rect 298462 164085 298990 164113
rect -958 164051 298990 164085
rect -958 164023 -430 164051
rect -402 164023 -368 164051
rect -340 164023 -306 164051
rect -278 164023 -244 164051
rect -216 164023 1625 164051
rect 1653 164023 1687 164051
rect 1715 164023 1749 164051
rect 1777 164023 1811 164051
rect 1839 164023 10625 164051
rect 10653 164023 10687 164051
rect 10715 164023 10749 164051
rect 10777 164023 10811 164051
rect 10839 164023 19625 164051
rect 19653 164023 19687 164051
rect 19715 164023 19749 164051
rect 19777 164023 19811 164051
rect 19839 164023 28625 164051
rect 28653 164023 28687 164051
rect 28715 164023 28749 164051
rect 28777 164023 28811 164051
rect 28839 164023 37625 164051
rect 37653 164023 37687 164051
rect 37715 164023 37749 164051
rect 37777 164023 37811 164051
rect 37839 164023 46625 164051
rect 46653 164023 46687 164051
rect 46715 164023 46749 164051
rect 46777 164023 46811 164051
rect 46839 164023 52259 164051
rect 52287 164023 52321 164051
rect 52349 164023 67619 164051
rect 67647 164023 67681 164051
rect 67709 164023 82979 164051
rect 83007 164023 83041 164051
rect 83069 164023 98339 164051
rect 98367 164023 98401 164051
rect 98429 164023 113699 164051
rect 113727 164023 113761 164051
rect 113789 164023 129059 164051
rect 129087 164023 129121 164051
rect 129149 164023 144419 164051
rect 144447 164023 144481 164051
rect 144509 164023 154625 164051
rect 154653 164023 154687 164051
rect 154715 164023 154749 164051
rect 154777 164023 154811 164051
rect 154839 164023 163625 164051
rect 163653 164023 163687 164051
rect 163715 164023 163749 164051
rect 163777 164023 163811 164051
rect 163839 164023 172625 164051
rect 172653 164023 172687 164051
rect 172715 164023 172749 164051
rect 172777 164023 172811 164051
rect 172839 164023 181625 164051
rect 181653 164023 181687 164051
rect 181715 164023 181749 164051
rect 181777 164023 181811 164051
rect 181839 164023 190625 164051
rect 190653 164023 190687 164051
rect 190715 164023 190749 164051
rect 190777 164023 190811 164051
rect 190839 164023 199625 164051
rect 199653 164023 199687 164051
rect 199715 164023 199749 164051
rect 199777 164023 199811 164051
rect 199839 164023 208625 164051
rect 208653 164023 208687 164051
rect 208715 164023 208749 164051
rect 208777 164023 208811 164051
rect 208839 164023 217625 164051
rect 217653 164023 217687 164051
rect 217715 164023 217749 164051
rect 217777 164023 217811 164051
rect 217839 164023 226625 164051
rect 226653 164023 226687 164051
rect 226715 164023 226749 164051
rect 226777 164023 226811 164051
rect 226839 164023 235625 164051
rect 235653 164023 235687 164051
rect 235715 164023 235749 164051
rect 235777 164023 235811 164051
rect 235839 164023 244625 164051
rect 244653 164023 244687 164051
rect 244715 164023 244749 164051
rect 244777 164023 244811 164051
rect 244839 164023 253625 164051
rect 253653 164023 253687 164051
rect 253715 164023 253749 164051
rect 253777 164023 253811 164051
rect 253839 164023 262625 164051
rect 262653 164023 262687 164051
rect 262715 164023 262749 164051
rect 262777 164023 262811 164051
rect 262839 164023 271625 164051
rect 271653 164023 271687 164051
rect 271715 164023 271749 164051
rect 271777 164023 271811 164051
rect 271839 164023 280625 164051
rect 280653 164023 280687 164051
rect 280715 164023 280749 164051
rect 280777 164023 280811 164051
rect 280839 164023 289625 164051
rect 289653 164023 289687 164051
rect 289715 164023 289749 164051
rect 289777 164023 289811 164051
rect 289839 164023 298248 164051
rect 298276 164023 298310 164051
rect 298338 164023 298372 164051
rect 298400 164023 298434 164051
rect 298462 164023 298990 164051
rect -958 163989 298990 164023
rect -958 163961 -430 163989
rect -402 163961 -368 163989
rect -340 163961 -306 163989
rect -278 163961 -244 163989
rect -216 163961 1625 163989
rect 1653 163961 1687 163989
rect 1715 163961 1749 163989
rect 1777 163961 1811 163989
rect 1839 163961 10625 163989
rect 10653 163961 10687 163989
rect 10715 163961 10749 163989
rect 10777 163961 10811 163989
rect 10839 163961 19625 163989
rect 19653 163961 19687 163989
rect 19715 163961 19749 163989
rect 19777 163961 19811 163989
rect 19839 163961 28625 163989
rect 28653 163961 28687 163989
rect 28715 163961 28749 163989
rect 28777 163961 28811 163989
rect 28839 163961 37625 163989
rect 37653 163961 37687 163989
rect 37715 163961 37749 163989
rect 37777 163961 37811 163989
rect 37839 163961 46625 163989
rect 46653 163961 46687 163989
rect 46715 163961 46749 163989
rect 46777 163961 46811 163989
rect 46839 163961 52259 163989
rect 52287 163961 52321 163989
rect 52349 163961 67619 163989
rect 67647 163961 67681 163989
rect 67709 163961 82979 163989
rect 83007 163961 83041 163989
rect 83069 163961 98339 163989
rect 98367 163961 98401 163989
rect 98429 163961 113699 163989
rect 113727 163961 113761 163989
rect 113789 163961 129059 163989
rect 129087 163961 129121 163989
rect 129149 163961 144419 163989
rect 144447 163961 144481 163989
rect 144509 163961 154625 163989
rect 154653 163961 154687 163989
rect 154715 163961 154749 163989
rect 154777 163961 154811 163989
rect 154839 163961 163625 163989
rect 163653 163961 163687 163989
rect 163715 163961 163749 163989
rect 163777 163961 163811 163989
rect 163839 163961 172625 163989
rect 172653 163961 172687 163989
rect 172715 163961 172749 163989
rect 172777 163961 172811 163989
rect 172839 163961 181625 163989
rect 181653 163961 181687 163989
rect 181715 163961 181749 163989
rect 181777 163961 181811 163989
rect 181839 163961 190625 163989
rect 190653 163961 190687 163989
rect 190715 163961 190749 163989
rect 190777 163961 190811 163989
rect 190839 163961 199625 163989
rect 199653 163961 199687 163989
rect 199715 163961 199749 163989
rect 199777 163961 199811 163989
rect 199839 163961 208625 163989
rect 208653 163961 208687 163989
rect 208715 163961 208749 163989
rect 208777 163961 208811 163989
rect 208839 163961 217625 163989
rect 217653 163961 217687 163989
rect 217715 163961 217749 163989
rect 217777 163961 217811 163989
rect 217839 163961 226625 163989
rect 226653 163961 226687 163989
rect 226715 163961 226749 163989
rect 226777 163961 226811 163989
rect 226839 163961 235625 163989
rect 235653 163961 235687 163989
rect 235715 163961 235749 163989
rect 235777 163961 235811 163989
rect 235839 163961 244625 163989
rect 244653 163961 244687 163989
rect 244715 163961 244749 163989
rect 244777 163961 244811 163989
rect 244839 163961 253625 163989
rect 253653 163961 253687 163989
rect 253715 163961 253749 163989
rect 253777 163961 253811 163989
rect 253839 163961 262625 163989
rect 262653 163961 262687 163989
rect 262715 163961 262749 163989
rect 262777 163961 262811 163989
rect 262839 163961 271625 163989
rect 271653 163961 271687 163989
rect 271715 163961 271749 163989
rect 271777 163961 271811 163989
rect 271839 163961 280625 163989
rect 280653 163961 280687 163989
rect 280715 163961 280749 163989
rect 280777 163961 280811 163989
rect 280839 163961 289625 163989
rect 289653 163961 289687 163989
rect 289715 163961 289749 163989
rect 289777 163961 289811 163989
rect 289839 163961 298248 163989
rect 298276 163961 298310 163989
rect 298338 163961 298372 163989
rect 298400 163961 298434 163989
rect 298462 163961 298990 163989
rect -958 163913 298990 163961
rect -958 158175 298990 158223
rect -958 158147 -910 158175
rect -882 158147 -848 158175
rect -820 158147 -786 158175
rect -758 158147 -724 158175
rect -696 158147 3485 158175
rect 3513 158147 3547 158175
rect 3575 158147 3609 158175
rect 3637 158147 3671 158175
rect 3699 158147 12485 158175
rect 12513 158147 12547 158175
rect 12575 158147 12609 158175
rect 12637 158147 12671 158175
rect 12699 158147 21485 158175
rect 21513 158147 21547 158175
rect 21575 158147 21609 158175
rect 21637 158147 21671 158175
rect 21699 158147 30485 158175
rect 30513 158147 30547 158175
rect 30575 158147 30609 158175
rect 30637 158147 30671 158175
rect 30699 158147 39485 158175
rect 39513 158147 39547 158175
rect 39575 158147 39609 158175
rect 39637 158147 39671 158175
rect 39699 158147 48485 158175
rect 48513 158147 48547 158175
rect 48575 158147 48609 158175
rect 48637 158147 48671 158175
rect 48699 158147 59939 158175
rect 59967 158147 60001 158175
rect 60029 158147 75299 158175
rect 75327 158147 75361 158175
rect 75389 158147 90659 158175
rect 90687 158147 90721 158175
rect 90749 158147 106019 158175
rect 106047 158147 106081 158175
rect 106109 158147 121379 158175
rect 121407 158147 121441 158175
rect 121469 158147 136739 158175
rect 136767 158147 136801 158175
rect 136829 158147 156485 158175
rect 156513 158147 156547 158175
rect 156575 158147 156609 158175
rect 156637 158147 156671 158175
rect 156699 158147 165485 158175
rect 165513 158147 165547 158175
rect 165575 158147 165609 158175
rect 165637 158147 165671 158175
rect 165699 158147 174485 158175
rect 174513 158147 174547 158175
rect 174575 158147 174609 158175
rect 174637 158147 174671 158175
rect 174699 158147 183485 158175
rect 183513 158147 183547 158175
rect 183575 158147 183609 158175
rect 183637 158147 183671 158175
rect 183699 158147 192485 158175
rect 192513 158147 192547 158175
rect 192575 158147 192609 158175
rect 192637 158147 192671 158175
rect 192699 158147 201485 158175
rect 201513 158147 201547 158175
rect 201575 158147 201609 158175
rect 201637 158147 201671 158175
rect 201699 158147 210485 158175
rect 210513 158147 210547 158175
rect 210575 158147 210609 158175
rect 210637 158147 210671 158175
rect 210699 158147 219485 158175
rect 219513 158147 219547 158175
rect 219575 158147 219609 158175
rect 219637 158147 219671 158175
rect 219699 158147 228485 158175
rect 228513 158147 228547 158175
rect 228575 158147 228609 158175
rect 228637 158147 228671 158175
rect 228699 158147 237485 158175
rect 237513 158147 237547 158175
rect 237575 158147 237609 158175
rect 237637 158147 237671 158175
rect 237699 158147 246485 158175
rect 246513 158147 246547 158175
rect 246575 158147 246609 158175
rect 246637 158147 246671 158175
rect 246699 158147 255485 158175
rect 255513 158147 255547 158175
rect 255575 158147 255609 158175
rect 255637 158147 255671 158175
rect 255699 158147 264485 158175
rect 264513 158147 264547 158175
rect 264575 158147 264609 158175
rect 264637 158147 264671 158175
rect 264699 158147 273485 158175
rect 273513 158147 273547 158175
rect 273575 158147 273609 158175
rect 273637 158147 273671 158175
rect 273699 158147 282485 158175
rect 282513 158147 282547 158175
rect 282575 158147 282609 158175
rect 282637 158147 282671 158175
rect 282699 158147 291485 158175
rect 291513 158147 291547 158175
rect 291575 158147 291609 158175
rect 291637 158147 291671 158175
rect 291699 158147 298728 158175
rect 298756 158147 298790 158175
rect 298818 158147 298852 158175
rect 298880 158147 298914 158175
rect 298942 158147 298990 158175
rect -958 158113 298990 158147
rect -958 158085 -910 158113
rect -882 158085 -848 158113
rect -820 158085 -786 158113
rect -758 158085 -724 158113
rect -696 158085 3485 158113
rect 3513 158085 3547 158113
rect 3575 158085 3609 158113
rect 3637 158085 3671 158113
rect 3699 158085 12485 158113
rect 12513 158085 12547 158113
rect 12575 158085 12609 158113
rect 12637 158085 12671 158113
rect 12699 158085 21485 158113
rect 21513 158085 21547 158113
rect 21575 158085 21609 158113
rect 21637 158085 21671 158113
rect 21699 158085 30485 158113
rect 30513 158085 30547 158113
rect 30575 158085 30609 158113
rect 30637 158085 30671 158113
rect 30699 158085 39485 158113
rect 39513 158085 39547 158113
rect 39575 158085 39609 158113
rect 39637 158085 39671 158113
rect 39699 158085 48485 158113
rect 48513 158085 48547 158113
rect 48575 158085 48609 158113
rect 48637 158085 48671 158113
rect 48699 158085 59939 158113
rect 59967 158085 60001 158113
rect 60029 158085 75299 158113
rect 75327 158085 75361 158113
rect 75389 158085 90659 158113
rect 90687 158085 90721 158113
rect 90749 158085 106019 158113
rect 106047 158085 106081 158113
rect 106109 158085 121379 158113
rect 121407 158085 121441 158113
rect 121469 158085 136739 158113
rect 136767 158085 136801 158113
rect 136829 158085 156485 158113
rect 156513 158085 156547 158113
rect 156575 158085 156609 158113
rect 156637 158085 156671 158113
rect 156699 158085 165485 158113
rect 165513 158085 165547 158113
rect 165575 158085 165609 158113
rect 165637 158085 165671 158113
rect 165699 158085 174485 158113
rect 174513 158085 174547 158113
rect 174575 158085 174609 158113
rect 174637 158085 174671 158113
rect 174699 158085 183485 158113
rect 183513 158085 183547 158113
rect 183575 158085 183609 158113
rect 183637 158085 183671 158113
rect 183699 158085 192485 158113
rect 192513 158085 192547 158113
rect 192575 158085 192609 158113
rect 192637 158085 192671 158113
rect 192699 158085 201485 158113
rect 201513 158085 201547 158113
rect 201575 158085 201609 158113
rect 201637 158085 201671 158113
rect 201699 158085 210485 158113
rect 210513 158085 210547 158113
rect 210575 158085 210609 158113
rect 210637 158085 210671 158113
rect 210699 158085 219485 158113
rect 219513 158085 219547 158113
rect 219575 158085 219609 158113
rect 219637 158085 219671 158113
rect 219699 158085 228485 158113
rect 228513 158085 228547 158113
rect 228575 158085 228609 158113
rect 228637 158085 228671 158113
rect 228699 158085 237485 158113
rect 237513 158085 237547 158113
rect 237575 158085 237609 158113
rect 237637 158085 237671 158113
rect 237699 158085 246485 158113
rect 246513 158085 246547 158113
rect 246575 158085 246609 158113
rect 246637 158085 246671 158113
rect 246699 158085 255485 158113
rect 255513 158085 255547 158113
rect 255575 158085 255609 158113
rect 255637 158085 255671 158113
rect 255699 158085 264485 158113
rect 264513 158085 264547 158113
rect 264575 158085 264609 158113
rect 264637 158085 264671 158113
rect 264699 158085 273485 158113
rect 273513 158085 273547 158113
rect 273575 158085 273609 158113
rect 273637 158085 273671 158113
rect 273699 158085 282485 158113
rect 282513 158085 282547 158113
rect 282575 158085 282609 158113
rect 282637 158085 282671 158113
rect 282699 158085 291485 158113
rect 291513 158085 291547 158113
rect 291575 158085 291609 158113
rect 291637 158085 291671 158113
rect 291699 158085 298728 158113
rect 298756 158085 298790 158113
rect 298818 158085 298852 158113
rect 298880 158085 298914 158113
rect 298942 158085 298990 158113
rect -958 158051 298990 158085
rect -958 158023 -910 158051
rect -882 158023 -848 158051
rect -820 158023 -786 158051
rect -758 158023 -724 158051
rect -696 158023 3485 158051
rect 3513 158023 3547 158051
rect 3575 158023 3609 158051
rect 3637 158023 3671 158051
rect 3699 158023 12485 158051
rect 12513 158023 12547 158051
rect 12575 158023 12609 158051
rect 12637 158023 12671 158051
rect 12699 158023 21485 158051
rect 21513 158023 21547 158051
rect 21575 158023 21609 158051
rect 21637 158023 21671 158051
rect 21699 158023 30485 158051
rect 30513 158023 30547 158051
rect 30575 158023 30609 158051
rect 30637 158023 30671 158051
rect 30699 158023 39485 158051
rect 39513 158023 39547 158051
rect 39575 158023 39609 158051
rect 39637 158023 39671 158051
rect 39699 158023 48485 158051
rect 48513 158023 48547 158051
rect 48575 158023 48609 158051
rect 48637 158023 48671 158051
rect 48699 158023 59939 158051
rect 59967 158023 60001 158051
rect 60029 158023 75299 158051
rect 75327 158023 75361 158051
rect 75389 158023 90659 158051
rect 90687 158023 90721 158051
rect 90749 158023 106019 158051
rect 106047 158023 106081 158051
rect 106109 158023 121379 158051
rect 121407 158023 121441 158051
rect 121469 158023 136739 158051
rect 136767 158023 136801 158051
rect 136829 158023 156485 158051
rect 156513 158023 156547 158051
rect 156575 158023 156609 158051
rect 156637 158023 156671 158051
rect 156699 158023 165485 158051
rect 165513 158023 165547 158051
rect 165575 158023 165609 158051
rect 165637 158023 165671 158051
rect 165699 158023 174485 158051
rect 174513 158023 174547 158051
rect 174575 158023 174609 158051
rect 174637 158023 174671 158051
rect 174699 158023 183485 158051
rect 183513 158023 183547 158051
rect 183575 158023 183609 158051
rect 183637 158023 183671 158051
rect 183699 158023 192485 158051
rect 192513 158023 192547 158051
rect 192575 158023 192609 158051
rect 192637 158023 192671 158051
rect 192699 158023 201485 158051
rect 201513 158023 201547 158051
rect 201575 158023 201609 158051
rect 201637 158023 201671 158051
rect 201699 158023 210485 158051
rect 210513 158023 210547 158051
rect 210575 158023 210609 158051
rect 210637 158023 210671 158051
rect 210699 158023 219485 158051
rect 219513 158023 219547 158051
rect 219575 158023 219609 158051
rect 219637 158023 219671 158051
rect 219699 158023 228485 158051
rect 228513 158023 228547 158051
rect 228575 158023 228609 158051
rect 228637 158023 228671 158051
rect 228699 158023 237485 158051
rect 237513 158023 237547 158051
rect 237575 158023 237609 158051
rect 237637 158023 237671 158051
rect 237699 158023 246485 158051
rect 246513 158023 246547 158051
rect 246575 158023 246609 158051
rect 246637 158023 246671 158051
rect 246699 158023 255485 158051
rect 255513 158023 255547 158051
rect 255575 158023 255609 158051
rect 255637 158023 255671 158051
rect 255699 158023 264485 158051
rect 264513 158023 264547 158051
rect 264575 158023 264609 158051
rect 264637 158023 264671 158051
rect 264699 158023 273485 158051
rect 273513 158023 273547 158051
rect 273575 158023 273609 158051
rect 273637 158023 273671 158051
rect 273699 158023 282485 158051
rect 282513 158023 282547 158051
rect 282575 158023 282609 158051
rect 282637 158023 282671 158051
rect 282699 158023 291485 158051
rect 291513 158023 291547 158051
rect 291575 158023 291609 158051
rect 291637 158023 291671 158051
rect 291699 158023 298728 158051
rect 298756 158023 298790 158051
rect 298818 158023 298852 158051
rect 298880 158023 298914 158051
rect 298942 158023 298990 158051
rect -958 157989 298990 158023
rect -958 157961 -910 157989
rect -882 157961 -848 157989
rect -820 157961 -786 157989
rect -758 157961 -724 157989
rect -696 157961 3485 157989
rect 3513 157961 3547 157989
rect 3575 157961 3609 157989
rect 3637 157961 3671 157989
rect 3699 157961 12485 157989
rect 12513 157961 12547 157989
rect 12575 157961 12609 157989
rect 12637 157961 12671 157989
rect 12699 157961 21485 157989
rect 21513 157961 21547 157989
rect 21575 157961 21609 157989
rect 21637 157961 21671 157989
rect 21699 157961 30485 157989
rect 30513 157961 30547 157989
rect 30575 157961 30609 157989
rect 30637 157961 30671 157989
rect 30699 157961 39485 157989
rect 39513 157961 39547 157989
rect 39575 157961 39609 157989
rect 39637 157961 39671 157989
rect 39699 157961 48485 157989
rect 48513 157961 48547 157989
rect 48575 157961 48609 157989
rect 48637 157961 48671 157989
rect 48699 157961 59939 157989
rect 59967 157961 60001 157989
rect 60029 157961 75299 157989
rect 75327 157961 75361 157989
rect 75389 157961 90659 157989
rect 90687 157961 90721 157989
rect 90749 157961 106019 157989
rect 106047 157961 106081 157989
rect 106109 157961 121379 157989
rect 121407 157961 121441 157989
rect 121469 157961 136739 157989
rect 136767 157961 136801 157989
rect 136829 157961 156485 157989
rect 156513 157961 156547 157989
rect 156575 157961 156609 157989
rect 156637 157961 156671 157989
rect 156699 157961 165485 157989
rect 165513 157961 165547 157989
rect 165575 157961 165609 157989
rect 165637 157961 165671 157989
rect 165699 157961 174485 157989
rect 174513 157961 174547 157989
rect 174575 157961 174609 157989
rect 174637 157961 174671 157989
rect 174699 157961 183485 157989
rect 183513 157961 183547 157989
rect 183575 157961 183609 157989
rect 183637 157961 183671 157989
rect 183699 157961 192485 157989
rect 192513 157961 192547 157989
rect 192575 157961 192609 157989
rect 192637 157961 192671 157989
rect 192699 157961 201485 157989
rect 201513 157961 201547 157989
rect 201575 157961 201609 157989
rect 201637 157961 201671 157989
rect 201699 157961 210485 157989
rect 210513 157961 210547 157989
rect 210575 157961 210609 157989
rect 210637 157961 210671 157989
rect 210699 157961 219485 157989
rect 219513 157961 219547 157989
rect 219575 157961 219609 157989
rect 219637 157961 219671 157989
rect 219699 157961 228485 157989
rect 228513 157961 228547 157989
rect 228575 157961 228609 157989
rect 228637 157961 228671 157989
rect 228699 157961 237485 157989
rect 237513 157961 237547 157989
rect 237575 157961 237609 157989
rect 237637 157961 237671 157989
rect 237699 157961 246485 157989
rect 246513 157961 246547 157989
rect 246575 157961 246609 157989
rect 246637 157961 246671 157989
rect 246699 157961 255485 157989
rect 255513 157961 255547 157989
rect 255575 157961 255609 157989
rect 255637 157961 255671 157989
rect 255699 157961 264485 157989
rect 264513 157961 264547 157989
rect 264575 157961 264609 157989
rect 264637 157961 264671 157989
rect 264699 157961 273485 157989
rect 273513 157961 273547 157989
rect 273575 157961 273609 157989
rect 273637 157961 273671 157989
rect 273699 157961 282485 157989
rect 282513 157961 282547 157989
rect 282575 157961 282609 157989
rect 282637 157961 282671 157989
rect 282699 157961 291485 157989
rect 291513 157961 291547 157989
rect 291575 157961 291609 157989
rect 291637 157961 291671 157989
rect 291699 157961 298728 157989
rect 298756 157961 298790 157989
rect 298818 157961 298852 157989
rect 298880 157961 298914 157989
rect 298942 157961 298990 157989
rect -958 157913 298990 157961
rect -958 155175 298990 155223
rect -958 155147 -430 155175
rect -402 155147 -368 155175
rect -340 155147 -306 155175
rect -278 155147 -244 155175
rect -216 155147 1625 155175
rect 1653 155147 1687 155175
rect 1715 155147 1749 155175
rect 1777 155147 1811 155175
rect 1839 155147 10625 155175
rect 10653 155147 10687 155175
rect 10715 155147 10749 155175
rect 10777 155147 10811 155175
rect 10839 155147 19625 155175
rect 19653 155147 19687 155175
rect 19715 155147 19749 155175
rect 19777 155147 19811 155175
rect 19839 155147 28625 155175
rect 28653 155147 28687 155175
rect 28715 155147 28749 155175
rect 28777 155147 28811 155175
rect 28839 155147 37625 155175
rect 37653 155147 37687 155175
rect 37715 155147 37749 155175
rect 37777 155147 37811 155175
rect 37839 155147 46625 155175
rect 46653 155147 46687 155175
rect 46715 155147 46749 155175
rect 46777 155147 46811 155175
rect 46839 155147 52259 155175
rect 52287 155147 52321 155175
rect 52349 155147 67619 155175
rect 67647 155147 67681 155175
rect 67709 155147 82979 155175
rect 83007 155147 83041 155175
rect 83069 155147 98339 155175
rect 98367 155147 98401 155175
rect 98429 155147 113699 155175
rect 113727 155147 113761 155175
rect 113789 155147 129059 155175
rect 129087 155147 129121 155175
rect 129149 155147 144419 155175
rect 144447 155147 144481 155175
rect 144509 155147 154625 155175
rect 154653 155147 154687 155175
rect 154715 155147 154749 155175
rect 154777 155147 154811 155175
rect 154839 155147 163625 155175
rect 163653 155147 163687 155175
rect 163715 155147 163749 155175
rect 163777 155147 163811 155175
rect 163839 155147 172625 155175
rect 172653 155147 172687 155175
rect 172715 155147 172749 155175
rect 172777 155147 172811 155175
rect 172839 155147 181625 155175
rect 181653 155147 181687 155175
rect 181715 155147 181749 155175
rect 181777 155147 181811 155175
rect 181839 155147 190625 155175
rect 190653 155147 190687 155175
rect 190715 155147 190749 155175
rect 190777 155147 190811 155175
rect 190839 155147 199625 155175
rect 199653 155147 199687 155175
rect 199715 155147 199749 155175
rect 199777 155147 199811 155175
rect 199839 155147 208625 155175
rect 208653 155147 208687 155175
rect 208715 155147 208749 155175
rect 208777 155147 208811 155175
rect 208839 155147 217625 155175
rect 217653 155147 217687 155175
rect 217715 155147 217749 155175
rect 217777 155147 217811 155175
rect 217839 155147 226625 155175
rect 226653 155147 226687 155175
rect 226715 155147 226749 155175
rect 226777 155147 226811 155175
rect 226839 155147 235625 155175
rect 235653 155147 235687 155175
rect 235715 155147 235749 155175
rect 235777 155147 235811 155175
rect 235839 155147 244625 155175
rect 244653 155147 244687 155175
rect 244715 155147 244749 155175
rect 244777 155147 244811 155175
rect 244839 155147 253625 155175
rect 253653 155147 253687 155175
rect 253715 155147 253749 155175
rect 253777 155147 253811 155175
rect 253839 155147 262625 155175
rect 262653 155147 262687 155175
rect 262715 155147 262749 155175
rect 262777 155147 262811 155175
rect 262839 155147 271625 155175
rect 271653 155147 271687 155175
rect 271715 155147 271749 155175
rect 271777 155147 271811 155175
rect 271839 155147 280625 155175
rect 280653 155147 280687 155175
rect 280715 155147 280749 155175
rect 280777 155147 280811 155175
rect 280839 155147 289625 155175
rect 289653 155147 289687 155175
rect 289715 155147 289749 155175
rect 289777 155147 289811 155175
rect 289839 155147 298248 155175
rect 298276 155147 298310 155175
rect 298338 155147 298372 155175
rect 298400 155147 298434 155175
rect 298462 155147 298990 155175
rect -958 155113 298990 155147
rect -958 155085 -430 155113
rect -402 155085 -368 155113
rect -340 155085 -306 155113
rect -278 155085 -244 155113
rect -216 155085 1625 155113
rect 1653 155085 1687 155113
rect 1715 155085 1749 155113
rect 1777 155085 1811 155113
rect 1839 155085 10625 155113
rect 10653 155085 10687 155113
rect 10715 155085 10749 155113
rect 10777 155085 10811 155113
rect 10839 155085 19625 155113
rect 19653 155085 19687 155113
rect 19715 155085 19749 155113
rect 19777 155085 19811 155113
rect 19839 155085 28625 155113
rect 28653 155085 28687 155113
rect 28715 155085 28749 155113
rect 28777 155085 28811 155113
rect 28839 155085 37625 155113
rect 37653 155085 37687 155113
rect 37715 155085 37749 155113
rect 37777 155085 37811 155113
rect 37839 155085 46625 155113
rect 46653 155085 46687 155113
rect 46715 155085 46749 155113
rect 46777 155085 46811 155113
rect 46839 155085 52259 155113
rect 52287 155085 52321 155113
rect 52349 155085 67619 155113
rect 67647 155085 67681 155113
rect 67709 155085 82979 155113
rect 83007 155085 83041 155113
rect 83069 155085 98339 155113
rect 98367 155085 98401 155113
rect 98429 155085 113699 155113
rect 113727 155085 113761 155113
rect 113789 155085 129059 155113
rect 129087 155085 129121 155113
rect 129149 155085 144419 155113
rect 144447 155085 144481 155113
rect 144509 155085 154625 155113
rect 154653 155085 154687 155113
rect 154715 155085 154749 155113
rect 154777 155085 154811 155113
rect 154839 155085 163625 155113
rect 163653 155085 163687 155113
rect 163715 155085 163749 155113
rect 163777 155085 163811 155113
rect 163839 155085 172625 155113
rect 172653 155085 172687 155113
rect 172715 155085 172749 155113
rect 172777 155085 172811 155113
rect 172839 155085 181625 155113
rect 181653 155085 181687 155113
rect 181715 155085 181749 155113
rect 181777 155085 181811 155113
rect 181839 155085 190625 155113
rect 190653 155085 190687 155113
rect 190715 155085 190749 155113
rect 190777 155085 190811 155113
rect 190839 155085 199625 155113
rect 199653 155085 199687 155113
rect 199715 155085 199749 155113
rect 199777 155085 199811 155113
rect 199839 155085 208625 155113
rect 208653 155085 208687 155113
rect 208715 155085 208749 155113
rect 208777 155085 208811 155113
rect 208839 155085 217625 155113
rect 217653 155085 217687 155113
rect 217715 155085 217749 155113
rect 217777 155085 217811 155113
rect 217839 155085 226625 155113
rect 226653 155085 226687 155113
rect 226715 155085 226749 155113
rect 226777 155085 226811 155113
rect 226839 155085 235625 155113
rect 235653 155085 235687 155113
rect 235715 155085 235749 155113
rect 235777 155085 235811 155113
rect 235839 155085 244625 155113
rect 244653 155085 244687 155113
rect 244715 155085 244749 155113
rect 244777 155085 244811 155113
rect 244839 155085 253625 155113
rect 253653 155085 253687 155113
rect 253715 155085 253749 155113
rect 253777 155085 253811 155113
rect 253839 155085 262625 155113
rect 262653 155085 262687 155113
rect 262715 155085 262749 155113
rect 262777 155085 262811 155113
rect 262839 155085 271625 155113
rect 271653 155085 271687 155113
rect 271715 155085 271749 155113
rect 271777 155085 271811 155113
rect 271839 155085 280625 155113
rect 280653 155085 280687 155113
rect 280715 155085 280749 155113
rect 280777 155085 280811 155113
rect 280839 155085 289625 155113
rect 289653 155085 289687 155113
rect 289715 155085 289749 155113
rect 289777 155085 289811 155113
rect 289839 155085 298248 155113
rect 298276 155085 298310 155113
rect 298338 155085 298372 155113
rect 298400 155085 298434 155113
rect 298462 155085 298990 155113
rect -958 155051 298990 155085
rect -958 155023 -430 155051
rect -402 155023 -368 155051
rect -340 155023 -306 155051
rect -278 155023 -244 155051
rect -216 155023 1625 155051
rect 1653 155023 1687 155051
rect 1715 155023 1749 155051
rect 1777 155023 1811 155051
rect 1839 155023 10625 155051
rect 10653 155023 10687 155051
rect 10715 155023 10749 155051
rect 10777 155023 10811 155051
rect 10839 155023 19625 155051
rect 19653 155023 19687 155051
rect 19715 155023 19749 155051
rect 19777 155023 19811 155051
rect 19839 155023 28625 155051
rect 28653 155023 28687 155051
rect 28715 155023 28749 155051
rect 28777 155023 28811 155051
rect 28839 155023 37625 155051
rect 37653 155023 37687 155051
rect 37715 155023 37749 155051
rect 37777 155023 37811 155051
rect 37839 155023 46625 155051
rect 46653 155023 46687 155051
rect 46715 155023 46749 155051
rect 46777 155023 46811 155051
rect 46839 155023 52259 155051
rect 52287 155023 52321 155051
rect 52349 155023 67619 155051
rect 67647 155023 67681 155051
rect 67709 155023 82979 155051
rect 83007 155023 83041 155051
rect 83069 155023 98339 155051
rect 98367 155023 98401 155051
rect 98429 155023 113699 155051
rect 113727 155023 113761 155051
rect 113789 155023 129059 155051
rect 129087 155023 129121 155051
rect 129149 155023 144419 155051
rect 144447 155023 144481 155051
rect 144509 155023 154625 155051
rect 154653 155023 154687 155051
rect 154715 155023 154749 155051
rect 154777 155023 154811 155051
rect 154839 155023 163625 155051
rect 163653 155023 163687 155051
rect 163715 155023 163749 155051
rect 163777 155023 163811 155051
rect 163839 155023 172625 155051
rect 172653 155023 172687 155051
rect 172715 155023 172749 155051
rect 172777 155023 172811 155051
rect 172839 155023 181625 155051
rect 181653 155023 181687 155051
rect 181715 155023 181749 155051
rect 181777 155023 181811 155051
rect 181839 155023 190625 155051
rect 190653 155023 190687 155051
rect 190715 155023 190749 155051
rect 190777 155023 190811 155051
rect 190839 155023 199625 155051
rect 199653 155023 199687 155051
rect 199715 155023 199749 155051
rect 199777 155023 199811 155051
rect 199839 155023 208625 155051
rect 208653 155023 208687 155051
rect 208715 155023 208749 155051
rect 208777 155023 208811 155051
rect 208839 155023 217625 155051
rect 217653 155023 217687 155051
rect 217715 155023 217749 155051
rect 217777 155023 217811 155051
rect 217839 155023 226625 155051
rect 226653 155023 226687 155051
rect 226715 155023 226749 155051
rect 226777 155023 226811 155051
rect 226839 155023 235625 155051
rect 235653 155023 235687 155051
rect 235715 155023 235749 155051
rect 235777 155023 235811 155051
rect 235839 155023 244625 155051
rect 244653 155023 244687 155051
rect 244715 155023 244749 155051
rect 244777 155023 244811 155051
rect 244839 155023 253625 155051
rect 253653 155023 253687 155051
rect 253715 155023 253749 155051
rect 253777 155023 253811 155051
rect 253839 155023 262625 155051
rect 262653 155023 262687 155051
rect 262715 155023 262749 155051
rect 262777 155023 262811 155051
rect 262839 155023 271625 155051
rect 271653 155023 271687 155051
rect 271715 155023 271749 155051
rect 271777 155023 271811 155051
rect 271839 155023 280625 155051
rect 280653 155023 280687 155051
rect 280715 155023 280749 155051
rect 280777 155023 280811 155051
rect 280839 155023 289625 155051
rect 289653 155023 289687 155051
rect 289715 155023 289749 155051
rect 289777 155023 289811 155051
rect 289839 155023 298248 155051
rect 298276 155023 298310 155051
rect 298338 155023 298372 155051
rect 298400 155023 298434 155051
rect 298462 155023 298990 155051
rect -958 154989 298990 155023
rect -958 154961 -430 154989
rect -402 154961 -368 154989
rect -340 154961 -306 154989
rect -278 154961 -244 154989
rect -216 154961 1625 154989
rect 1653 154961 1687 154989
rect 1715 154961 1749 154989
rect 1777 154961 1811 154989
rect 1839 154961 10625 154989
rect 10653 154961 10687 154989
rect 10715 154961 10749 154989
rect 10777 154961 10811 154989
rect 10839 154961 19625 154989
rect 19653 154961 19687 154989
rect 19715 154961 19749 154989
rect 19777 154961 19811 154989
rect 19839 154961 28625 154989
rect 28653 154961 28687 154989
rect 28715 154961 28749 154989
rect 28777 154961 28811 154989
rect 28839 154961 37625 154989
rect 37653 154961 37687 154989
rect 37715 154961 37749 154989
rect 37777 154961 37811 154989
rect 37839 154961 46625 154989
rect 46653 154961 46687 154989
rect 46715 154961 46749 154989
rect 46777 154961 46811 154989
rect 46839 154961 52259 154989
rect 52287 154961 52321 154989
rect 52349 154961 67619 154989
rect 67647 154961 67681 154989
rect 67709 154961 82979 154989
rect 83007 154961 83041 154989
rect 83069 154961 98339 154989
rect 98367 154961 98401 154989
rect 98429 154961 113699 154989
rect 113727 154961 113761 154989
rect 113789 154961 129059 154989
rect 129087 154961 129121 154989
rect 129149 154961 144419 154989
rect 144447 154961 144481 154989
rect 144509 154961 154625 154989
rect 154653 154961 154687 154989
rect 154715 154961 154749 154989
rect 154777 154961 154811 154989
rect 154839 154961 163625 154989
rect 163653 154961 163687 154989
rect 163715 154961 163749 154989
rect 163777 154961 163811 154989
rect 163839 154961 172625 154989
rect 172653 154961 172687 154989
rect 172715 154961 172749 154989
rect 172777 154961 172811 154989
rect 172839 154961 181625 154989
rect 181653 154961 181687 154989
rect 181715 154961 181749 154989
rect 181777 154961 181811 154989
rect 181839 154961 190625 154989
rect 190653 154961 190687 154989
rect 190715 154961 190749 154989
rect 190777 154961 190811 154989
rect 190839 154961 199625 154989
rect 199653 154961 199687 154989
rect 199715 154961 199749 154989
rect 199777 154961 199811 154989
rect 199839 154961 208625 154989
rect 208653 154961 208687 154989
rect 208715 154961 208749 154989
rect 208777 154961 208811 154989
rect 208839 154961 217625 154989
rect 217653 154961 217687 154989
rect 217715 154961 217749 154989
rect 217777 154961 217811 154989
rect 217839 154961 226625 154989
rect 226653 154961 226687 154989
rect 226715 154961 226749 154989
rect 226777 154961 226811 154989
rect 226839 154961 235625 154989
rect 235653 154961 235687 154989
rect 235715 154961 235749 154989
rect 235777 154961 235811 154989
rect 235839 154961 244625 154989
rect 244653 154961 244687 154989
rect 244715 154961 244749 154989
rect 244777 154961 244811 154989
rect 244839 154961 253625 154989
rect 253653 154961 253687 154989
rect 253715 154961 253749 154989
rect 253777 154961 253811 154989
rect 253839 154961 262625 154989
rect 262653 154961 262687 154989
rect 262715 154961 262749 154989
rect 262777 154961 262811 154989
rect 262839 154961 271625 154989
rect 271653 154961 271687 154989
rect 271715 154961 271749 154989
rect 271777 154961 271811 154989
rect 271839 154961 280625 154989
rect 280653 154961 280687 154989
rect 280715 154961 280749 154989
rect 280777 154961 280811 154989
rect 280839 154961 289625 154989
rect 289653 154961 289687 154989
rect 289715 154961 289749 154989
rect 289777 154961 289811 154989
rect 289839 154961 298248 154989
rect 298276 154961 298310 154989
rect 298338 154961 298372 154989
rect 298400 154961 298434 154989
rect 298462 154961 298990 154989
rect -958 154913 298990 154961
rect -958 149175 298990 149223
rect -958 149147 -910 149175
rect -882 149147 -848 149175
rect -820 149147 -786 149175
rect -758 149147 -724 149175
rect -696 149147 3485 149175
rect 3513 149147 3547 149175
rect 3575 149147 3609 149175
rect 3637 149147 3671 149175
rect 3699 149147 12485 149175
rect 12513 149147 12547 149175
rect 12575 149147 12609 149175
rect 12637 149147 12671 149175
rect 12699 149147 21485 149175
rect 21513 149147 21547 149175
rect 21575 149147 21609 149175
rect 21637 149147 21671 149175
rect 21699 149147 30485 149175
rect 30513 149147 30547 149175
rect 30575 149147 30609 149175
rect 30637 149147 30671 149175
rect 30699 149147 39485 149175
rect 39513 149147 39547 149175
rect 39575 149147 39609 149175
rect 39637 149147 39671 149175
rect 39699 149147 48485 149175
rect 48513 149147 48547 149175
rect 48575 149147 48609 149175
rect 48637 149147 48671 149175
rect 48699 149147 59939 149175
rect 59967 149147 60001 149175
rect 60029 149147 75299 149175
rect 75327 149147 75361 149175
rect 75389 149147 90659 149175
rect 90687 149147 90721 149175
rect 90749 149147 106019 149175
rect 106047 149147 106081 149175
rect 106109 149147 121379 149175
rect 121407 149147 121441 149175
rect 121469 149147 136739 149175
rect 136767 149147 136801 149175
rect 136829 149147 156485 149175
rect 156513 149147 156547 149175
rect 156575 149147 156609 149175
rect 156637 149147 156671 149175
rect 156699 149147 165485 149175
rect 165513 149147 165547 149175
rect 165575 149147 165609 149175
rect 165637 149147 165671 149175
rect 165699 149147 174485 149175
rect 174513 149147 174547 149175
rect 174575 149147 174609 149175
rect 174637 149147 174671 149175
rect 174699 149147 183485 149175
rect 183513 149147 183547 149175
rect 183575 149147 183609 149175
rect 183637 149147 183671 149175
rect 183699 149147 192485 149175
rect 192513 149147 192547 149175
rect 192575 149147 192609 149175
rect 192637 149147 192671 149175
rect 192699 149147 201485 149175
rect 201513 149147 201547 149175
rect 201575 149147 201609 149175
rect 201637 149147 201671 149175
rect 201699 149147 210485 149175
rect 210513 149147 210547 149175
rect 210575 149147 210609 149175
rect 210637 149147 210671 149175
rect 210699 149147 219485 149175
rect 219513 149147 219547 149175
rect 219575 149147 219609 149175
rect 219637 149147 219671 149175
rect 219699 149147 228485 149175
rect 228513 149147 228547 149175
rect 228575 149147 228609 149175
rect 228637 149147 228671 149175
rect 228699 149147 237485 149175
rect 237513 149147 237547 149175
rect 237575 149147 237609 149175
rect 237637 149147 237671 149175
rect 237699 149147 246485 149175
rect 246513 149147 246547 149175
rect 246575 149147 246609 149175
rect 246637 149147 246671 149175
rect 246699 149147 255485 149175
rect 255513 149147 255547 149175
rect 255575 149147 255609 149175
rect 255637 149147 255671 149175
rect 255699 149147 264485 149175
rect 264513 149147 264547 149175
rect 264575 149147 264609 149175
rect 264637 149147 264671 149175
rect 264699 149147 273485 149175
rect 273513 149147 273547 149175
rect 273575 149147 273609 149175
rect 273637 149147 273671 149175
rect 273699 149147 282485 149175
rect 282513 149147 282547 149175
rect 282575 149147 282609 149175
rect 282637 149147 282671 149175
rect 282699 149147 291485 149175
rect 291513 149147 291547 149175
rect 291575 149147 291609 149175
rect 291637 149147 291671 149175
rect 291699 149147 298728 149175
rect 298756 149147 298790 149175
rect 298818 149147 298852 149175
rect 298880 149147 298914 149175
rect 298942 149147 298990 149175
rect -958 149113 298990 149147
rect -958 149085 -910 149113
rect -882 149085 -848 149113
rect -820 149085 -786 149113
rect -758 149085 -724 149113
rect -696 149085 3485 149113
rect 3513 149085 3547 149113
rect 3575 149085 3609 149113
rect 3637 149085 3671 149113
rect 3699 149085 12485 149113
rect 12513 149085 12547 149113
rect 12575 149085 12609 149113
rect 12637 149085 12671 149113
rect 12699 149085 21485 149113
rect 21513 149085 21547 149113
rect 21575 149085 21609 149113
rect 21637 149085 21671 149113
rect 21699 149085 30485 149113
rect 30513 149085 30547 149113
rect 30575 149085 30609 149113
rect 30637 149085 30671 149113
rect 30699 149085 39485 149113
rect 39513 149085 39547 149113
rect 39575 149085 39609 149113
rect 39637 149085 39671 149113
rect 39699 149085 48485 149113
rect 48513 149085 48547 149113
rect 48575 149085 48609 149113
rect 48637 149085 48671 149113
rect 48699 149085 59939 149113
rect 59967 149085 60001 149113
rect 60029 149085 75299 149113
rect 75327 149085 75361 149113
rect 75389 149085 90659 149113
rect 90687 149085 90721 149113
rect 90749 149085 106019 149113
rect 106047 149085 106081 149113
rect 106109 149085 121379 149113
rect 121407 149085 121441 149113
rect 121469 149085 136739 149113
rect 136767 149085 136801 149113
rect 136829 149085 156485 149113
rect 156513 149085 156547 149113
rect 156575 149085 156609 149113
rect 156637 149085 156671 149113
rect 156699 149085 165485 149113
rect 165513 149085 165547 149113
rect 165575 149085 165609 149113
rect 165637 149085 165671 149113
rect 165699 149085 174485 149113
rect 174513 149085 174547 149113
rect 174575 149085 174609 149113
rect 174637 149085 174671 149113
rect 174699 149085 183485 149113
rect 183513 149085 183547 149113
rect 183575 149085 183609 149113
rect 183637 149085 183671 149113
rect 183699 149085 192485 149113
rect 192513 149085 192547 149113
rect 192575 149085 192609 149113
rect 192637 149085 192671 149113
rect 192699 149085 201485 149113
rect 201513 149085 201547 149113
rect 201575 149085 201609 149113
rect 201637 149085 201671 149113
rect 201699 149085 210485 149113
rect 210513 149085 210547 149113
rect 210575 149085 210609 149113
rect 210637 149085 210671 149113
rect 210699 149085 219485 149113
rect 219513 149085 219547 149113
rect 219575 149085 219609 149113
rect 219637 149085 219671 149113
rect 219699 149085 228485 149113
rect 228513 149085 228547 149113
rect 228575 149085 228609 149113
rect 228637 149085 228671 149113
rect 228699 149085 237485 149113
rect 237513 149085 237547 149113
rect 237575 149085 237609 149113
rect 237637 149085 237671 149113
rect 237699 149085 246485 149113
rect 246513 149085 246547 149113
rect 246575 149085 246609 149113
rect 246637 149085 246671 149113
rect 246699 149085 255485 149113
rect 255513 149085 255547 149113
rect 255575 149085 255609 149113
rect 255637 149085 255671 149113
rect 255699 149085 264485 149113
rect 264513 149085 264547 149113
rect 264575 149085 264609 149113
rect 264637 149085 264671 149113
rect 264699 149085 273485 149113
rect 273513 149085 273547 149113
rect 273575 149085 273609 149113
rect 273637 149085 273671 149113
rect 273699 149085 282485 149113
rect 282513 149085 282547 149113
rect 282575 149085 282609 149113
rect 282637 149085 282671 149113
rect 282699 149085 291485 149113
rect 291513 149085 291547 149113
rect 291575 149085 291609 149113
rect 291637 149085 291671 149113
rect 291699 149085 298728 149113
rect 298756 149085 298790 149113
rect 298818 149085 298852 149113
rect 298880 149085 298914 149113
rect 298942 149085 298990 149113
rect -958 149051 298990 149085
rect -958 149023 -910 149051
rect -882 149023 -848 149051
rect -820 149023 -786 149051
rect -758 149023 -724 149051
rect -696 149023 3485 149051
rect 3513 149023 3547 149051
rect 3575 149023 3609 149051
rect 3637 149023 3671 149051
rect 3699 149023 12485 149051
rect 12513 149023 12547 149051
rect 12575 149023 12609 149051
rect 12637 149023 12671 149051
rect 12699 149023 21485 149051
rect 21513 149023 21547 149051
rect 21575 149023 21609 149051
rect 21637 149023 21671 149051
rect 21699 149023 30485 149051
rect 30513 149023 30547 149051
rect 30575 149023 30609 149051
rect 30637 149023 30671 149051
rect 30699 149023 39485 149051
rect 39513 149023 39547 149051
rect 39575 149023 39609 149051
rect 39637 149023 39671 149051
rect 39699 149023 48485 149051
rect 48513 149023 48547 149051
rect 48575 149023 48609 149051
rect 48637 149023 48671 149051
rect 48699 149023 59939 149051
rect 59967 149023 60001 149051
rect 60029 149023 75299 149051
rect 75327 149023 75361 149051
rect 75389 149023 90659 149051
rect 90687 149023 90721 149051
rect 90749 149023 106019 149051
rect 106047 149023 106081 149051
rect 106109 149023 121379 149051
rect 121407 149023 121441 149051
rect 121469 149023 136739 149051
rect 136767 149023 136801 149051
rect 136829 149023 156485 149051
rect 156513 149023 156547 149051
rect 156575 149023 156609 149051
rect 156637 149023 156671 149051
rect 156699 149023 165485 149051
rect 165513 149023 165547 149051
rect 165575 149023 165609 149051
rect 165637 149023 165671 149051
rect 165699 149023 174485 149051
rect 174513 149023 174547 149051
rect 174575 149023 174609 149051
rect 174637 149023 174671 149051
rect 174699 149023 183485 149051
rect 183513 149023 183547 149051
rect 183575 149023 183609 149051
rect 183637 149023 183671 149051
rect 183699 149023 192485 149051
rect 192513 149023 192547 149051
rect 192575 149023 192609 149051
rect 192637 149023 192671 149051
rect 192699 149023 201485 149051
rect 201513 149023 201547 149051
rect 201575 149023 201609 149051
rect 201637 149023 201671 149051
rect 201699 149023 210485 149051
rect 210513 149023 210547 149051
rect 210575 149023 210609 149051
rect 210637 149023 210671 149051
rect 210699 149023 219485 149051
rect 219513 149023 219547 149051
rect 219575 149023 219609 149051
rect 219637 149023 219671 149051
rect 219699 149023 228485 149051
rect 228513 149023 228547 149051
rect 228575 149023 228609 149051
rect 228637 149023 228671 149051
rect 228699 149023 237485 149051
rect 237513 149023 237547 149051
rect 237575 149023 237609 149051
rect 237637 149023 237671 149051
rect 237699 149023 246485 149051
rect 246513 149023 246547 149051
rect 246575 149023 246609 149051
rect 246637 149023 246671 149051
rect 246699 149023 255485 149051
rect 255513 149023 255547 149051
rect 255575 149023 255609 149051
rect 255637 149023 255671 149051
rect 255699 149023 264485 149051
rect 264513 149023 264547 149051
rect 264575 149023 264609 149051
rect 264637 149023 264671 149051
rect 264699 149023 273485 149051
rect 273513 149023 273547 149051
rect 273575 149023 273609 149051
rect 273637 149023 273671 149051
rect 273699 149023 282485 149051
rect 282513 149023 282547 149051
rect 282575 149023 282609 149051
rect 282637 149023 282671 149051
rect 282699 149023 291485 149051
rect 291513 149023 291547 149051
rect 291575 149023 291609 149051
rect 291637 149023 291671 149051
rect 291699 149023 298728 149051
rect 298756 149023 298790 149051
rect 298818 149023 298852 149051
rect 298880 149023 298914 149051
rect 298942 149023 298990 149051
rect -958 148989 298990 149023
rect -958 148961 -910 148989
rect -882 148961 -848 148989
rect -820 148961 -786 148989
rect -758 148961 -724 148989
rect -696 148961 3485 148989
rect 3513 148961 3547 148989
rect 3575 148961 3609 148989
rect 3637 148961 3671 148989
rect 3699 148961 12485 148989
rect 12513 148961 12547 148989
rect 12575 148961 12609 148989
rect 12637 148961 12671 148989
rect 12699 148961 21485 148989
rect 21513 148961 21547 148989
rect 21575 148961 21609 148989
rect 21637 148961 21671 148989
rect 21699 148961 30485 148989
rect 30513 148961 30547 148989
rect 30575 148961 30609 148989
rect 30637 148961 30671 148989
rect 30699 148961 39485 148989
rect 39513 148961 39547 148989
rect 39575 148961 39609 148989
rect 39637 148961 39671 148989
rect 39699 148961 48485 148989
rect 48513 148961 48547 148989
rect 48575 148961 48609 148989
rect 48637 148961 48671 148989
rect 48699 148961 59939 148989
rect 59967 148961 60001 148989
rect 60029 148961 75299 148989
rect 75327 148961 75361 148989
rect 75389 148961 90659 148989
rect 90687 148961 90721 148989
rect 90749 148961 106019 148989
rect 106047 148961 106081 148989
rect 106109 148961 121379 148989
rect 121407 148961 121441 148989
rect 121469 148961 136739 148989
rect 136767 148961 136801 148989
rect 136829 148961 156485 148989
rect 156513 148961 156547 148989
rect 156575 148961 156609 148989
rect 156637 148961 156671 148989
rect 156699 148961 165485 148989
rect 165513 148961 165547 148989
rect 165575 148961 165609 148989
rect 165637 148961 165671 148989
rect 165699 148961 174485 148989
rect 174513 148961 174547 148989
rect 174575 148961 174609 148989
rect 174637 148961 174671 148989
rect 174699 148961 183485 148989
rect 183513 148961 183547 148989
rect 183575 148961 183609 148989
rect 183637 148961 183671 148989
rect 183699 148961 192485 148989
rect 192513 148961 192547 148989
rect 192575 148961 192609 148989
rect 192637 148961 192671 148989
rect 192699 148961 201485 148989
rect 201513 148961 201547 148989
rect 201575 148961 201609 148989
rect 201637 148961 201671 148989
rect 201699 148961 210485 148989
rect 210513 148961 210547 148989
rect 210575 148961 210609 148989
rect 210637 148961 210671 148989
rect 210699 148961 219485 148989
rect 219513 148961 219547 148989
rect 219575 148961 219609 148989
rect 219637 148961 219671 148989
rect 219699 148961 228485 148989
rect 228513 148961 228547 148989
rect 228575 148961 228609 148989
rect 228637 148961 228671 148989
rect 228699 148961 237485 148989
rect 237513 148961 237547 148989
rect 237575 148961 237609 148989
rect 237637 148961 237671 148989
rect 237699 148961 246485 148989
rect 246513 148961 246547 148989
rect 246575 148961 246609 148989
rect 246637 148961 246671 148989
rect 246699 148961 255485 148989
rect 255513 148961 255547 148989
rect 255575 148961 255609 148989
rect 255637 148961 255671 148989
rect 255699 148961 264485 148989
rect 264513 148961 264547 148989
rect 264575 148961 264609 148989
rect 264637 148961 264671 148989
rect 264699 148961 273485 148989
rect 273513 148961 273547 148989
rect 273575 148961 273609 148989
rect 273637 148961 273671 148989
rect 273699 148961 282485 148989
rect 282513 148961 282547 148989
rect 282575 148961 282609 148989
rect 282637 148961 282671 148989
rect 282699 148961 291485 148989
rect 291513 148961 291547 148989
rect 291575 148961 291609 148989
rect 291637 148961 291671 148989
rect 291699 148961 298728 148989
rect 298756 148961 298790 148989
rect 298818 148961 298852 148989
rect 298880 148961 298914 148989
rect 298942 148961 298990 148989
rect -958 148913 298990 148961
rect -958 146175 298990 146223
rect -958 146147 -430 146175
rect -402 146147 -368 146175
rect -340 146147 -306 146175
rect -278 146147 -244 146175
rect -216 146147 1625 146175
rect 1653 146147 1687 146175
rect 1715 146147 1749 146175
rect 1777 146147 1811 146175
rect 1839 146147 10625 146175
rect 10653 146147 10687 146175
rect 10715 146147 10749 146175
rect 10777 146147 10811 146175
rect 10839 146147 19625 146175
rect 19653 146147 19687 146175
rect 19715 146147 19749 146175
rect 19777 146147 19811 146175
rect 19839 146147 28625 146175
rect 28653 146147 28687 146175
rect 28715 146147 28749 146175
rect 28777 146147 28811 146175
rect 28839 146147 37625 146175
rect 37653 146147 37687 146175
rect 37715 146147 37749 146175
rect 37777 146147 37811 146175
rect 37839 146147 46625 146175
rect 46653 146147 46687 146175
rect 46715 146147 46749 146175
rect 46777 146147 46811 146175
rect 46839 146147 52259 146175
rect 52287 146147 52321 146175
rect 52349 146147 67619 146175
rect 67647 146147 67681 146175
rect 67709 146147 82979 146175
rect 83007 146147 83041 146175
rect 83069 146147 98339 146175
rect 98367 146147 98401 146175
rect 98429 146147 113699 146175
rect 113727 146147 113761 146175
rect 113789 146147 129059 146175
rect 129087 146147 129121 146175
rect 129149 146147 144419 146175
rect 144447 146147 144481 146175
rect 144509 146147 154625 146175
rect 154653 146147 154687 146175
rect 154715 146147 154749 146175
rect 154777 146147 154811 146175
rect 154839 146147 163625 146175
rect 163653 146147 163687 146175
rect 163715 146147 163749 146175
rect 163777 146147 163811 146175
rect 163839 146147 172625 146175
rect 172653 146147 172687 146175
rect 172715 146147 172749 146175
rect 172777 146147 172811 146175
rect 172839 146147 181625 146175
rect 181653 146147 181687 146175
rect 181715 146147 181749 146175
rect 181777 146147 181811 146175
rect 181839 146147 190625 146175
rect 190653 146147 190687 146175
rect 190715 146147 190749 146175
rect 190777 146147 190811 146175
rect 190839 146147 199625 146175
rect 199653 146147 199687 146175
rect 199715 146147 199749 146175
rect 199777 146147 199811 146175
rect 199839 146147 208625 146175
rect 208653 146147 208687 146175
rect 208715 146147 208749 146175
rect 208777 146147 208811 146175
rect 208839 146147 217625 146175
rect 217653 146147 217687 146175
rect 217715 146147 217749 146175
rect 217777 146147 217811 146175
rect 217839 146147 226625 146175
rect 226653 146147 226687 146175
rect 226715 146147 226749 146175
rect 226777 146147 226811 146175
rect 226839 146147 235625 146175
rect 235653 146147 235687 146175
rect 235715 146147 235749 146175
rect 235777 146147 235811 146175
rect 235839 146147 244625 146175
rect 244653 146147 244687 146175
rect 244715 146147 244749 146175
rect 244777 146147 244811 146175
rect 244839 146147 253625 146175
rect 253653 146147 253687 146175
rect 253715 146147 253749 146175
rect 253777 146147 253811 146175
rect 253839 146147 262625 146175
rect 262653 146147 262687 146175
rect 262715 146147 262749 146175
rect 262777 146147 262811 146175
rect 262839 146147 271625 146175
rect 271653 146147 271687 146175
rect 271715 146147 271749 146175
rect 271777 146147 271811 146175
rect 271839 146147 280625 146175
rect 280653 146147 280687 146175
rect 280715 146147 280749 146175
rect 280777 146147 280811 146175
rect 280839 146147 289625 146175
rect 289653 146147 289687 146175
rect 289715 146147 289749 146175
rect 289777 146147 289811 146175
rect 289839 146147 298248 146175
rect 298276 146147 298310 146175
rect 298338 146147 298372 146175
rect 298400 146147 298434 146175
rect 298462 146147 298990 146175
rect -958 146113 298990 146147
rect -958 146085 -430 146113
rect -402 146085 -368 146113
rect -340 146085 -306 146113
rect -278 146085 -244 146113
rect -216 146085 1625 146113
rect 1653 146085 1687 146113
rect 1715 146085 1749 146113
rect 1777 146085 1811 146113
rect 1839 146085 10625 146113
rect 10653 146085 10687 146113
rect 10715 146085 10749 146113
rect 10777 146085 10811 146113
rect 10839 146085 19625 146113
rect 19653 146085 19687 146113
rect 19715 146085 19749 146113
rect 19777 146085 19811 146113
rect 19839 146085 28625 146113
rect 28653 146085 28687 146113
rect 28715 146085 28749 146113
rect 28777 146085 28811 146113
rect 28839 146085 37625 146113
rect 37653 146085 37687 146113
rect 37715 146085 37749 146113
rect 37777 146085 37811 146113
rect 37839 146085 46625 146113
rect 46653 146085 46687 146113
rect 46715 146085 46749 146113
rect 46777 146085 46811 146113
rect 46839 146085 52259 146113
rect 52287 146085 52321 146113
rect 52349 146085 67619 146113
rect 67647 146085 67681 146113
rect 67709 146085 82979 146113
rect 83007 146085 83041 146113
rect 83069 146085 98339 146113
rect 98367 146085 98401 146113
rect 98429 146085 113699 146113
rect 113727 146085 113761 146113
rect 113789 146085 129059 146113
rect 129087 146085 129121 146113
rect 129149 146085 144419 146113
rect 144447 146085 144481 146113
rect 144509 146085 154625 146113
rect 154653 146085 154687 146113
rect 154715 146085 154749 146113
rect 154777 146085 154811 146113
rect 154839 146085 163625 146113
rect 163653 146085 163687 146113
rect 163715 146085 163749 146113
rect 163777 146085 163811 146113
rect 163839 146085 172625 146113
rect 172653 146085 172687 146113
rect 172715 146085 172749 146113
rect 172777 146085 172811 146113
rect 172839 146085 181625 146113
rect 181653 146085 181687 146113
rect 181715 146085 181749 146113
rect 181777 146085 181811 146113
rect 181839 146085 190625 146113
rect 190653 146085 190687 146113
rect 190715 146085 190749 146113
rect 190777 146085 190811 146113
rect 190839 146085 199625 146113
rect 199653 146085 199687 146113
rect 199715 146085 199749 146113
rect 199777 146085 199811 146113
rect 199839 146085 208625 146113
rect 208653 146085 208687 146113
rect 208715 146085 208749 146113
rect 208777 146085 208811 146113
rect 208839 146085 217625 146113
rect 217653 146085 217687 146113
rect 217715 146085 217749 146113
rect 217777 146085 217811 146113
rect 217839 146085 226625 146113
rect 226653 146085 226687 146113
rect 226715 146085 226749 146113
rect 226777 146085 226811 146113
rect 226839 146085 235625 146113
rect 235653 146085 235687 146113
rect 235715 146085 235749 146113
rect 235777 146085 235811 146113
rect 235839 146085 244625 146113
rect 244653 146085 244687 146113
rect 244715 146085 244749 146113
rect 244777 146085 244811 146113
rect 244839 146085 253625 146113
rect 253653 146085 253687 146113
rect 253715 146085 253749 146113
rect 253777 146085 253811 146113
rect 253839 146085 262625 146113
rect 262653 146085 262687 146113
rect 262715 146085 262749 146113
rect 262777 146085 262811 146113
rect 262839 146085 271625 146113
rect 271653 146085 271687 146113
rect 271715 146085 271749 146113
rect 271777 146085 271811 146113
rect 271839 146085 280625 146113
rect 280653 146085 280687 146113
rect 280715 146085 280749 146113
rect 280777 146085 280811 146113
rect 280839 146085 289625 146113
rect 289653 146085 289687 146113
rect 289715 146085 289749 146113
rect 289777 146085 289811 146113
rect 289839 146085 298248 146113
rect 298276 146085 298310 146113
rect 298338 146085 298372 146113
rect 298400 146085 298434 146113
rect 298462 146085 298990 146113
rect -958 146051 298990 146085
rect -958 146023 -430 146051
rect -402 146023 -368 146051
rect -340 146023 -306 146051
rect -278 146023 -244 146051
rect -216 146023 1625 146051
rect 1653 146023 1687 146051
rect 1715 146023 1749 146051
rect 1777 146023 1811 146051
rect 1839 146023 10625 146051
rect 10653 146023 10687 146051
rect 10715 146023 10749 146051
rect 10777 146023 10811 146051
rect 10839 146023 19625 146051
rect 19653 146023 19687 146051
rect 19715 146023 19749 146051
rect 19777 146023 19811 146051
rect 19839 146023 28625 146051
rect 28653 146023 28687 146051
rect 28715 146023 28749 146051
rect 28777 146023 28811 146051
rect 28839 146023 37625 146051
rect 37653 146023 37687 146051
rect 37715 146023 37749 146051
rect 37777 146023 37811 146051
rect 37839 146023 46625 146051
rect 46653 146023 46687 146051
rect 46715 146023 46749 146051
rect 46777 146023 46811 146051
rect 46839 146023 52259 146051
rect 52287 146023 52321 146051
rect 52349 146023 67619 146051
rect 67647 146023 67681 146051
rect 67709 146023 82979 146051
rect 83007 146023 83041 146051
rect 83069 146023 98339 146051
rect 98367 146023 98401 146051
rect 98429 146023 113699 146051
rect 113727 146023 113761 146051
rect 113789 146023 129059 146051
rect 129087 146023 129121 146051
rect 129149 146023 144419 146051
rect 144447 146023 144481 146051
rect 144509 146023 154625 146051
rect 154653 146023 154687 146051
rect 154715 146023 154749 146051
rect 154777 146023 154811 146051
rect 154839 146023 163625 146051
rect 163653 146023 163687 146051
rect 163715 146023 163749 146051
rect 163777 146023 163811 146051
rect 163839 146023 172625 146051
rect 172653 146023 172687 146051
rect 172715 146023 172749 146051
rect 172777 146023 172811 146051
rect 172839 146023 181625 146051
rect 181653 146023 181687 146051
rect 181715 146023 181749 146051
rect 181777 146023 181811 146051
rect 181839 146023 190625 146051
rect 190653 146023 190687 146051
rect 190715 146023 190749 146051
rect 190777 146023 190811 146051
rect 190839 146023 199625 146051
rect 199653 146023 199687 146051
rect 199715 146023 199749 146051
rect 199777 146023 199811 146051
rect 199839 146023 208625 146051
rect 208653 146023 208687 146051
rect 208715 146023 208749 146051
rect 208777 146023 208811 146051
rect 208839 146023 217625 146051
rect 217653 146023 217687 146051
rect 217715 146023 217749 146051
rect 217777 146023 217811 146051
rect 217839 146023 226625 146051
rect 226653 146023 226687 146051
rect 226715 146023 226749 146051
rect 226777 146023 226811 146051
rect 226839 146023 235625 146051
rect 235653 146023 235687 146051
rect 235715 146023 235749 146051
rect 235777 146023 235811 146051
rect 235839 146023 244625 146051
rect 244653 146023 244687 146051
rect 244715 146023 244749 146051
rect 244777 146023 244811 146051
rect 244839 146023 253625 146051
rect 253653 146023 253687 146051
rect 253715 146023 253749 146051
rect 253777 146023 253811 146051
rect 253839 146023 262625 146051
rect 262653 146023 262687 146051
rect 262715 146023 262749 146051
rect 262777 146023 262811 146051
rect 262839 146023 271625 146051
rect 271653 146023 271687 146051
rect 271715 146023 271749 146051
rect 271777 146023 271811 146051
rect 271839 146023 280625 146051
rect 280653 146023 280687 146051
rect 280715 146023 280749 146051
rect 280777 146023 280811 146051
rect 280839 146023 289625 146051
rect 289653 146023 289687 146051
rect 289715 146023 289749 146051
rect 289777 146023 289811 146051
rect 289839 146023 298248 146051
rect 298276 146023 298310 146051
rect 298338 146023 298372 146051
rect 298400 146023 298434 146051
rect 298462 146023 298990 146051
rect -958 145989 298990 146023
rect -958 145961 -430 145989
rect -402 145961 -368 145989
rect -340 145961 -306 145989
rect -278 145961 -244 145989
rect -216 145961 1625 145989
rect 1653 145961 1687 145989
rect 1715 145961 1749 145989
rect 1777 145961 1811 145989
rect 1839 145961 10625 145989
rect 10653 145961 10687 145989
rect 10715 145961 10749 145989
rect 10777 145961 10811 145989
rect 10839 145961 19625 145989
rect 19653 145961 19687 145989
rect 19715 145961 19749 145989
rect 19777 145961 19811 145989
rect 19839 145961 28625 145989
rect 28653 145961 28687 145989
rect 28715 145961 28749 145989
rect 28777 145961 28811 145989
rect 28839 145961 37625 145989
rect 37653 145961 37687 145989
rect 37715 145961 37749 145989
rect 37777 145961 37811 145989
rect 37839 145961 46625 145989
rect 46653 145961 46687 145989
rect 46715 145961 46749 145989
rect 46777 145961 46811 145989
rect 46839 145961 52259 145989
rect 52287 145961 52321 145989
rect 52349 145961 67619 145989
rect 67647 145961 67681 145989
rect 67709 145961 82979 145989
rect 83007 145961 83041 145989
rect 83069 145961 98339 145989
rect 98367 145961 98401 145989
rect 98429 145961 113699 145989
rect 113727 145961 113761 145989
rect 113789 145961 129059 145989
rect 129087 145961 129121 145989
rect 129149 145961 144419 145989
rect 144447 145961 144481 145989
rect 144509 145961 154625 145989
rect 154653 145961 154687 145989
rect 154715 145961 154749 145989
rect 154777 145961 154811 145989
rect 154839 145961 163625 145989
rect 163653 145961 163687 145989
rect 163715 145961 163749 145989
rect 163777 145961 163811 145989
rect 163839 145961 172625 145989
rect 172653 145961 172687 145989
rect 172715 145961 172749 145989
rect 172777 145961 172811 145989
rect 172839 145961 181625 145989
rect 181653 145961 181687 145989
rect 181715 145961 181749 145989
rect 181777 145961 181811 145989
rect 181839 145961 190625 145989
rect 190653 145961 190687 145989
rect 190715 145961 190749 145989
rect 190777 145961 190811 145989
rect 190839 145961 199625 145989
rect 199653 145961 199687 145989
rect 199715 145961 199749 145989
rect 199777 145961 199811 145989
rect 199839 145961 208625 145989
rect 208653 145961 208687 145989
rect 208715 145961 208749 145989
rect 208777 145961 208811 145989
rect 208839 145961 217625 145989
rect 217653 145961 217687 145989
rect 217715 145961 217749 145989
rect 217777 145961 217811 145989
rect 217839 145961 226625 145989
rect 226653 145961 226687 145989
rect 226715 145961 226749 145989
rect 226777 145961 226811 145989
rect 226839 145961 235625 145989
rect 235653 145961 235687 145989
rect 235715 145961 235749 145989
rect 235777 145961 235811 145989
rect 235839 145961 244625 145989
rect 244653 145961 244687 145989
rect 244715 145961 244749 145989
rect 244777 145961 244811 145989
rect 244839 145961 253625 145989
rect 253653 145961 253687 145989
rect 253715 145961 253749 145989
rect 253777 145961 253811 145989
rect 253839 145961 262625 145989
rect 262653 145961 262687 145989
rect 262715 145961 262749 145989
rect 262777 145961 262811 145989
rect 262839 145961 271625 145989
rect 271653 145961 271687 145989
rect 271715 145961 271749 145989
rect 271777 145961 271811 145989
rect 271839 145961 280625 145989
rect 280653 145961 280687 145989
rect 280715 145961 280749 145989
rect 280777 145961 280811 145989
rect 280839 145961 289625 145989
rect 289653 145961 289687 145989
rect 289715 145961 289749 145989
rect 289777 145961 289811 145989
rect 289839 145961 298248 145989
rect 298276 145961 298310 145989
rect 298338 145961 298372 145989
rect 298400 145961 298434 145989
rect 298462 145961 298990 145989
rect -958 145913 298990 145961
rect -958 140175 298990 140223
rect -958 140147 -910 140175
rect -882 140147 -848 140175
rect -820 140147 -786 140175
rect -758 140147 -724 140175
rect -696 140147 3485 140175
rect 3513 140147 3547 140175
rect 3575 140147 3609 140175
rect 3637 140147 3671 140175
rect 3699 140147 12485 140175
rect 12513 140147 12547 140175
rect 12575 140147 12609 140175
rect 12637 140147 12671 140175
rect 12699 140147 21485 140175
rect 21513 140147 21547 140175
rect 21575 140147 21609 140175
rect 21637 140147 21671 140175
rect 21699 140147 30485 140175
rect 30513 140147 30547 140175
rect 30575 140147 30609 140175
rect 30637 140147 30671 140175
rect 30699 140147 39485 140175
rect 39513 140147 39547 140175
rect 39575 140147 39609 140175
rect 39637 140147 39671 140175
rect 39699 140147 48485 140175
rect 48513 140147 48547 140175
rect 48575 140147 48609 140175
rect 48637 140147 48671 140175
rect 48699 140147 59939 140175
rect 59967 140147 60001 140175
rect 60029 140147 75299 140175
rect 75327 140147 75361 140175
rect 75389 140147 90659 140175
rect 90687 140147 90721 140175
rect 90749 140147 106019 140175
rect 106047 140147 106081 140175
rect 106109 140147 121379 140175
rect 121407 140147 121441 140175
rect 121469 140147 136739 140175
rect 136767 140147 136801 140175
rect 136829 140147 156485 140175
rect 156513 140147 156547 140175
rect 156575 140147 156609 140175
rect 156637 140147 156671 140175
rect 156699 140147 165485 140175
rect 165513 140147 165547 140175
rect 165575 140147 165609 140175
rect 165637 140147 165671 140175
rect 165699 140147 174485 140175
rect 174513 140147 174547 140175
rect 174575 140147 174609 140175
rect 174637 140147 174671 140175
rect 174699 140147 183485 140175
rect 183513 140147 183547 140175
rect 183575 140147 183609 140175
rect 183637 140147 183671 140175
rect 183699 140147 192485 140175
rect 192513 140147 192547 140175
rect 192575 140147 192609 140175
rect 192637 140147 192671 140175
rect 192699 140147 201485 140175
rect 201513 140147 201547 140175
rect 201575 140147 201609 140175
rect 201637 140147 201671 140175
rect 201699 140147 210485 140175
rect 210513 140147 210547 140175
rect 210575 140147 210609 140175
rect 210637 140147 210671 140175
rect 210699 140147 219485 140175
rect 219513 140147 219547 140175
rect 219575 140147 219609 140175
rect 219637 140147 219671 140175
rect 219699 140147 228485 140175
rect 228513 140147 228547 140175
rect 228575 140147 228609 140175
rect 228637 140147 228671 140175
rect 228699 140147 237485 140175
rect 237513 140147 237547 140175
rect 237575 140147 237609 140175
rect 237637 140147 237671 140175
rect 237699 140147 246485 140175
rect 246513 140147 246547 140175
rect 246575 140147 246609 140175
rect 246637 140147 246671 140175
rect 246699 140147 255485 140175
rect 255513 140147 255547 140175
rect 255575 140147 255609 140175
rect 255637 140147 255671 140175
rect 255699 140147 264485 140175
rect 264513 140147 264547 140175
rect 264575 140147 264609 140175
rect 264637 140147 264671 140175
rect 264699 140147 273485 140175
rect 273513 140147 273547 140175
rect 273575 140147 273609 140175
rect 273637 140147 273671 140175
rect 273699 140147 282485 140175
rect 282513 140147 282547 140175
rect 282575 140147 282609 140175
rect 282637 140147 282671 140175
rect 282699 140147 291485 140175
rect 291513 140147 291547 140175
rect 291575 140147 291609 140175
rect 291637 140147 291671 140175
rect 291699 140147 298728 140175
rect 298756 140147 298790 140175
rect 298818 140147 298852 140175
rect 298880 140147 298914 140175
rect 298942 140147 298990 140175
rect -958 140113 298990 140147
rect -958 140085 -910 140113
rect -882 140085 -848 140113
rect -820 140085 -786 140113
rect -758 140085 -724 140113
rect -696 140085 3485 140113
rect 3513 140085 3547 140113
rect 3575 140085 3609 140113
rect 3637 140085 3671 140113
rect 3699 140085 12485 140113
rect 12513 140085 12547 140113
rect 12575 140085 12609 140113
rect 12637 140085 12671 140113
rect 12699 140085 21485 140113
rect 21513 140085 21547 140113
rect 21575 140085 21609 140113
rect 21637 140085 21671 140113
rect 21699 140085 30485 140113
rect 30513 140085 30547 140113
rect 30575 140085 30609 140113
rect 30637 140085 30671 140113
rect 30699 140085 39485 140113
rect 39513 140085 39547 140113
rect 39575 140085 39609 140113
rect 39637 140085 39671 140113
rect 39699 140085 48485 140113
rect 48513 140085 48547 140113
rect 48575 140085 48609 140113
rect 48637 140085 48671 140113
rect 48699 140085 59939 140113
rect 59967 140085 60001 140113
rect 60029 140085 75299 140113
rect 75327 140085 75361 140113
rect 75389 140085 90659 140113
rect 90687 140085 90721 140113
rect 90749 140085 106019 140113
rect 106047 140085 106081 140113
rect 106109 140085 121379 140113
rect 121407 140085 121441 140113
rect 121469 140085 136739 140113
rect 136767 140085 136801 140113
rect 136829 140085 156485 140113
rect 156513 140085 156547 140113
rect 156575 140085 156609 140113
rect 156637 140085 156671 140113
rect 156699 140085 165485 140113
rect 165513 140085 165547 140113
rect 165575 140085 165609 140113
rect 165637 140085 165671 140113
rect 165699 140085 174485 140113
rect 174513 140085 174547 140113
rect 174575 140085 174609 140113
rect 174637 140085 174671 140113
rect 174699 140085 183485 140113
rect 183513 140085 183547 140113
rect 183575 140085 183609 140113
rect 183637 140085 183671 140113
rect 183699 140085 192485 140113
rect 192513 140085 192547 140113
rect 192575 140085 192609 140113
rect 192637 140085 192671 140113
rect 192699 140085 201485 140113
rect 201513 140085 201547 140113
rect 201575 140085 201609 140113
rect 201637 140085 201671 140113
rect 201699 140085 210485 140113
rect 210513 140085 210547 140113
rect 210575 140085 210609 140113
rect 210637 140085 210671 140113
rect 210699 140085 219485 140113
rect 219513 140085 219547 140113
rect 219575 140085 219609 140113
rect 219637 140085 219671 140113
rect 219699 140085 228485 140113
rect 228513 140085 228547 140113
rect 228575 140085 228609 140113
rect 228637 140085 228671 140113
rect 228699 140085 237485 140113
rect 237513 140085 237547 140113
rect 237575 140085 237609 140113
rect 237637 140085 237671 140113
rect 237699 140085 246485 140113
rect 246513 140085 246547 140113
rect 246575 140085 246609 140113
rect 246637 140085 246671 140113
rect 246699 140085 255485 140113
rect 255513 140085 255547 140113
rect 255575 140085 255609 140113
rect 255637 140085 255671 140113
rect 255699 140085 264485 140113
rect 264513 140085 264547 140113
rect 264575 140085 264609 140113
rect 264637 140085 264671 140113
rect 264699 140085 273485 140113
rect 273513 140085 273547 140113
rect 273575 140085 273609 140113
rect 273637 140085 273671 140113
rect 273699 140085 282485 140113
rect 282513 140085 282547 140113
rect 282575 140085 282609 140113
rect 282637 140085 282671 140113
rect 282699 140085 291485 140113
rect 291513 140085 291547 140113
rect 291575 140085 291609 140113
rect 291637 140085 291671 140113
rect 291699 140085 298728 140113
rect 298756 140085 298790 140113
rect 298818 140085 298852 140113
rect 298880 140085 298914 140113
rect 298942 140085 298990 140113
rect -958 140051 298990 140085
rect -958 140023 -910 140051
rect -882 140023 -848 140051
rect -820 140023 -786 140051
rect -758 140023 -724 140051
rect -696 140023 3485 140051
rect 3513 140023 3547 140051
rect 3575 140023 3609 140051
rect 3637 140023 3671 140051
rect 3699 140023 12485 140051
rect 12513 140023 12547 140051
rect 12575 140023 12609 140051
rect 12637 140023 12671 140051
rect 12699 140023 21485 140051
rect 21513 140023 21547 140051
rect 21575 140023 21609 140051
rect 21637 140023 21671 140051
rect 21699 140023 30485 140051
rect 30513 140023 30547 140051
rect 30575 140023 30609 140051
rect 30637 140023 30671 140051
rect 30699 140023 39485 140051
rect 39513 140023 39547 140051
rect 39575 140023 39609 140051
rect 39637 140023 39671 140051
rect 39699 140023 48485 140051
rect 48513 140023 48547 140051
rect 48575 140023 48609 140051
rect 48637 140023 48671 140051
rect 48699 140023 59939 140051
rect 59967 140023 60001 140051
rect 60029 140023 75299 140051
rect 75327 140023 75361 140051
rect 75389 140023 90659 140051
rect 90687 140023 90721 140051
rect 90749 140023 106019 140051
rect 106047 140023 106081 140051
rect 106109 140023 121379 140051
rect 121407 140023 121441 140051
rect 121469 140023 136739 140051
rect 136767 140023 136801 140051
rect 136829 140023 156485 140051
rect 156513 140023 156547 140051
rect 156575 140023 156609 140051
rect 156637 140023 156671 140051
rect 156699 140023 165485 140051
rect 165513 140023 165547 140051
rect 165575 140023 165609 140051
rect 165637 140023 165671 140051
rect 165699 140023 174485 140051
rect 174513 140023 174547 140051
rect 174575 140023 174609 140051
rect 174637 140023 174671 140051
rect 174699 140023 183485 140051
rect 183513 140023 183547 140051
rect 183575 140023 183609 140051
rect 183637 140023 183671 140051
rect 183699 140023 192485 140051
rect 192513 140023 192547 140051
rect 192575 140023 192609 140051
rect 192637 140023 192671 140051
rect 192699 140023 201485 140051
rect 201513 140023 201547 140051
rect 201575 140023 201609 140051
rect 201637 140023 201671 140051
rect 201699 140023 210485 140051
rect 210513 140023 210547 140051
rect 210575 140023 210609 140051
rect 210637 140023 210671 140051
rect 210699 140023 219485 140051
rect 219513 140023 219547 140051
rect 219575 140023 219609 140051
rect 219637 140023 219671 140051
rect 219699 140023 228485 140051
rect 228513 140023 228547 140051
rect 228575 140023 228609 140051
rect 228637 140023 228671 140051
rect 228699 140023 237485 140051
rect 237513 140023 237547 140051
rect 237575 140023 237609 140051
rect 237637 140023 237671 140051
rect 237699 140023 246485 140051
rect 246513 140023 246547 140051
rect 246575 140023 246609 140051
rect 246637 140023 246671 140051
rect 246699 140023 255485 140051
rect 255513 140023 255547 140051
rect 255575 140023 255609 140051
rect 255637 140023 255671 140051
rect 255699 140023 264485 140051
rect 264513 140023 264547 140051
rect 264575 140023 264609 140051
rect 264637 140023 264671 140051
rect 264699 140023 273485 140051
rect 273513 140023 273547 140051
rect 273575 140023 273609 140051
rect 273637 140023 273671 140051
rect 273699 140023 282485 140051
rect 282513 140023 282547 140051
rect 282575 140023 282609 140051
rect 282637 140023 282671 140051
rect 282699 140023 291485 140051
rect 291513 140023 291547 140051
rect 291575 140023 291609 140051
rect 291637 140023 291671 140051
rect 291699 140023 298728 140051
rect 298756 140023 298790 140051
rect 298818 140023 298852 140051
rect 298880 140023 298914 140051
rect 298942 140023 298990 140051
rect -958 139989 298990 140023
rect -958 139961 -910 139989
rect -882 139961 -848 139989
rect -820 139961 -786 139989
rect -758 139961 -724 139989
rect -696 139961 3485 139989
rect 3513 139961 3547 139989
rect 3575 139961 3609 139989
rect 3637 139961 3671 139989
rect 3699 139961 12485 139989
rect 12513 139961 12547 139989
rect 12575 139961 12609 139989
rect 12637 139961 12671 139989
rect 12699 139961 21485 139989
rect 21513 139961 21547 139989
rect 21575 139961 21609 139989
rect 21637 139961 21671 139989
rect 21699 139961 30485 139989
rect 30513 139961 30547 139989
rect 30575 139961 30609 139989
rect 30637 139961 30671 139989
rect 30699 139961 39485 139989
rect 39513 139961 39547 139989
rect 39575 139961 39609 139989
rect 39637 139961 39671 139989
rect 39699 139961 48485 139989
rect 48513 139961 48547 139989
rect 48575 139961 48609 139989
rect 48637 139961 48671 139989
rect 48699 139961 59939 139989
rect 59967 139961 60001 139989
rect 60029 139961 75299 139989
rect 75327 139961 75361 139989
rect 75389 139961 90659 139989
rect 90687 139961 90721 139989
rect 90749 139961 106019 139989
rect 106047 139961 106081 139989
rect 106109 139961 121379 139989
rect 121407 139961 121441 139989
rect 121469 139961 136739 139989
rect 136767 139961 136801 139989
rect 136829 139961 156485 139989
rect 156513 139961 156547 139989
rect 156575 139961 156609 139989
rect 156637 139961 156671 139989
rect 156699 139961 165485 139989
rect 165513 139961 165547 139989
rect 165575 139961 165609 139989
rect 165637 139961 165671 139989
rect 165699 139961 174485 139989
rect 174513 139961 174547 139989
rect 174575 139961 174609 139989
rect 174637 139961 174671 139989
rect 174699 139961 183485 139989
rect 183513 139961 183547 139989
rect 183575 139961 183609 139989
rect 183637 139961 183671 139989
rect 183699 139961 192485 139989
rect 192513 139961 192547 139989
rect 192575 139961 192609 139989
rect 192637 139961 192671 139989
rect 192699 139961 201485 139989
rect 201513 139961 201547 139989
rect 201575 139961 201609 139989
rect 201637 139961 201671 139989
rect 201699 139961 210485 139989
rect 210513 139961 210547 139989
rect 210575 139961 210609 139989
rect 210637 139961 210671 139989
rect 210699 139961 219485 139989
rect 219513 139961 219547 139989
rect 219575 139961 219609 139989
rect 219637 139961 219671 139989
rect 219699 139961 228485 139989
rect 228513 139961 228547 139989
rect 228575 139961 228609 139989
rect 228637 139961 228671 139989
rect 228699 139961 237485 139989
rect 237513 139961 237547 139989
rect 237575 139961 237609 139989
rect 237637 139961 237671 139989
rect 237699 139961 246485 139989
rect 246513 139961 246547 139989
rect 246575 139961 246609 139989
rect 246637 139961 246671 139989
rect 246699 139961 255485 139989
rect 255513 139961 255547 139989
rect 255575 139961 255609 139989
rect 255637 139961 255671 139989
rect 255699 139961 264485 139989
rect 264513 139961 264547 139989
rect 264575 139961 264609 139989
rect 264637 139961 264671 139989
rect 264699 139961 273485 139989
rect 273513 139961 273547 139989
rect 273575 139961 273609 139989
rect 273637 139961 273671 139989
rect 273699 139961 282485 139989
rect 282513 139961 282547 139989
rect 282575 139961 282609 139989
rect 282637 139961 282671 139989
rect 282699 139961 291485 139989
rect 291513 139961 291547 139989
rect 291575 139961 291609 139989
rect 291637 139961 291671 139989
rect 291699 139961 298728 139989
rect 298756 139961 298790 139989
rect 298818 139961 298852 139989
rect 298880 139961 298914 139989
rect 298942 139961 298990 139989
rect -958 139913 298990 139961
rect -958 137175 298990 137223
rect -958 137147 -430 137175
rect -402 137147 -368 137175
rect -340 137147 -306 137175
rect -278 137147 -244 137175
rect -216 137147 1625 137175
rect 1653 137147 1687 137175
rect 1715 137147 1749 137175
rect 1777 137147 1811 137175
rect 1839 137147 10625 137175
rect 10653 137147 10687 137175
rect 10715 137147 10749 137175
rect 10777 137147 10811 137175
rect 10839 137147 19625 137175
rect 19653 137147 19687 137175
rect 19715 137147 19749 137175
rect 19777 137147 19811 137175
rect 19839 137147 28625 137175
rect 28653 137147 28687 137175
rect 28715 137147 28749 137175
rect 28777 137147 28811 137175
rect 28839 137147 37625 137175
rect 37653 137147 37687 137175
rect 37715 137147 37749 137175
rect 37777 137147 37811 137175
rect 37839 137147 46625 137175
rect 46653 137147 46687 137175
rect 46715 137147 46749 137175
rect 46777 137147 46811 137175
rect 46839 137147 52259 137175
rect 52287 137147 52321 137175
rect 52349 137147 67619 137175
rect 67647 137147 67681 137175
rect 67709 137147 82979 137175
rect 83007 137147 83041 137175
rect 83069 137147 98339 137175
rect 98367 137147 98401 137175
rect 98429 137147 113699 137175
rect 113727 137147 113761 137175
rect 113789 137147 129059 137175
rect 129087 137147 129121 137175
rect 129149 137147 144419 137175
rect 144447 137147 144481 137175
rect 144509 137147 154625 137175
rect 154653 137147 154687 137175
rect 154715 137147 154749 137175
rect 154777 137147 154811 137175
rect 154839 137147 163625 137175
rect 163653 137147 163687 137175
rect 163715 137147 163749 137175
rect 163777 137147 163811 137175
rect 163839 137147 172625 137175
rect 172653 137147 172687 137175
rect 172715 137147 172749 137175
rect 172777 137147 172811 137175
rect 172839 137147 181625 137175
rect 181653 137147 181687 137175
rect 181715 137147 181749 137175
rect 181777 137147 181811 137175
rect 181839 137147 190625 137175
rect 190653 137147 190687 137175
rect 190715 137147 190749 137175
rect 190777 137147 190811 137175
rect 190839 137147 199625 137175
rect 199653 137147 199687 137175
rect 199715 137147 199749 137175
rect 199777 137147 199811 137175
rect 199839 137147 208625 137175
rect 208653 137147 208687 137175
rect 208715 137147 208749 137175
rect 208777 137147 208811 137175
rect 208839 137147 217625 137175
rect 217653 137147 217687 137175
rect 217715 137147 217749 137175
rect 217777 137147 217811 137175
rect 217839 137147 226625 137175
rect 226653 137147 226687 137175
rect 226715 137147 226749 137175
rect 226777 137147 226811 137175
rect 226839 137147 235625 137175
rect 235653 137147 235687 137175
rect 235715 137147 235749 137175
rect 235777 137147 235811 137175
rect 235839 137147 244625 137175
rect 244653 137147 244687 137175
rect 244715 137147 244749 137175
rect 244777 137147 244811 137175
rect 244839 137147 253625 137175
rect 253653 137147 253687 137175
rect 253715 137147 253749 137175
rect 253777 137147 253811 137175
rect 253839 137147 262625 137175
rect 262653 137147 262687 137175
rect 262715 137147 262749 137175
rect 262777 137147 262811 137175
rect 262839 137147 271625 137175
rect 271653 137147 271687 137175
rect 271715 137147 271749 137175
rect 271777 137147 271811 137175
rect 271839 137147 280625 137175
rect 280653 137147 280687 137175
rect 280715 137147 280749 137175
rect 280777 137147 280811 137175
rect 280839 137147 289625 137175
rect 289653 137147 289687 137175
rect 289715 137147 289749 137175
rect 289777 137147 289811 137175
rect 289839 137147 298248 137175
rect 298276 137147 298310 137175
rect 298338 137147 298372 137175
rect 298400 137147 298434 137175
rect 298462 137147 298990 137175
rect -958 137113 298990 137147
rect -958 137085 -430 137113
rect -402 137085 -368 137113
rect -340 137085 -306 137113
rect -278 137085 -244 137113
rect -216 137085 1625 137113
rect 1653 137085 1687 137113
rect 1715 137085 1749 137113
rect 1777 137085 1811 137113
rect 1839 137085 10625 137113
rect 10653 137085 10687 137113
rect 10715 137085 10749 137113
rect 10777 137085 10811 137113
rect 10839 137085 19625 137113
rect 19653 137085 19687 137113
rect 19715 137085 19749 137113
rect 19777 137085 19811 137113
rect 19839 137085 28625 137113
rect 28653 137085 28687 137113
rect 28715 137085 28749 137113
rect 28777 137085 28811 137113
rect 28839 137085 37625 137113
rect 37653 137085 37687 137113
rect 37715 137085 37749 137113
rect 37777 137085 37811 137113
rect 37839 137085 46625 137113
rect 46653 137085 46687 137113
rect 46715 137085 46749 137113
rect 46777 137085 46811 137113
rect 46839 137085 52259 137113
rect 52287 137085 52321 137113
rect 52349 137085 67619 137113
rect 67647 137085 67681 137113
rect 67709 137085 82979 137113
rect 83007 137085 83041 137113
rect 83069 137085 98339 137113
rect 98367 137085 98401 137113
rect 98429 137085 113699 137113
rect 113727 137085 113761 137113
rect 113789 137085 129059 137113
rect 129087 137085 129121 137113
rect 129149 137085 144419 137113
rect 144447 137085 144481 137113
rect 144509 137085 154625 137113
rect 154653 137085 154687 137113
rect 154715 137085 154749 137113
rect 154777 137085 154811 137113
rect 154839 137085 163625 137113
rect 163653 137085 163687 137113
rect 163715 137085 163749 137113
rect 163777 137085 163811 137113
rect 163839 137085 172625 137113
rect 172653 137085 172687 137113
rect 172715 137085 172749 137113
rect 172777 137085 172811 137113
rect 172839 137085 181625 137113
rect 181653 137085 181687 137113
rect 181715 137085 181749 137113
rect 181777 137085 181811 137113
rect 181839 137085 190625 137113
rect 190653 137085 190687 137113
rect 190715 137085 190749 137113
rect 190777 137085 190811 137113
rect 190839 137085 199625 137113
rect 199653 137085 199687 137113
rect 199715 137085 199749 137113
rect 199777 137085 199811 137113
rect 199839 137085 208625 137113
rect 208653 137085 208687 137113
rect 208715 137085 208749 137113
rect 208777 137085 208811 137113
rect 208839 137085 217625 137113
rect 217653 137085 217687 137113
rect 217715 137085 217749 137113
rect 217777 137085 217811 137113
rect 217839 137085 226625 137113
rect 226653 137085 226687 137113
rect 226715 137085 226749 137113
rect 226777 137085 226811 137113
rect 226839 137085 235625 137113
rect 235653 137085 235687 137113
rect 235715 137085 235749 137113
rect 235777 137085 235811 137113
rect 235839 137085 244625 137113
rect 244653 137085 244687 137113
rect 244715 137085 244749 137113
rect 244777 137085 244811 137113
rect 244839 137085 253625 137113
rect 253653 137085 253687 137113
rect 253715 137085 253749 137113
rect 253777 137085 253811 137113
rect 253839 137085 262625 137113
rect 262653 137085 262687 137113
rect 262715 137085 262749 137113
rect 262777 137085 262811 137113
rect 262839 137085 271625 137113
rect 271653 137085 271687 137113
rect 271715 137085 271749 137113
rect 271777 137085 271811 137113
rect 271839 137085 280625 137113
rect 280653 137085 280687 137113
rect 280715 137085 280749 137113
rect 280777 137085 280811 137113
rect 280839 137085 289625 137113
rect 289653 137085 289687 137113
rect 289715 137085 289749 137113
rect 289777 137085 289811 137113
rect 289839 137085 298248 137113
rect 298276 137085 298310 137113
rect 298338 137085 298372 137113
rect 298400 137085 298434 137113
rect 298462 137085 298990 137113
rect -958 137051 298990 137085
rect -958 137023 -430 137051
rect -402 137023 -368 137051
rect -340 137023 -306 137051
rect -278 137023 -244 137051
rect -216 137023 1625 137051
rect 1653 137023 1687 137051
rect 1715 137023 1749 137051
rect 1777 137023 1811 137051
rect 1839 137023 10625 137051
rect 10653 137023 10687 137051
rect 10715 137023 10749 137051
rect 10777 137023 10811 137051
rect 10839 137023 19625 137051
rect 19653 137023 19687 137051
rect 19715 137023 19749 137051
rect 19777 137023 19811 137051
rect 19839 137023 28625 137051
rect 28653 137023 28687 137051
rect 28715 137023 28749 137051
rect 28777 137023 28811 137051
rect 28839 137023 37625 137051
rect 37653 137023 37687 137051
rect 37715 137023 37749 137051
rect 37777 137023 37811 137051
rect 37839 137023 46625 137051
rect 46653 137023 46687 137051
rect 46715 137023 46749 137051
rect 46777 137023 46811 137051
rect 46839 137023 52259 137051
rect 52287 137023 52321 137051
rect 52349 137023 67619 137051
rect 67647 137023 67681 137051
rect 67709 137023 82979 137051
rect 83007 137023 83041 137051
rect 83069 137023 98339 137051
rect 98367 137023 98401 137051
rect 98429 137023 113699 137051
rect 113727 137023 113761 137051
rect 113789 137023 129059 137051
rect 129087 137023 129121 137051
rect 129149 137023 144419 137051
rect 144447 137023 144481 137051
rect 144509 137023 154625 137051
rect 154653 137023 154687 137051
rect 154715 137023 154749 137051
rect 154777 137023 154811 137051
rect 154839 137023 163625 137051
rect 163653 137023 163687 137051
rect 163715 137023 163749 137051
rect 163777 137023 163811 137051
rect 163839 137023 172625 137051
rect 172653 137023 172687 137051
rect 172715 137023 172749 137051
rect 172777 137023 172811 137051
rect 172839 137023 181625 137051
rect 181653 137023 181687 137051
rect 181715 137023 181749 137051
rect 181777 137023 181811 137051
rect 181839 137023 190625 137051
rect 190653 137023 190687 137051
rect 190715 137023 190749 137051
rect 190777 137023 190811 137051
rect 190839 137023 199625 137051
rect 199653 137023 199687 137051
rect 199715 137023 199749 137051
rect 199777 137023 199811 137051
rect 199839 137023 208625 137051
rect 208653 137023 208687 137051
rect 208715 137023 208749 137051
rect 208777 137023 208811 137051
rect 208839 137023 217625 137051
rect 217653 137023 217687 137051
rect 217715 137023 217749 137051
rect 217777 137023 217811 137051
rect 217839 137023 226625 137051
rect 226653 137023 226687 137051
rect 226715 137023 226749 137051
rect 226777 137023 226811 137051
rect 226839 137023 235625 137051
rect 235653 137023 235687 137051
rect 235715 137023 235749 137051
rect 235777 137023 235811 137051
rect 235839 137023 244625 137051
rect 244653 137023 244687 137051
rect 244715 137023 244749 137051
rect 244777 137023 244811 137051
rect 244839 137023 253625 137051
rect 253653 137023 253687 137051
rect 253715 137023 253749 137051
rect 253777 137023 253811 137051
rect 253839 137023 262625 137051
rect 262653 137023 262687 137051
rect 262715 137023 262749 137051
rect 262777 137023 262811 137051
rect 262839 137023 271625 137051
rect 271653 137023 271687 137051
rect 271715 137023 271749 137051
rect 271777 137023 271811 137051
rect 271839 137023 280625 137051
rect 280653 137023 280687 137051
rect 280715 137023 280749 137051
rect 280777 137023 280811 137051
rect 280839 137023 289625 137051
rect 289653 137023 289687 137051
rect 289715 137023 289749 137051
rect 289777 137023 289811 137051
rect 289839 137023 298248 137051
rect 298276 137023 298310 137051
rect 298338 137023 298372 137051
rect 298400 137023 298434 137051
rect 298462 137023 298990 137051
rect -958 136989 298990 137023
rect -958 136961 -430 136989
rect -402 136961 -368 136989
rect -340 136961 -306 136989
rect -278 136961 -244 136989
rect -216 136961 1625 136989
rect 1653 136961 1687 136989
rect 1715 136961 1749 136989
rect 1777 136961 1811 136989
rect 1839 136961 10625 136989
rect 10653 136961 10687 136989
rect 10715 136961 10749 136989
rect 10777 136961 10811 136989
rect 10839 136961 19625 136989
rect 19653 136961 19687 136989
rect 19715 136961 19749 136989
rect 19777 136961 19811 136989
rect 19839 136961 28625 136989
rect 28653 136961 28687 136989
rect 28715 136961 28749 136989
rect 28777 136961 28811 136989
rect 28839 136961 37625 136989
rect 37653 136961 37687 136989
rect 37715 136961 37749 136989
rect 37777 136961 37811 136989
rect 37839 136961 46625 136989
rect 46653 136961 46687 136989
rect 46715 136961 46749 136989
rect 46777 136961 46811 136989
rect 46839 136961 52259 136989
rect 52287 136961 52321 136989
rect 52349 136961 67619 136989
rect 67647 136961 67681 136989
rect 67709 136961 82979 136989
rect 83007 136961 83041 136989
rect 83069 136961 98339 136989
rect 98367 136961 98401 136989
rect 98429 136961 113699 136989
rect 113727 136961 113761 136989
rect 113789 136961 129059 136989
rect 129087 136961 129121 136989
rect 129149 136961 144419 136989
rect 144447 136961 144481 136989
rect 144509 136961 154625 136989
rect 154653 136961 154687 136989
rect 154715 136961 154749 136989
rect 154777 136961 154811 136989
rect 154839 136961 163625 136989
rect 163653 136961 163687 136989
rect 163715 136961 163749 136989
rect 163777 136961 163811 136989
rect 163839 136961 172625 136989
rect 172653 136961 172687 136989
rect 172715 136961 172749 136989
rect 172777 136961 172811 136989
rect 172839 136961 181625 136989
rect 181653 136961 181687 136989
rect 181715 136961 181749 136989
rect 181777 136961 181811 136989
rect 181839 136961 190625 136989
rect 190653 136961 190687 136989
rect 190715 136961 190749 136989
rect 190777 136961 190811 136989
rect 190839 136961 199625 136989
rect 199653 136961 199687 136989
rect 199715 136961 199749 136989
rect 199777 136961 199811 136989
rect 199839 136961 208625 136989
rect 208653 136961 208687 136989
rect 208715 136961 208749 136989
rect 208777 136961 208811 136989
rect 208839 136961 217625 136989
rect 217653 136961 217687 136989
rect 217715 136961 217749 136989
rect 217777 136961 217811 136989
rect 217839 136961 226625 136989
rect 226653 136961 226687 136989
rect 226715 136961 226749 136989
rect 226777 136961 226811 136989
rect 226839 136961 235625 136989
rect 235653 136961 235687 136989
rect 235715 136961 235749 136989
rect 235777 136961 235811 136989
rect 235839 136961 244625 136989
rect 244653 136961 244687 136989
rect 244715 136961 244749 136989
rect 244777 136961 244811 136989
rect 244839 136961 253625 136989
rect 253653 136961 253687 136989
rect 253715 136961 253749 136989
rect 253777 136961 253811 136989
rect 253839 136961 262625 136989
rect 262653 136961 262687 136989
rect 262715 136961 262749 136989
rect 262777 136961 262811 136989
rect 262839 136961 271625 136989
rect 271653 136961 271687 136989
rect 271715 136961 271749 136989
rect 271777 136961 271811 136989
rect 271839 136961 280625 136989
rect 280653 136961 280687 136989
rect 280715 136961 280749 136989
rect 280777 136961 280811 136989
rect 280839 136961 289625 136989
rect 289653 136961 289687 136989
rect 289715 136961 289749 136989
rect 289777 136961 289811 136989
rect 289839 136961 298248 136989
rect 298276 136961 298310 136989
rect 298338 136961 298372 136989
rect 298400 136961 298434 136989
rect 298462 136961 298990 136989
rect -958 136913 298990 136961
rect -958 131175 298990 131223
rect -958 131147 -910 131175
rect -882 131147 -848 131175
rect -820 131147 -786 131175
rect -758 131147 -724 131175
rect -696 131147 3485 131175
rect 3513 131147 3547 131175
rect 3575 131147 3609 131175
rect 3637 131147 3671 131175
rect 3699 131147 12485 131175
rect 12513 131147 12547 131175
rect 12575 131147 12609 131175
rect 12637 131147 12671 131175
rect 12699 131147 21485 131175
rect 21513 131147 21547 131175
rect 21575 131147 21609 131175
rect 21637 131147 21671 131175
rect 21699 131147 30485 131175
rect 30513 131147 30547 131175
rect 30575 131147 30609 131175
rect 30637 131147 30671 131175
rect 30699 131147 39485 131175
rect 39513 131147 39547 131175
rect 39575 131147 39609 131175
rect 39637 131147 39671 131175
rect 39699 131147 48485 131175
rect 48513 131147 48547 131175
rect 48575 131147 48609 131175
rect 48637 131147 48671 131175
rect 48699 131147 59939 131175
rect 59967 131147 60001 131175
rect 60029 131147 75299 131175
rect 75327 131147 75361 131175
rect 75389 131147 90659 131175
rect 90687 131147 90721 131175
rect 90749 131147 106019 131175
rect 106047 131147 106081 131175
rect 106109 131147 121379 131175
rect 121407 131147 121441 131175
rect 121469 131147 136739 131175
rect 136767 131147 136801 131175
rect 136829 131147 156485 131175
rect 156513 131147 156547 131175
rect 156575 131147 156609 131175
rect 156637 131147 156671 131175
rect 156699 131147 165485 131175
rect 165513 131147 165547 131175
rect 165575 131147 165609 131175
rect 165637 131147 165671 131175
rect 165699 131147 174485 131175
rect 174513 131147 174547 131175
rect 174575 131147 174609 131175
rect 174637 131147 174671 131175
rect 174699 131147 183485 131175
rect 183513 131147 183547 131175
rect 183575 131147 183609 131175
rect 183637 131147 183671 131175
rect 183699 131147 192485 131175
rect 192513 131147 192547 131175
rect 192575 131147 192609 131175
rect 192637 131147 192671 131175
rect 192699 131147 201485 131175
rect 201513 131147 201547 131175
rect 201575 131147 201609 131175
rect 201637 131147 201671 131175
rect 201699 131147 210485 131175
rect 210513 131147 210547 131175
rect 210575 131147 210609 131175
rect 210637 131147 210671 131175
rect 210699 131147 219485 131175
rect 219513 131147 219547 131175
rect 219575 131147 219609 131175
rect 219637 131147 219671 131175
rect 219699 131147 228485 131175
rect 228513 131147 228547 131175
rect 228575 131147 228609 131175
rect 228637 131147 228671 131175
rect 228699 131147 237485 131175
rect 237513 131147 237547 131175
rect 237575 131147 237609 131175
rect 237637 131147 237671 131175
rect 237699 131147 246485 131175
rect 246513 131147 246547 131175
rect 246575 131147 246609 131175
rect 246637 131147 246671 131175
rect 246699 131147 255485 131175
rect 255513 131147 255547 131175
rect 255575 131147 255609 131175
rect 255637 131147 255671 131175
rect 255699 131147 264485 131175
rect 264513 131147 264547 131175
rect 264575 131147 264609 131175
rect 264637 131147 264671 131175
rect 264699 131147 273485 131175
rect 273513 131147 273547 131175
rect 273575 131147 273609 131175
rect 273637 131147 273671 131175
rect 273699 131147 282485 131175
rect 282513 131147 282547 131175
rect 282575 131147 282609 131175
rect 282637 131147 282671 131175
rect 282699 131147 291485 131175
rect 291513 131147 291547 131175
rect 291575 131147 291609 131175
rect 291637 131147 291671 131175
rect 291699 131147 298728 131175
rect 298756 131147 298790 131175
rect 298818 131147 298852 131175
rect 298880 131147 298914 131175
rect 298942 131147 298990 131175
rect -958 131113 298990 131147
rect -958 131085 -910 131113
rect -882 131085 -848 131113
rect -820 131085 -786 131113
rect -758 131085 -724 131113
rect -696 131085 3485 131113
rect 3513 131085 3547 131113
rect 3575 131085 3609 131113
rect 3637 131085 3671 131113
rect 3699 131085 12485 131113
rect 12513 131085 12547 131113
rect 12575 131085 12609 131113
rect 12637 131085 12671 131113
rect 12699 131085 21485 131113
rect 21513 131085 21547 131113
rect 21575 131085 21609 131113
rect 21637 131085 21671 131113
rect 21699 131085 30485 131113
rect 30513 131085 30547 131113
rect 30575 131085 30609 131113
rect 30637 131085 30671 131113
rect 30699 131085 39485 131113
rect 39513 131085 39547 131113
rect 39575 131085 39609 131113
rect 39637 131085 39671 131113
rect 39699 131085 48485 131113
rect 48513 131085 48547 131113
rect 48575 131085 48609 131113
rect 48637 131085 48671 131113
rect 48699 131085 59939 131113
rect 59967 131085 60001 131113
rect 60029 131085 75299 131113
rect 75327 131085 75361 131113
rect 75389 131085 90659 131113
rect 90687 131085 90721 131113
rect 90749 131085 106019 131113
rect 106047 131085 106081 131113
rect 106109 131085 121379 131113
rect 121407 131085 121441 131113
rect 121469 131085 136739 131113
rect 136767 131085 136801 131113
rect 136829 131085 156485 131113
rect 156513 131085 156547 131113
rect 156575 131085 156609 131113
rect 156637 131085 156671 131113
rect 156699 131085 165485 131113
rect 165513 131085 165547 131113
rect 165575 131085 165609 131113
rect 165637 131085 165671 131113
rect 165699 131085 174485 131113
rect 174513 131085 174547 131113
rect 174575 131085 174609 131113
rect 174637 131085 174671 131113
rect 174699 131085 183485 131113
rect 183513 131085 183547 131113
rect 183575 131085 183609 131113
rect 183637 131085 183671 131113
rect 183699 131085 192485 131113
rect 192513 131085 192547 131113
rect 192575 131085 192609 131113
rect 192637 131085 192671 131113
rect 192699 131085 201485 131113
rect 201513 131085 201547 131113
rect 201575 131085 201609 131113
rect 201637 131085 201671 131113
rect 201699 131085 210485 131113
rect 210513 131085 210547 131113
rect 210575 131085 210609 131113
rect 210637 131085 210671 131113
rect 210699 131085 219485 131113
rect 219513 131085 219547 131113
rect 219575 131085 219609 131113
rect 219637 131085 219671 131113
rect 219699 131085 228485 131113
rect 228513 131085 228547 131113
rect 228575 131085 228609 131113
rect 228637 131085 228671 131113
rect 228699 131085 237485 131113
rect 237513 131085 237547 131113
rect 237575 131085 237609 131113
rect 237637 131085 237671 131113
rect 237699 131085 246485 131113
rect 246513 131085 246547 131113
rect 246575 131085 246609 131113
rect 246637 131085 246671 131113
rect 246699 131085 255485 131113
rect 255513 131085 255547 131113
rect 255575 131085 255609 131113
rect 255637 131085 255671 131113
rect 255699 131085 264485 131113
rect 264513 131085 264547 131113
rect 264575 131085 264609 131113
rect 264637 131085 264671 131113
rect 264699 131085 273485 131113
rect 273513 131085 273547 131113
rect 273575 131085 273609 131113
rect 273637 131085 273671 131113
rect 273699 131085 282485 131113
rect 282513 131085 282547 131113
rect 282575 131085 282609 131113
rect 282637 131085 282671 131113
rect 282699 131085 291485 131113
rect 291513 131085 291547 131113
rect 291575 131085 291609 131113
rect 291637 131085 291671 131113
rect 291699 131085 298728 131113
rect 298756 131085 298790 131113
rect 298818 131085 298852 131113
rect 298880 131085 298914 131113
rect 298942 131085 298990 131113
rect -958 131051 298990 131085
rect -958 131023 -910 131051
rect -882 131023 -848 131051
rect -820 131023 -786 131051
rect -758 131023 -724 131051
rect -696 131023 3485 131051
rect 3513 131023 3547 131051
rect 3575 131023 3609 131051
rect 3637 131023 3671 131051
rect 3699 131023 12485 131051
rect 12513 131023 12547 131051
rect 12575 131023 12609 131051
rect 12637 131023 12671 131051
rect 12699 131023 21485 131051
rect 21513 131023 21547 131051
rect 21575 131023 21609 131051
rect 21637 131023 21671 131051
rect 21699 131023 30485 131051
rect 30513 131023 30547 131051
rect 30575 131023 30609 131051
rect 30637 131023 30671 131051
rect 30699 131023 39485 131051
rect 39513 131023 39547 131051
rect 39575 131023 39609 131051
rect 39637 131023 39671 131051
rect 39699 131023 48485 131051
rect 48513 131023 48547 131051
rect 48575 131023 48609 131051
rect 48637 131023 48671 131051
rect 48699 131023 59939 131051
rect 59967 131023 60001 131051
rect 60029 131023 75299 131051
rect 75327 131023 75361 131051
rect 75389 131023 90659 131051
rect 90687 131023 90721 131051
rect 90749 131023 106019 131051
rect 106047 131023 106081 131051
rect 106109 131023 121379 131051
rect 121407 131023 121441 131051
rect 121469 131023 136739 131051
rect 136767 131023 136801 131051
rect 136829 131023 156485 131051
rect 156513 131023 156547 131051
rect 156575 131023 156609 131051
rect 156637 131023 156671 131051
rect 156699 131023 165485 131051
rect 165513 131023 165547 131051
rect 165575 131023 165609 131051
rect 165637 131023 165671 131051
rect 165699 131023 174485 131051
rect 174513 131023 174547 131051
rect 174575 131023 174609 131051
rect 174637 131023 174671 131051
rect 174699 131023 183485 131051
rect 183513 131023 183547 131051
rect 183575 131023 183609 131051
rect 183637 131023 183671 131051
rect 183699 131023 192485 131051
rect 192513 131023 192547 131051
rect 192575 131023 192609 131051
rect 192637 131023 192671 131051
rect 192699 131023 201485 131051
rect 201513 131023 201547 131051
rect 201575 131023 201609 131051
rect 201637 131023 201671 131051
rect 201699 131023 210485 131051
rect 210513 131023 210547 131051
rect 210575 131023 210609 131051
rect 210637 131023 210671 131051
rect 210699 131023 219485 131051
rect 219513 131023 219547 131051
rect 219575 131023 219609 131051
rect 219637 131023 219671 131051
rect 219699 131023 228485 131051
rect 228513 131023 228547 131051
rect 228575 131023 228609 131051
rect 228637 131023 228671 131051
rect 228699 131023 237485 131051
rect 237513 131023 237547 131051
rect 237575 131023 237609 131051
rect 237637 131023 237671 131051
rect 237699 131023 246485 131051
rect 246513 131023 246547 131051
rect 246575 131023 246609 131051
rect 246637 131023 246671 131051
rect 246699 131023 255485 131051
rect 255513 131023 255547 131051
rect 255575 131023 255609 131051
rect 255637 131023 255671 131051
rect 255699 131023 264485 131051
rect 264513 131023 264547 131051
rect 264575 131023 264609 131051
rect 264637 131023 264671 131051
rect 264699 131023 273485 131051
rect 273513 131023 273547 131051
rect 273575 131023 273609 131051
rect 273637 131023 273671 131051
rect 273699 131023 282485 131051
rect 282513 131023 282547 131051
rect 282575 131023 282609 131051
rect 282637 131023 282671 131051
rect 282699 131023 291485 131051
rect 291513 131023 291547 131051
rect 291575 131023 291609 131051
rect 291637 131023 291671 131051
rect 291699 131023 298728 131051
rect 298756 131023 298790 131051
rect 298818 131023 298852 131051
rect 298880 131023 298914 131051
rect 298942 131023 298990 131051
rect -958 130989 298990 131023
rect -958 130961 -910 130989
rect -882 130961 -848 130989
rect -820 130961 -786 130989
rect -758 130961 -724 130989
rect -696 130961 3485 130989
rect 3513 130961 3547 130989
rect 3575 130961 3609 130989
rect 3637 130961 3671 130989
rect 3699 130961 12485 130989
rect 12513 130961 12547 130989
rect 12575 130961 12609 130989
rect 12637 130961 12671 130989
rect 12699 130961 21485 130989
rect 21513 130961 21547 130989
rect 21575 130961 21609 130989
rect 21637 130961 21671 130989
rect 21699 130961 30485 130989
rect 30513 130961 30547 130989
rect 30575 130961 30609 130989
rect 30637 130961 30671 130989
rect 30699 130961 39485 130989
rect 39513 130961 39547 130989
rect 39575 130961 39609 130989
rect 39637 130961 39671 130989
rect 39699 130961 48485 130989
rect 48513 130961 48547 130989
rect 48575 130961 48609 130989
rect 48637 130961 48671 130989
rect 48699 130961 59939 130989
rect 59967 130961 60001 130989
rect 60029 130961 75299 130989
rect 75327 130961 75361 130989
rect 75389 130961 90659 130989
rect 90687 130961 90721 130989
rect 90749 130961 106019 130989
rect 106047 130961 106081 130989
rect 106109 130961 121379 130989
rect 121407 130961 121441 130989
rect 121469 130961 136739 130989
rect 136767 130961 136801 130989
rect 136829 130961 156485 130989
rect 156513 130961 156547 130989
rect 156575 130961 156609 130989
rect 156637 130961 156671 130989
rect 156699 130961 165485 130989
rect 165513 130961 165547 130989
rect 165575 130961 165609 130989
rect 165637 130961 165671 130989
rect 165699 130961 174485 130989
rect 174513 130961 174547 130989
rect 174575 130961 174609 130989
rect 174637 130961 174671 130989
rect 174699 130961 183485 130989
rect 183513 130961 183547 130989
rect 183575 130961 183609 130989
rect 183637 130961 183671 130989
rect 183699 130961 192485 130989
rect 192513 130961 192547 130989
rect 192575 130961 192609 130989
rect 192637 130961 192671 130989
rect 192699 130961 201485 130989
rect 201513 130961 201547 130989
rect 201575 130961 201609 130989
rect 201637 130961 201671 130989
rect 201699 130961 210485 130989
rect 210513 130961 210547 130989
rect 210575 130961 210609 130989
rect 210637 130961 210671 130989
rect 210699 130961 219485 130989
rect 219513 130961 219547 130989
rect 219575 130961 219609 130989
rect 219637 130961 219671 130989
rect 219699 130961 228485 130989
rect 228513 130961 228547 130989
rect 228575 130961 228609 130989
rect 228637 130961 228671 130989
rect 228699 130961 237485 130989
rect 237513 130961 237547 130989
rect 237575 130961 237609 130989
rect 237637 130961 237671 130989
rect 237699 130961 246485 130989
rect 246513 130961 246547 130989
rect 246575 130961 246609 130989
rect 246637 130961 246671 130989
rect 246699 130961 255485 130989
rect 255513 130961 255547 130989
rect 255575 130961 255609 130989
rect 255637 130961 255671 130989
rect 255699 130961 264485 130989
rect 264513 130961 264547 130989
rect 264575 130961 264609 130989
rect 264637 130961 264671 130989
rect 264699 130961 273485 130989
rect 273513 130961 273547 130989
rect 273575 130961 273609 130989
rect 273637 130961 273671 130989
rect 273699 130961 282485 130989
rect 282513 130961 282547 130989
rect 282575 130961 282609 130989
rect 282637 130961 282671 130989
rect 282699 130961 291485 130989
rect 291513 130961 291547 130989
rect 291575 130961 291609 130989
rect 291637 130961 291671 130989
rect 291699 130961 298728 130989
rect 298756 130961 298790 130989
rect 298818 130961 298852 130989
rect 298880 130961 298914 130989
rect 298942 130961 298990 130989
rect -958 130913 298990 130961
rect -958 128175 298990 128223
rect -958 128147 -430 128175
rect -402 128147 -368 128175
rect -340 128147 -306 128175
rect -278 128147 -244 128175
rect -216 128147 1625 128175
rect 1653 128147 1687 128175
rect 1715 128147 1749 128175
rect 1777 128147 1811 128175
rect 1839 128147 10625 128175
rect 10653 128147 10687 128175
rect 10715 128147 10749 128175
rect 10777 128147 10811 128175
rect 10839 128147 19625 128175
rect 19653 128147 19687 128175
rect 19715 128147 19749 128175
rect 19777 128147 19811 128175
rect 19839 128147 28625 128175
rect 28653 128147 28687 128175
rect 28715 128147 28749 128175
rect 28777 128147 28811 128175
rect 28839 128147 37625 128175
rect 37653 128147 37687 128175
rect 37715 128147 37749 128175
rect 37777 128147 37811 128175
rect 37839 128147 46625 128175
rect 46653 128147 46687 128175
rect 46715 128147 46749 128175
rect 46777 128147 46811 128175
rect 46839 128147 52259 128175
rect 52287 128147 52321 128175
rect 52349 128147 67619 128175
rect 67647 128147 67681 128175
rect 67709 128147 82979 128175
rect 83007 128147 83041 128175
rect 83069 128147 98339 128175
rect 98367 128147 98401 128175
rect 98429 128147 113699 128175
rect 113727 128147 113761 128175
rect 113789 128147 129059 128175
rect 129087 128147 129121 128175
rect 129149 128147 144419 128175
rect 144447 128147 144481 128175
rect 144509 128147 154625 128175
rect 154653 128147 154687 128175
rect 154715 128147 154749 128175
rect 154777 128147 154811 128175
rect 154839 128147 163625 128175
rect 163653 128147 163687 128175
rect 163715 128147 163749 128175
rect 163777 128147 163811 128175
rect 163839 128147 172625 128175
rect 172653 128147 172687 128175
rect 172715 128147 172749 128175
rect 172777 128147 172811 128175
rect 172839 128147 181625 128175
rect 181653 128147 181687 128175
rect 181715 128147 181749 128175
rect 181777 128147 181811 128175
rect 181839 128147 190625 128175
rect 190653 128147 190687 128175
rect 190715 128147 190749 128175
rect 190777 128147 190811 128175
rect 190839 128147 199625 128175
rect 199653 128147 199687 128175
rect 199715 128147 199749 128175
rect 199777 128147 199811 128175
rect 199839 128147 208625 128175
rect 208653 128147 208687 128175
rect 208715 128147 208749 128175
rect 208777 128147 208811 128175
rect 208839 128147 217625 128175
rect 217653 128147 217687 128175
rect 217715 128147 217749 128175
rect 217777 128147 217811 128175
rect 217839 128147 226625 128175
rect 226653 128147 226687 128175
rect 226715 128147 226749 128175
rect 226777 128147 226811 128175
rect 226839 128147 235625 128175
rect 235653 128147 235687 128175
rect 235715 128147 235749 128175
rect 235777 128147 235811 128175
rect 235839 128147 244625 128175
rect 244653 128147 244687 128175
rect 244715 128147 244749 128175
rect 244777 128147 244811 128175
rect 244839 128147 253625 128175
rect 253653 128147 253687 128175
rect 253715 128147 253749 128175
rect 253777 128147 253811 128175
rect 253839 128147 262625 128175
rect 262653 128147 262687 128175
rect 262715 128147 262749 128175
rect 262777 128147 262811 128175
rect 262839 128147 271625 128175
rect 271653 128147 271687 128175
rect 271715 128147 271749 128175
rect 271777 128147 271811 128175
rect 271839 128147 280625 128175
rect 280653 128147 280687 128175
rect 280715 128147 280749 128175
rect 280777 128147 280811 128175
rect 280839 128147 289625 128175
rect 289653 128147 289687 128175
rect 289715 128147 289749 128175
rect 289777 128147 289811 128175
rect 289839 128147 298248 128175
rect 298276 128147 298310 128175
rect 298338 128147 298372 128175
rect 298400 128147 298434 128175
rect 298462 128147 298990 128175
rect -958 128113 298990 128147
rect -958 128085 -430 128113
rect -402 128085 -368 128113
rect -340 128085 -306 128113
rect -278 128085 -244 128113
rect -216 128085 1625 128113
rect 1653 128085 1687 128113
rect 1715 128085 1749 128113
rect 1777 128085 1811 128113
rect 1839 128085 10625 128113
rect 10653 128085 10687 128113
rect 10715 128085 10749 128113
rect 10777 128085 10811 128113
rect 10839 128085 19625 128113
rect 19653 128085 19687 128113
rect 19715 128085 19749 128113
rect 19777 128085 19811 128113
rect 19839 128085 28625 128113
rect 28653 128085 28687 128113
rect 28715 128085 28749 128113
rect 28777 128085 28811 128113
rect 28839 128085 37625 128113
rect 37653 128085 37687 128113
rect 37715 128085 37749 128113
rect 37777 128085 37811 128113
rect 37839 128085 46625 128113
rect 46653 128085 46687 128113
rect 46715 128085 46749 128113
rect 46777 128085 46811 128113
rect 46839 128085 52259 128113
rect 52287 128085 52321 128113
rect 52349 128085 67619 128113
rect 67647 128085 67681 128113
rect 67709 128085 82979 128113
rect 83007 128085 83041 128113
rect 83069 128085 98339 128113
rect 98367 128085 98401 128113
rect 98429 128085 113699 128113
rect 113727 128085 113761 128113
rect 113789 128085 129059 128113
rect 129087 128085 129121 128113
rect 129149 128085 144419 128113
rect 144447 128085 144481 128113
rect 144509 128085 154625 128113
rect 154653 128085 154687 128113
rect 154715 128085 154749 128113
rect 154777 128085 154811 128113
rect 154839 128085 163625 128113
rect 163653 128085 163687 128113
rect 163715 128085 163749 128113
rect 163777 128085 163811 128113
rect 163839 128085 172625 128113
rect 172653 128085 172687 128113
rect 172715 128085 172749 128113
rect 172777 128085 172811 128113
rect 172839 128085 181625 128113
rect 181653 128085 181687 128113
rect 181715 128085 181749 128113
rect 181777 128085 181811 128113
rect 181839 128085 190625 128113
rect 190653 128085 190687 128113
rect 190715 128085 190749 128113
rect 190777 128085 190811 128113
rect 190839 128085 199625 128113
rect 199653 128085 199687 128113
rect 199715 128085 199749 128113
rect 199777 128085 199811 128113
rect 199839 128085 208625 128113
rect 208653 128085 208687 128113
rect 208715 128085 208749 128113
rect 208777 128085 208811 128113
rect 208839 128085 217625 128113
rect 217653 128085 217687 128113
rect 217715 128085 217749 128113
rect 217777 128085 217811 128113
rect 217839 128085 226625 128113
rect 226653 128085 226687 128113
rect 226715 128085 226749 128113
rect 226777 128085 226811 128113
rect 226839 128085 235625 128113
rect 235653 128085 235687 128113
rect 235715 128085 235749 128113
rect 235777 128085 235811 128113
rect 235839 128085 244625 128113
rect 244653 128085 244687 128113
rect 244715 128085 244749 128113
rect 244777 128085 244811 128113
rect 244839 128085 253625 128113
rect 253653 128085 253687 128113
rect 253715 128085 253749 128113
rect 253777 128085 253811 128113
rect 253839 128085 262625 128113
rect 262653 128085 262687 128113
rect 262715 128085 262749 128113
rect 262777 128085 262811 128113
rect 262839 128085 271625 128113
rect 271653 128085 271687 128113
rect 271715 128085 271749 128113
rect 271777 128085 271811 128113
rect 271839 128085 280625 128113
rect 280653 128085 280687 128113
rect 280715 128085 280749 128113
rect 280777 128085 280811 128113
rect 280839 128085 289625 128113
rect 289653 128085 289687 128113
rect 289715 128085 289749 128113
rect 289777 128085 289811 128113
rect 289839 128085 298248 128113
rect 298276 128085 298310 128113
rect 298338 128085 298372 128113
rect 298400 128085 298434 128113
rect 298462 128085 298990 128113
rect -958 128051 298990 128085
rect -958 128023 -430 128051
rect -402 128023 -368 128051
rect -340 128023 -306 128051
rect -278 128023 -244 128051
rect -216 128023 1625 128051
rect 1653 128023 1687 128051
rect 1715 128023 1749 128051
rect 1777 128023 1811 128051
rect 1839 128023 10625 128051
rect 10653 128023 10687 128051
rect 10715 128023 10749 128051
rect 10777 128023 10811 128051
rect 10839 128023 19625 128051
rect 19653 128023 19687 128051
rect 19715 128023 19749 128051
rect 19777 128023 19811 128051
rect 19839 128023 28625 128051
rect 28653 128023 28687 128051
rect 28715 128023 28749 128051
rect 28777 128023 28811 128051
rect 28839 128023 37625 128051
rect 37653 128023 37687 128051
rect 37715 128023 37749 128051
rect 37777 128023 37811 128051
rect 37839 128023 46625 128051
rect 46653 128023 46687 128051
rect 46715 128023 46749 128051
rect 46777 128023 46811 128051
rect 46839 128023 52259 128051
rect 52287 128023 52321 128051
rect 52349 128023 67619 128051
rect 67647 128023 67681 128051
rect 67709 128023 82979 128051
rect 83007 128023 83041 128051
rect 83069 128023 98339 128051
rect 98367 128023 98401 128051
rect 98429 128023 113699 128051
rect 113727 128023 113761 128051
rect 113789 128023 129059 128051
rect 129087 128023 129121 128051
rect 129149 128023 144419 128051
rect 144447 128023 144481 128051
rect 144509 128023 154625 128051
rect 154653 128023 154687 128051
rect 154715 128023 154749 128051
rect 154777 128023 154811 128051
rect 154839 128023 163625 128051
rect 163653 128023 163687 128051
rect 163715 128023 163749 128051
rect 163777 128023 163811 128051
rect 163839 128023 172625 128051
rect 172653 128023 172687 128051
rect 172715 128023 172749 128051
rect 172777 128023 172811 128051
rect 172839 128023 181625 128051
rect 181653 128023 181687 128051
rect 181715 128023 181749 128051
rect 181777 128023 181811 128051
rect 181839 128023 190625 128051
rect 190653 128023 190687 128051
rect 190715 128023 190749 128051
rect 190777 128023 190811 128051
rect 190839 128023 199625 128051
rect 199653 128023 199687 128051
rect 199715 128023 199749 128051
rect 199777 128023 199811 128051
rect 199839 128023 208625 128051
rect 208653 128023 208687 128051
rect 208715 128023 208749 128051
rect 208777 128023 208811 128051
rect 208839 128023 217625 128051
rect 217653 128023 217687 128051
rect 217715 128023 217749 128051
rect 217777 128023 217811 128051
rect 217839 128023 226625 128051
rect 226653 128023 226687 128051
rect 226715 128023 226749 128051
rect 226777 128023 226811 128051
rect 226839 128023 235625 128051
rect 235653 128023 235687 128051
rect 235715 128023 235749 128051
rect 235777 128023 235811 128051
rect 235839 128023 244625 128051
rect 244653 128023 244687 128051
rect 244715 128023 244749 128051
rect 244777 128023 244811 128051
rect 244839 128023 253625 128051
rect 253653 128023 253687 128051
rect 253715 128023 253749 128051
rect 253777 128023 253811 128051
rect 253839 128023 262625 128051
rect 262653 128023 262687 128051
rect 262715 128023 262749 128051
rect 262777 128023 262811 128051
rect 262839 128023 271625 128051
rect 271653 128023 271687 128051
rect 271715 128023 271749 128051
rect 271777 128023 271811 128051
rect 271839 128023 280625 128051
rect 280653 128023 280687 128051
rect 280715 128023 280749 128051
rect 280777 128023 280811 128051
rect 280839 128023 289625 128051
rect 289653 128023 289687 128051
rect 289715 128023 289749 128051
rect 289777 128023 289811 128051
rect 289839 128023 298248 128051
rect 298276 128023 298310 128051
rect 298338 128023 298372 128051
rect 298400 128023 298434 128051
rect 298462 128023 298990 128051
rect -958 127989 298990 128023
rect -958 127961 -430 127989
rect -402 127961 -368 127989
rect -340 127961 -306 127989
rect -278 127961 -244 127989
rect -216 127961 1625 127989
rect 1653 127961 1687 127989
rect 1715 127961 1749 127989
rect 1777 127961 1811 127989
rect 1839 127961 10625 127989
rect 10653 127961 10687 127989
rect 10715 127961 10749 127989
rect 10777 127961 10811 127989
rect 10839 127961 19625 127989
rect 19653 127961 19687 127989
rect 19715 127961 19749 127989
rect 19777 127961 19811 127989
rect 19839 127961 28625 127989
rect 28653 127961 28687 127989
rect 28715 127961 28749 127989
rect 28777 127961 28811 127989
rect 28839 127961 37625 127989
rect 37653 127961 37687 127989
rect 37715 127961 37749 127989
rect 37777 127961 37811 127989
rect 37839 127961 46625 127989
rect 46653 127961 46687 127989
rect 46715 127961 46749 127989
rect 46777 127961 46811 127989
rect 46839 127961 52259 127989
rect 52287 127961 52321 127989
rect 52349 127961 67619 127989
rect 67647 127961 67681 127989
rect 67709 127961 82979 127989
rect 83007 127961 83041 127989
rect 83069 127961 98339 127989
rect 98367 127961 98401 127989
rect 98429 127961 113699 127989
rect 113727 127961 113761 127989
rect 113789 127961 129059 127989
rect 129087 127961 129121 127989
rect 129149 127961 144419 127989
rect 144447 127961 144481 127989
rect 144509 127961 154625 127989
rect 154653 127961 154687 127989
rect 154715 127961 154749 127989
rect 154777 127961 154811 127989
rect 154839 127961 163625 127989
rect 163653 127961 163687 127989
rect 163715 127961 163749 127989
rect 163777 127961 163811 127989
rect 163839 127961 172625 127989
rect 172653 127961 172687 127989
rect 172715 127961 172749 127989
rect 172777 127961 172811 127989
rect 172839 127961 181625 127989
rect 181653 127961 181687 127989
rect 181715 127961 181749 127989
rect 181777 127961 181811 127989
rect 181839 127961 190625 127989
rect 190653 127961 190687 127989
rect 190715 127961 190749 127989
rect 190777 127961 190811 127989
rect 190839 127961 199625 127989
rect 199653 127961 199687 127989
rect 199715 127961 199749 127989
rect 199777 127961 199811 127989
rect 199839 127961 208625 127989
rect 208653 127961 208687 127989
rect 208715 127961 208749 127989
rect 208777 127961 208811 127989
rect 208839 127961 217625 127989
rect 217653 127961 217687 127989
rect 217715 127961 217749 127989
rect 217777 127961 217811 127989
rect 217839 127961 226625 127989
rect 226653 127961 226687 127989
rect 226715 127961 226749 127989
rect 226777 127961 226811 127989
rect 226839 127961 235625 127989
rect 235653 127961 235687 127989
rect 235715 127961 235749 127989
rect 235777 127961 235811 127989
rect 235839 127961 244625 127989
rect 244653 127961 244687 127989
rect 244715 127961 244749 127989
rect 244777 127961 244811 127989
rect 244839 127961 253625 127989
rect 253653 127961 253687 127989
rect 253715 127961 253749 127989
rect 253777 127961 253811 127989
rect 253839 127961 262625 127989
rect 262653 127961 262687 127989
rect 262715 127961 262749 127989
rect 262777 127961 262811 127989
rect 262839 127961 271625 127989
rect 271653 127961 271687 127989
rect 271715 127961 271749 127989
rect 271777 127961 271811 127989
rect 271839 127961 280625 127989
rect 280653 127961 280687 127989
rect 280715 127961 280749 127989
rect 280777 127961 280811 127989
rect 280839 127961 289625 127989
rect 289653 127961 289687 127989
rect 289715 127961 289749 127989
rect 289777 127961 289811 127989
rect 289839 127961 298248 127989
rect 298276 127961 298310 127989
rect 298338 127961 298372 127989
rect 298400 127961 298434 127989
rect 298462 127961 298990 127989
rect -958 127913 298990 127961
rect -958 122175 298990 122223
rect -958 122147 -910 122175
rect -882 122147 -848 122175
rect -820 122147 -786 122175
rect -758 122147 -724 122175
rect -696 122147 3485 122175
rect 3513 122147 3547 122175
rect 3575 122147 3609 122175
rect 3637 122147 3671 122175
rect 3699 122147 12485 122175
rect 12513 122147 12547 122175
rect 12575 122147 12609 122175
rect 12637 122147 12671 122175
rect 12699 122147 21485 122175
rect 21513 122147 21547 122175
rect 21575 122147 21609 122175
rect 21637 122147 21671 122175
rect 21699 122147 30485 122175
rect 30513 122147 30547 122175
rect 30575 122147 30609 122175
rect 30637 122147 30671 122175
rect 30699 122147 39485 122175
rect 39513 122147 39547 122175
rect 39575 122147 39609 122175
rect 39637 122147 39671 122175
rect 39699 122147 48485 122175
rect 48513 122147 48547 122175
rect 48575 122147 48609 122175
rect 48637 122147 48671 122175
rect 48699 122147 57485 122175
rect 57513 122147 57547 122175
rect 57575 122147 57609 122175
rect 57637 122147 57671 122175
rect 57699 122147 66485 122175
rect 66513 122147 66547 122175
rect 66575 122147 66609 122175
rect 66637 122147 66671 122175
rect 66699 122147 75485 122175
rect 75513 122147 75547 122175
rect 75575 122147 75609 122175
rect 75637 122147 75671 122175
rect 75699 122147 84485 122175
rect 84513 122147 84547 122175
rect 84575 122147 84609 122175
rect 84637 122147 84671 122175
rect 84699 122147 93485 122175
rect 93513 122147 93547 122175
rect 93575 122147 93609 122175
rect 93637 122147 93671 122175
rect 93699 122147 102485 122175
rect 102513 122147 102547 122175
rect 102575 122147 102609 122175
rect 102637 122147 102671 122175
rect 102699 122147 111485 122175
rect 111513 122147 111547 122175
rect 111575 122147 111609 122175
rect 111637 122147 111671 122175
rect 111699 122147 120485 122175
rect 120513 122147 120547 122175
rect 120575 122147 120609 122175
rect 120637 122147 120671 122175
rect 120699 122147 129485 122175
rect 129513 122147 129547 122175
rect 129575 122147 129609 122175
rect 129637 122147 129671 122175
rect 129699 122147 138485 122175
rect 138513 122147 138547 122175
rect 138575 122147 138609 122175
rect 138637 122147 138671 122175
rect 138699 122147 147485 122175
rect 147513 122147 147547 122175
rect 147575 122147 147609 122175
rect 147637 122147 147671 122175
rect 147699 122147 156485 122175
rect 156513 122147 156547 122175
rect 156575 122147 156609 122175
rect 156637 122147 156671 122175
rect 156699 122147 165485 122175
rect 165513 122147 165547 122175
rect 165575 122147 165609 122175
rect 165637 122147 165671 122175
rect 165699 122147 174485 122175
rect 174513 122147 174547 122175
rect 174575 122147 174609 122175
rect 174637 122147 174671 122175
rect 174699 122147 183485 122175
rect 183513 122147 183547 122175
rect 183575 122147 183609 122175
rect 183637 122147 183671 122175
rect 183699 122147 192485 122175
rect 192513 122147 192547 122175
rect 192575 122147 192609 122175
rect 192637 122147 192671 122175
rect 192699 122147 201485 122175
rect 201513 122147 201547 122175
rect 201575 122147 201609 122175
rect 201637 122147 201671 122175
rect 201699 122147 210485 122175
rect 210513 122147 210547 122175
rect 210575 122147 210609 122175
rect 210637 122147 210671 122175
rect 210699 122147 219485 122175
rect 219513 122147 219547 122175
rect 219575 122147 219609 122175
rect 219637 122147 219671 122175
rect 219699 122147 228485 122175
rect 228513 122147 228547 122175
rect 228575 122147 228609 122175
rect 228637 122147 228671 122175
rect 228699 122147 237485 122175
rect 237513 122147 237547 122175
rect 237575 122147 237609 122175
rect 237637 122147 237671 122175
rect 237699 122147 246485 122175
rect 246513 122147 246547 122175
rect 246575 122147 246609 122175
rect 246637 122147 246671 122175
rect 246699 122147 255485 122175
rect 255513 122147 255547 122175
rect 255575 122147 255609 122175
rect 255637 122147 255671 122175
rect 255699 122147 264485 122175
rect 264513 122147 264547 122175
rect 264575 122147 264609 122175
rect 264637 122147 264671 122175
rect 264699 122147 273485 122175
rect 273513 122147 273547 122175
rect 273575 122147 273609 122175
rect 273637 122147 273671 122175
rect 273699 122147 282485 122175
rect 282513 122147 282547 122175
rect 282575 122147 282609 122175
rect 282637 122147 282671 122175
rect 282699 122147 291485 122175
rect 291513 122147 291547 122175
rect 291575 122147 291609 122175
rect 291637 122147 291671 122175
rect 291699 122147 298728 122175
rect 298756 122147 298790 122175
rect 298818 122147 298852 122175
rect 298880 122147 298914 122175
rect 298942 122147 298990 122175
rect -958 122113 298990 122147
rect -958 122085 -910 122113
rect -882 122085 -848 122113
rect -820 122085 -786 122113
rect -758 122085 -724 122113
rect -696 122085 3485 122113
rect 3513 122085 3547 122113
rect 3575 122085 3609 122113
rect 3637 122085 3671 122113
rect 3699 122085 12485 122113
rect 12513 122085 12547 122113
rect 12575 122085 12609 122113
rect 12637 122085 12671 122113
rect 12699 122085 21485 122113
rect 21513 122085 21547 122113
rect 21575 122085 21609 122113
rect 21637 122085 21671 122113
rect 21699 122085 30485 122113
rect 30513 122085 30547 122113
rect 30575 122085 30609 122113
rect 30637 122085 30671 122113
rect 30699 122085 39485 122113
rect 39513 122085 39547 122113
rect 39575 122085 39609 122113
rect 39637 122085 39671 122113
rect 39699 122085 48485 122113
rect 48513 122085 48547 122113
rect 48575 122085 48609 122113
rect 48637 122085 48671 122113
rect 48699 122085 57485 122113
rect 57513 122085 57547 122113
rect 57575 122085 57609 122113
rect 57637 122085 57671 122113
rect 57699 122085 66485 122113
rect 66513 122085 66547 122113
rect 66575 122085 66609 122113
rect 66637 122085 66671 122113
rect 66699 122085 75485 122113
rect 75513 122085 75547 122113
rect 75575 122085 75609 122113
rect 75637 122085 75671 122113
rect 75699 122085 84485 122113
rect 84513 122085 84547 122113
rect 84575 122085 84609 122113
rect 84637 122085 84671 122113
rect 84699 122085 93485 122113
rect 93513 122085 93547 122113
rect 93575 122085 93609 122113
rect 93637 122085 93671 122113
rect 93699 122085 102485 122113
rect 102513 122085 102547 122113
rect 102575 122085 102609 122113
rect 102637 122085 102671 122113
rect 102699 122085 111485 122113
rect 111513 122085 111547 122113
rect 111575 122085 111609 122113
rect 111637 122085 111671 122113
rect 111699 122085 120485 122113
rect 120513 122085 120547 122113
rect 120575 122085 120609 122113
rect 120637 122085 120671 122113
rect 120699 122085 129485 122113
rect 129513 122085 129547 122113
rect 129575 122085 129609 122113
rect 129637 122085 129671 122113
rect 129699 122085 138485 122113
rect 138513 122085 138547 122113
rect 138575 122085 138609 122113
rect 138637 122085 138671 122113
rect 138699 122085 147485 122113
rect 147513 122085 147547 122113
rect 147575 122085 147609 122113
rect 147637 122085 147671 122113
rect 147699 122085 156485 122113
rect 156513 122085 156547 122113
rect 156575 122085 156609 122113
rect 156637 122085 156671 122113
rect 156699 122085 165485 122113
rect 165513 122085 165547 122113
rect 165575 122085 165609 122113
rect 165637 122085 165671 122113
rect 165699 122085 174485 122113
rect 174513 122085 174547 122113
rect 174575 122085 174609 122113
rect 174637 122085 174671 122113
rect 174699 122085 183485 122113
rect 183513 122085 183547 122113
rect 183575 122085 183609 122113
rect 183637 122085 183671 122113
rect 183699 122085 192485 122113
rect 192513 122085 192547 122113
rect 192575 122085 192609 122113
rect 192637 122085 192671 122113
rect 192699 122085 201485 122113
rect 201513 122085 201547 122113
rect 201575 122085 201609 122113
rect 201637 122085 201671 122113
rect 201699 122085 210485 122113
rect 210513 122085 210547 122113
rect 210575 122085 210609 122113
rect 210637 122085 210671 122113
rect 210699 122085 219485 122113
rect 219513 122085 219547 122113
rect 219575 122085 219609 122113
rect 219637 122085 219671 122113
rect 219699 122085 228485 122113
rect 228513 122085 228547 122113
rect 228575 122085 228609 122113
rect 228637 122085 228671 122113
rect 228699 122085 237485 122113
rect 237513 122085 237547 122113
rect 237575 122085 237609 122113
rect 237637 122085 237671 122113
rect 237699 122085 246485 122113
rect 246513 122085 246547 122113
rect 246575 122085 246609 122113
rect 246637 122085 246671 122113
rect 246699 122085 255485 122113
rect 255513 122085 255547 122113
rect 255575 122085 255609 122113
rect 255637 122085 255671 122113
rect 255699 122085 264485 122113
rect 264513 122085 264547 122113
rect 264575 122085 264609 122113
rect 264637 122085 264671 122113
rect 264699 122085 273485 122113
rect 273513 122085 273547 122113
rect 273575 122085 273609 122113
rect 273637 122085 273671 122113
rect 273699 122085 282485 122113
rect 282513 122085 282547 122113
rect 282575 122085 282609 122113
rect 282637 122085 282671 122113
rect 282699 122085 291485 122113
rect 291513 122085 291547 122113
rect 291575 122085 291609 122113
rect 291637 122085 291671 122113
rect 291699 122085 298728 122113
rect 298756 122085 298790 122113
rect 298818 122085 298852 122113
rect 298880 122085 298914 122113
rect 298942 122085 298990 122113
rect -958 122051 298990 122085
rect -958 122023 -910 122051
rect -882 122023 -848 122051
rect -820 122023 -786 122051
rect -758 122023 -724 122051
rect -696 122023 3485 122051
rect 3513 122023 3547 122051
rect 3575 122023 3609 122051
rect 3637 122023 3671 122051
rect 3699 122023 12485 122051
rect 12513 122023 12547 122051
rect 12575 122023 12609 122051
rect 12637 122023 12671 122051
rect 12699 122023 21485 122051
rect 21513 122023 21547 122051
rect 21575 122023 21609 122051
rect 21637 122023 21671 122051
rect 21699 122023 30485 122051
rect 30513 122023 30547 122051
rect 30575 122023 30609 122051
rect 30637 122023 30671 122051
rect 30699 122023 39485 122051
rect 39513 122023 39547 122051
rect 39575 122023 39609 122051
rect 39637 122023 39671 122051
rect 39699 122023 48485 122051
rect 48513 122023 48547 122051
rect 48575 122023 48609 122051
rect 48637 122023 48671 122051
rect 48699 122023 57485 122051
rect 57513 122023 57547 122051
rect 57575 122023 57609 122051
rect 57637 122023 57671 122051
rect 57699 122023 66485 122051
rect 66513 122023 66547 122051
rect 66575 122023 66609 122051
rect 66637 122023 66671 122051
rect 66699 122023 75485 122051
rect 75513 122023 75547 122051
rect 75575 122023 75609 122051
rect 75637 122023 75671 122051
rect 75699 122023 84485 122051
rect 84513 122023 84547 122051
rect 84575 122023 84609 122051
rect 84637 122023 84671 122051
rect 84699 122023 93485 122051
rect 93513 122023 93547 122051
rect 93575 122023 93609 122051
rect 93637 122023 93671 122051
rect 93699 122023 102485 122051
rect 102513 122023 102547 122051
rect 102575 122023 102609 122051
rect 102637 122023 102671 122051
rect 102699 122023 111485 122051
rect 111513 122023 111547 122051
rect 111575 122023 111609 122051
rect 111637 122023 111671 122051
rect 111699 122023 120485 122051
rect 120513 122023 120547 122051
rect 120575 122023 120609 122051
rect 120637 122023 120671 122051
rect 120699 122023 129485 122051
rect 129513 122023 129547 122051
rect 129575 122023 129609 122051
rect 129637 122023 129671 122051
rect 129699 122023 138485 122051
rect 138513 122023 138547 122051
rect 138575 122023 138609 122051
rect 138637 122023 138671 122051
rect 138699 122023 147485 122051
rect 147513 122023 147547 122051
rect 147575 122023 147609 122051
rect 147637 122023 147671 122051
rect 147699 122023 156485 122051
rect 156513 122023 156547 122051
rect 156575 122023 156609 122051
rect 156637 122023 156671 122051
rect 156699 122023 165485 122051
rect 165513 122023 165547 122051
rect 165575 122023 165609 122051
rect 165637 122023 165671 122051
rect 165699 122023 174485 122051
rect 174513 122023 174547 122051
rect 174575 122023 174609 122051
rect 174637 122023 174671 122051
rect 174699 122023 183485 122051
rect 183513 122023 183547 122051
rect 183575 122023 183609 122051
rect 183637 122023 183671 122051
rect 183699 122023 192485 122051
rect 192513 122023 192547 122051
rect 192575 122023 192609 122051
rect 192637 122023 192671 122051
rect 192699 122023 201485 122051
rect 201513 122023 201547 122051
rect 201575 122023 201609 122051
rect 201637 122023 201671 122051
rect 201699 122023 210485 122051
rect 210513 122023 210547 122051
rect 210575 122023 210609 122051
rect 210637 122023 210671 122051
rect 210699 122023 219485 122051
rect 219513 122023 219547 122051
rect 219575 122023 219609 122051
rect 219637 122023 219671 122051
rect 219699 122023 228485 122051
rect 228513 122023 228547 122051
rect 228575 122023 228609 122051
rect 228637 122023 228671 122051
rect 228699 122023 237485 122051
rect 237513 122023 237547 122051
rect 237575 122023 237609 122051
rect 237637 122023 237671 122051
rect 237699 122023 246485 122051
rect 246513 122023 246547 122051
rect 246575 122023 246609 122051
rect 246637 122023 246671 122051
rect 246699 122023 255485 122051
rect 255513 122023 255547 122051
rect 255575 122023 255609 122051
rect 255637 122023 255671 122051
rect 255699 122023 264485 122051
rect 264513 122023 264547 122051
rect 264575 122023 264609 122051
rect 264637 122023 264671 122051
rect 264699 122023 273485 122051
rect 273513 122023 273547 122051
rect 273575 122023 273609 122051
rect 273637 122023 273671 122051
rect 273699 122023 282485 122051
rect 282513 122023 282547 122051
rect 282575 122023 282609 122051
rect 282637 122023 282671 122051
rect 282699 122023 291485 122051
rect 291513 122023 291547 122051
rect 291575 122023 291609 122051
rect 291637 122023 291671 122051
rect 291699 122023 298728 122051
rect 298756 122023 298790 122051
rect 298818 122023 298852 122051
rect 298880 122023 298914 122051
rect 298942 122023 298990 122051
rect -958 121989 298990 122023
rect -958 121961 -910 121989
rect -882 121961 -848 121989
rect -820 121961 -786 121989
rect -758 121961 -724 121989
rect -696 121961 3485 121989
rect 3513 121961 3547 121989
rect 3575 121961 3609 121989
rect 3637 121961 3671 121989
rect 3699 121961 12485 121989
rect 12513 121961 12547 121989
rect 12575 121961 12609 121989
rect 12637 121961 12671 121989
rect 12699 121961 21485 121989
rect 21513 121961 21547 121989
rect 21575 121961 21609 121989
rect 21637 121961 21671 121989
rect 21699 121961 30485 121989
rect 30513 121961 30547 121989
rect 30575 121961 30609 121989
rect 30637 121961 30671 121989
rect 30699 121961 39485 121989
rect 39513 121961 39547 121989
rect 39575 121961 39609 121989
rect 39637 121961 39671 121989
rect 39699 121961 48485 121989
rect 48513 121961 48547 121989
rect 48575 121961 48609 121989
rect 48637 121961 48671 121989
rect 48699 121961 57485 121989
rect 57513 121961 57547 121989
rect 57575 121961 57609 121989
rect 57637 121961 57671 121989
rect 57699 121961 66485 121989
rect 66513 121961 66547 121989
rect 66575 121961 66609 121989
rect 66637 121961 66671 121989
rect 66699 121961 75485 121989
rect 75513 121961 75547 121989
rect 75575 121961 75609 121989
rect 75637 121961 75671 121989
rect 75699 121961 84485 121989
rect 84513 121961 84547 121989
rect 84575 121961 84609 121989
rect 84637 121961 84671 121989
rect 84699 121961 93485 121989
rect 93513 121961 93547 121989
rect 93575 121961 93609 121989
rect 93637 121961 93671 121989
rect 93699 121961 102485 121989
rect 102513 121961 102547 121989
rect 102575 121961 102609 121989
rect 102637 121961 102671 121989
rect 102699 121961 111485 121989
rect 111513 121961 111547 121989
rect 111575 121961 111609 121989
rect 111637 121961 111671 121989
rect 111699 121961 120485 121989
rect 120513 121961 120547 121989
rect 120575 121961 120609 121989
rect 120637 121961 120671 121989
rect 120699 121961 129485 121989
rect 129513 121961 129547 121989
rect 129575 121961 129609 121989
rect 129637 121961 129671 121989
rect 129699 121961 138485 121989
rect 138513 121961 138547 121989
rect 138575 121961 138609 121989
rect 138637 121961 138671 121989
rect 138699 121961 147485 121989
rect 147513 121961 147547 121989
rect 147575 121961 147609 121989
rect 147637 121961 147671 121989
rect 147699 121961 156485 121989
rect 156513 121961 156547 121989
rect 156575 121961 156609 121989
rect 156637 121961 156671 121989
rect 156699 121961 165485 121989
rect 165513 121961 165547 121989
rect 165575 121961 165609 121989
rect 165637 121961 165671 121989
rect 165699 121961 174485 121989
rect 174513 121961 174547 121989
rect 174575 121961 174609 121989
rect 174637 121961 174671 121989
rect 174699 121961 183485 121989
rect 183513 121961 183547 121989
rect 183575 121961 183609 121989
rect 183637 121961 183671 121989
rect 183699 121961 192485 121989
rect 192513 121961 192547 121989
rect 192575 121961 192609 121989
rect 192637 121961 192671 121989
rect 192699 121961 201485 121989
rect 201513 121961 201547 121989
rect 201575 121961 201609 121989
rect 201637 121961 201671 121989
rect 201699 121961 210485 121989
rect 210513 121961 210547 121989
rect 210575 121961 210609 121989
rect 210637 121961 210671 121989
rect 210699 121961 219485 121989
rect 219513 121961 219547 121989
rect 219575 121961 219609 121989
rect 219637 121961 219671 121989
rect 219699 121961 228485 121989
rect 228513 121961 228547 121989
rect 228575 121961 228609 121989
rect 228637 121961 228671 121989
rect 228699 121961 237485 121989
rect 237513 121961 237547 121989
rect 237575 121961 237609 121989
rect 237637 121961 237671 121989
rect 237699 121961 246485 121989
rect 246513 121961 246547 121989
rect 246575 121961 246609 121989
rect 246637 121961 246671 121989
rect 246699 121961 255485 121989
rect 255513 121961 255547 121989
rect 255575 121961 255609 121989
rect 255637 121961 255671 121989
rect 255699 121961 264485 121989
rect 264513 121961 264547 121989
rect 264575 121961 264609 121989
rect 264637 121961 264671 121989
rect 264699 121961 273485 121989
rect 273513 121961 273547 121989
rect 273575 121961 273609 121989
rect 273637 121961 273671 121989
rect 273699 121961 282485 121989
rect 282513 121961 282547 121989
rect 282575 121961 282609 121989
rect 282637 121961 282671 121989
rect 282699 121961 291485 121989
rect 291513 121961 291547 121989
rect 291575 121961 291609 121989
rect 291637 121961 291671 121989
rect 291699 121961 298728 121989
rect 298756 121961 298790 121989
rect 298818 121961 298852 121989
rect 298880 121961 298914 121989
rect 298942 121961 298990 121989
rect -958 121913 298990 121961
rect -958 119175 298990 119223
rect -958 119147 -430 119175
rect -402 119147 -368 119175
rect -340 119147 -306 119175
rect -278 119147 -244 119175
rect -216 119147 1625 119175
rect 1653 119147 1687 119175
rect 1715 119147 1749 119175
rect 1777 119147 1811 119175
rect 1839 119147 10625 119175
rect 10653 119147 10687 119175
rect 10715 119147 10749 119175
rect 10777 119147 10811 119175
rect 10839 119147 19625 119175
rect 19653 119147 19687 119175
rect 19715 119147 19749 119175
rect 19777 119147 19811 119175
rect 19839 119147 28625 119175
rect 28653 119147 28687 119175
rect 28715 119147 28749 119175
rect 28777 119147 28811 119175
rect 28839 119147 37625 119175
rect 37653 119147 37687 119175
rect 37715 119147 37749 119175
rect 37777 119147 37811 119175
rect 37839 119147 46625 119175
rect 46653 119147 46687 119175
rect 46715 119147 46749 119175
rect 46777 119147 46811 119175
rect 46839 119147 55625 119175
rect 55653 119147 55687 119175
rect 55715 119147 55749 119175
rect 55777 119147 55811 119175
rect 55839 119147 64625 119175
rect 64653 119147 64687 119175
rect 64715 119147 64749 119175
rect 64777 119147 64811 119175
rect 64839 119147 73625 119175
rect 73653 119147 73687 119175
rect 73715 119147 73749 119175
rect 73777 119147 73811 119175
rect 73839 119147 82625 119175
rect 82653 119147 82687 119175
rect 82715 119147 82749 119175
rect 82777 119147 82811 119175
rect 82839 119147 91625 119175
rect 91653 119147 91687 119175
rect 91715 119147 91749 119175
rect 91777 119147 91811 119175
rect 91839 119147 100625 119175
rect 100653 119147 100687 119175
rect 100715 119147 100749 119175
rect 100777 119147 100811 119175
rect 100839 119147 109625 119175
rect 109653 119147 109687 119175
rect 109715 119147 109749 119175
rect 109777 119147 109811 119175
rect 109839 119147 118625 119175
rect 118653 119147 118687 119175
rect 118715 119147 118749 119175
rect 118777 119147 118811 119175
rect 118839 119147 127625 119175
rect 127653 119147 127687 119175
rect 127715 119147 127749 119175
rect 127777 119147 127811 119175
rect 127839 119147 136625 119175
rect 136653 119147 136687 119175
rect 136715 119147 136749 119175
rect 136777 119147 136811 119175
rect 136839 119147 145625 119175
rect 145653 119147 145687 119175
rect 145715 119147 145749 119175
rect 145777 119147 145811 119175
rect 145839 119147 154625 119175
rect 154653 119147 154687 119175
rect 154715 119147 154749 119175
rect 154777 119147 154811 119175
rect 154839 119147 163625 119175
rect 163653 119147 163687 119175
rect 163715 119147 163749 119175
rect 163777 119147 163811 119175
rect 163839 119147 172625 119175
rect 172653 119147 172687 119175
rect 172715 119147 172749 119175
rect 172777 119147 172811 119175
rect 172839 119147 181625 119175
rect 181653 119147 181687 119175
rect 181715 119147 181749 119175
rect 181777 119147 181811 119175
rect 181839 119147 190625 119175
rect 190653 119147 190687 119175
rect 190715 119147 190749 119175
rect 190777 119147 190811 119175
rect 190839 119147 199625 119175
rect 199653 119147 199687 119175
rect 199715 119147 199749 119175
rect 199777 119147 199811 119175
rect 199839 119147 208625 119175
rect 208653 119147 208687 119175
rect 208715 119147 208749 119175
rect 208777 119147 208811 119175
rect 208839 119147 217625 119175
rect 217653 119147 217687 119175
rect 217715 119147 217749 119175
rect 217777 119147 217811 119175
rect 217839 119147 226625 119175
rect 226653 119147 226687 119175
rect 226715 119147 226749 119175
rect 226777 119147 226811 119175
rect 226839 119147 235625 119175
rect 235653 119147 235687 119175
rect 235715 119147 235749 119175
rect 235777 119147 235811 119175
rect 235839 119147 244625 119175
rect 244653 119147 244687 119175
rect 244715 119147 244749 119175
rect 244777 119147 244811 119175
rect 244839 119147 253625 119175
rect 253653 119147 253687 119175
rect 253715 119147 253749 119175
rect 253777 119147 253811 119175
rect 253839 119147 262625 119175
rect 262653 119147 262687 119175
rect 262715 119147 262749 119175
rect 262777 119147 262811 119175
rect 262839 119147 271625 119175
rect 271653 119147 271687 119175
rect 271715 119147 271749 119175
rect 271777 119147 271811 119175
rect 271839 119147 280625 119175
rect 280653 119147 280687 119175
rect 280715 119147 280749 119175
rect 280777 119147 280811 119175
rect 280839 119147 289625 119175
rect 289653 119147 289687 119175
rect 289715 119147 289749 119175
rect 289777 119147 289811 119175
rect 289839 119147 298248 119175
rect 298276 119147 298310 119175
rect 298338 119147 298372 119175
rect 298400 119147 298434 119175
rect 298462 119147 298990 119175
rect -958 119113 298990 119147
rect -958 119085 -430 119113
rect -402 119085 -368 119113
rect -340 119085 -306 119113
rect -278 119085 -244 119113
rect -216 119085 1625 119113
rect 1653 119085 1687 119113
rect 1715 119085 1749 119113
rect 1777 119085 1811 119113
rect 1839 119085 10625 119113
rect 10653 119085 10687 119113
rect 10715 119085 10749 119113
rect 10777 119085 10811 119113
rect 10839 119085 19625 119113
rect 19653 119085 19687 119113
rect 19715 119085 19749 119113
rect 19777 119085 19811 119113
rect 19839 119085 28625 119113
rect 28653 119085 28687 119113
rect 28715 119085 28749 119113
rect 28777 119085 28811 119113
rect 28839 119085 37625 119113
rect 37653 119085 37687 119113
rect 37715 119085 37749 119113
rect 37777 119085 37811 119113
rect 37839 119085 46625 119113
rect 46653 119085 46687 119113
rect 46715 119085 46749 119113
rect 46777 119085 46811 119113
rect 46839 119085 55625 119113
rect 55653 119085 55687 119113
rect 55715 119085 55749 119113
rect 55777 119085 55811 119113
rect 55839 119085 64625 119113
rect 64653 119085 64687 119113
rect 64715 119085 64749 119113
rect 64777 119085 64811 119113
rect 64839 119085 73625 119113
rect 73653 119085 73687 119113
rect 73715 119085 73749 119113
rect 73777 119085 73811 119113
rect 73839 119085 82625 119113
rect 82653 119085 82687 119113
rect 82715 119085 82749 119113
rect 82777 119085 82811 119113
rect 82839 119085 91625 119113
rect 91653 119085 91687 119113
rect 91715 119085 91749 119113
rect 91777 119085 91811 119113
rect 91839 119085 100625 119113
rect 100653 119085 100687 119113
rect 100715 119085 100749 119113
rect 100777 119085 100811 119113
rect 100839 119085 109625 119113
rect 109653 119085 109687 119113
rect 109715 119085 109749 119113
rect 109777 119085 109811 119113
rect 109839 119085 118625 119113
rect 118653 119085 118687 119113
rect 118715 119085 118749 119113
rect 118777 119085 118811 119113
rect 118839 119085 127625 119113
rect 127653 119085 127687 119113
rect 127715 119085 127749 119113
rect 127777 119085 127811 119113
rect 127839 119085 136625 119113
rect 136653 119085 136687 119113
rect 136715 119085 136749 119113
rect 136777 119085 136811 119113
rect 136839 119085 145625 119113
rect 145653 119085 145687 119113
rect 145715 119085 145749 119113
rect 145777 119085 145811 119113
rect 145839 119085 154625 119113
rect 154653 119085 154687 119113
rect 154715 119085 154749 119113
rect 154777 119085 154811 119113
rect 154839 119085 163625 119113
rect 163653 119085 163687 119113
rect 163715 119085 163749 119113
rect 163777 119085 163811 119113
rect 163839 119085 172625 119113
rect 172653 119085 172687 119113
rect 172715 119085 172749 119113
rect 172777 119085 172811 119113
rect 172839 119085 181625 119113
rect 181653 119085 181687 119113
rect 181715 119085 181749 119113
rect 181777 119085 181811 119113
rect 181839 119085 190625 119113
rect 190653 119085 190687 119113
rect 190715 119085 190749 119113
rect 190777 119085 190811 119113
rect 190839 119085 199625 119113
rect 199653 119085 199687 119113
rect 199715 119085 199749 119113
rect 199777 119085 199811 119113
rect 199839 119085 208625 119113
rect 208653 119085 208687 119113
rect 208715 119085 208749 119113
rect 208777 119085 208811 119113
rect 208839 119085 217625 119113
rect 217653 119085 217687 119113
rect 217715 119085 217749 119113
rect 217777 119085 217811 119113
rect 217839 119085 226625 119113
rect 226653 119085 226687 119113
rect 226715 119085 226749 119113
rect 226777 119085 226811 119113
rect 226839 119085 235625 119113
rect 235653 119085 235687 119113
rect 235715 119085 235749 119113
rect 235777 119085 235811 119113
rect 235839 119085 244625 119113
rect 244653 119085 244687 119113
rect 244715 119085 244749 119113
rect 244777 119085 244811 119113
rect 244839 119085 253625 119113
rect 253653 119085 253687 119113
rect 253715 119085 253749 119113
rect 253777 119085 253811 119113
rect 253839 119085 262625 119113
rect 262653 119085 262687 119113
rect 262715 119085 262749 119113
rect 262777 119085 262811 119113
rect 262839 119085 271625 119113
rect 271653 119085 271687 119113
rect 271715 119085 271749 119113
rect 271777 119085 271811 119113
rect 271839 119085 280625 119113
rect 280653 119085 280687 119113
rect 280715 119085 280749 119113
rect 280777 119085 280811 119113
rect 280839 119085 289625 119113
rect 289653 119085 289687 119113
rect 289715 119085 289749 119113
rect 289777 119085 289811 119113
rect 289839 119085 298248 119113
rect 298276 119085 298310 119113
rect 298338 119085 298372 119113
rect 298400 119085 298434 119113
rect 298462 119085 298990 119113
rect -958 119051 298990 119085
rect -958 119023 -430 119051
rect -402 119023 -368 119051
rect -340 119023 -306 119051
rect -278 119023 -244 119051
rect -216 119023 1625 119051
rect 1653 119023 1687 119051
rect 1715 119023 1749 119051
rect 1777 119023 1811 119051
rect 1839 119023 10625 119051
rect 10653 119023 10687 119051
rect 10715 119023 10749 119051
rect 10777 119023 10811 119051
rect 10839 119023 19625 119051
rect 19653 119023 19687 119051
rect 19715 119023 19749 119051
rect 19777 119023 19811 119051
rect 19839 119023 28625 119051
rect 28653 119023 28687 119051
rect 28715 119023 28749 119051
rect 28777 119023 28811 119051
rect 28839 119023 37625 119051
rect 37653 119023 37687 119051
rect 37715 119023 37749 119051
rect 37777 119023 37811 119051
rect 37839 119023 46625 119051
rect 46653 119023 46687 119051
rect 46715 119023 46749 119051
rect 46777 119023 46811 119051
rect 46839 119023 55625 119051
rect 55653 119023 55687 119051
rect 55715 119023 55749 119051
rect 55777 119023 55811 119051
rect 55839 119023 64625 119051
rect 64653 119023 64687 119051
rect 64715 119023 64749 119051
rect 64777 119023 64811 119051
rect 64839 119023 73625 119051
rect 73653 119023 73687 119051
rect 73715 119023 73749 119051
rect 73777 119023 73811 119051
rect 73839 119023 82625 119051
rect 82653 119023 82687 119051
rect 82715 119023 82749 119051
rect 82777 119023 82811 119051
rect 82839 119023 91625 119051
rect 91653 119023 91687 119051
rect 91715 119023 91749 119051
rect 91777 119023 91811 119051
rect 91839 119023 100625 119051
rect 100653 119023 100687 119051
rect 100715 119023 100749 119051
rect 100777 119023 100811 119051
rect 100839 119023 109625 119051
rect 109653 119023 109687 119051
rect 109715 119023 109749 119051
rect 109777 119023 109811 119051
rect 109839 119023 118625 119051
rect 118653 119023 118687 119051
rect 118715 119023 118749 119051
rect 118777 119023 118811 119051
rect 118839 119023 127625 119051
rect 127653 119023 127687 119051
rect 127715 119023 127749 119051
rect 127777 119023 127811 119051
rect 127839 119023 136625 119051
rect 136653 119023 136687 119051
rect 136715 119023 136749 119051
rect 136777 119023 136811 119051
rect 136839 119023 145625 119051
rect 145653 119023 145687 119051
rect 145715 119023 145749 119051
rect 145777 119023 145811 119051
rect 145839 119023 154625 119051
rect 154653 119023 154687 119051
rect 154715 119023 154749 119051
rect 154777 119023 154811 119051
rect 154839 119023 163625 119051
rect 163653 119023 163687 119051
rect 163715 119023 163749 119051
rect 163777 119023 163811 119051
rect 163839 119023 172625 119051
rect 172653 119023 172687 119051
rect 172715 119023 172749 119051
rect 172777 119023 172811 119051
rect 172839 119023 181625 119051
rect 181653 119023 181687 119051
rect 181715 119023 181749 119051
rect 181777 119023 181811 119051
rect 181839 119023 190625 119051
rect 190653 119023 190687 119051
rect 190715 119023 190749 119051
rect 190777 119023 190811 119051
rect 190839 119023 199625 119051
rect 199653 119023 199687 119051
rect 199715 119023 199749 119051
rect 199777 119023 199811 119051
rect 199839 119023 208625 119051
rect 208653 119023 208687 119051
rect 208715 119023 208749 119051
rect 208777 119023 208811 119051
rect 208839 119023 217625 119051
rect 217653 119023 217687 119051
rect 217715 119023 217749 119051
rect 217777 119023 217811 119051
rect 217839 119023 226625 119051
rect 226653 119023 226687 119051
rect 226715 119023 226749 119051
rect 226777 119023 226811 119051
rect 226839 119023 235625 119051
rect 235653 119023 235687 119051
rect 235715 119023 235749 119051
rect 235777 119023 235811 119051
rect 235839 119023 244625 119051
rect 244653 119023 244687 119051
rect 244715 119023 244749 119051
rect 244777 119023 244811 119051
rect 244839 119023 253625 119051
rect 253653 119023 253687 119051
rect 253715 119023 253749 119051
rect 253777 119023 253811 119051
rect 253839 119023 262625 119051
rect 262653 119023 262687 119051
rect 262715 119023 262749 119051
rect 262777 119023 262811 119051
rect 262839 119023 271625 119051
rect 271653 119023 271687 119051
rect 271715 119023 271749 119051
rect 271777 119023 271811 119051
rect 271839 119023 280625 119051
rect 280653 119023 280687 119051
rect 280715 119023 280749 119051
rect 280777 119023 280811 119051
rect 280839 119023 289625 119051
rect 289653 119023 289687 119051
rect 289715 119023 289749 119051
rect 289777 119023 289811 119051
rect 289839 119023 298248 119051
rect 298276 119023 298310 119051
rect 298338 119023 298372 119051
rect 298400 119023 298434 119051
rect 298462 119023 298990 119051
rect -958 118989 298990 119023
rect -958 118961 -430 118989
rect -402 118961 -368 118989
rect -340 118961 -306 118989
rect -278 118961 -244 118989
rect -216 118961 1625 118989
rect 1653 118961 1687 118989
rect 1715 118961 1749 118989
rect 1777 118961 1811 118989
rect 1839 118961 10625 118989
rect 10653 118961 10687 118989
rect 10715 118961 10749 118989
rect 10777 118961 10811 118989
rect 10839 118961 19625 118989
rect 19653 118961 19687 118989
rect 19715 118961 19749 118989
rect 19777 118961 19811 118989
rect 19839 118961 28625 118989
rect 28653 118961 28687 118989
rect 28715 118961 28749 118989
rect 28777 118961 28811 118989
rect 28839 118961 37625 118989
rect 37653 118961 37687 118989
rect 37715 118961 37749 118989
rect 37777 118961 37811 118989
rect 37839 118961 46625 118989
rect 46653 118961 46687 118989
rect 46715 118961 46749 118989
rect 46777 118961 46811 118989
rect 46839 118961 55625 118989
rect 55653 118961 55687 118989
rect 55715 118961 55749 118989
rect 55777 118961 55811 118989
rect 55839 118961 64625 118989
rect 64653 118961 64687 118989
rect 64715 118961 64749 118989
rect 64777 118961 64811 118989
rect 64839 118961 73625 118989
rect 73653 118961 73687 118989
rect 73715 118961 73749 118989
rect 73777 118961 73811 118989
rect 73839 118961 82625 118989
rect 82653 118961 82687 118989
rect 82715 118961 82749 118989
rect 82777 118961 82811 118989
rect 82839 118961 91625 118989
rect 91653 118961 91687 118989
rect 91715 118961 91749 118989
rect 91777 118961 91811 118989
rect 91839 118961 100625 118989
rect 100653 118961 100687 118989
rect 100715 118961 100749 118989
rect 100777 118961 100811 118989
rect 100839 118961 109625 118989
rect 109653 118961 109687 118989
rect 109715 118961 109749 118989
rect 109777 118961 109811 118989
rect 109839 118961 118625 118989
rect 118653 118961 118687 118989
rect 118715 118961 118749 118989
rect 118777 118961 118811 118989
rect 118839 118961 127625 118989
rect 127653 118961 127687 118989
rect 127715 118961 127749 118989
rect 127777 118961 127811 118989
rect 127839 118961 136625 118989
rect 136653 118961 136687 118989
rect 136715 118961 136749 118989
rect 136777 118961 136811 118989
rect 136839 118961 145625 118989
rect 145653 118961 145687 118989
rect 145715 118961 145749 118989
rect 145777 118961 145811 118989
rect 145839 118961 154625 118989
rect 154653 118961 154687 118989
rect 154715 118961 154749 118989
rect 154777 118961 154811 118989
rect 154839 118961 163625 118989
rect 163653 118961 163687 118989
rect 163715 118961 163749 118989
rect 163777 118961 163811 118989
rect 163839 118961 172625 118989
rect 172653 118961 172687 118989
rect 172715 118961 172749 118989
rect 172777 118961 172811 118989
rect 172839 118961 181625 118989
rect 181653 118961 181687 118989
rect 181715 118961 181749 118989
rect 181777 118961 181811 118989
rect 181839 118961 190625 118989
rect 190653 118961 190687 118989
rect 190715 118961 190749 118989
rect 190777 118961 190811 118989
rect 190839 118961 199625 118989
rect 199653 118961 199687 118989
rect 199715 118961 199749 118989
rect 199777 118961 199811 118989
rect 199839 118961 208625 118989
rect 208653 118961 208687 118989
rect 208715 118961 208749 118989
rect 208777 118961 208811 118989
rect 208839 118961 217625 118989
rect 217653 118961 217687 118989
rect 217715 118961 217749 118989
rect 217777 118961 217811 118989
rect 217839 118961 226625 118989
rect 226653 118961 226687 118989
rect 226715 118961 226749 118989
rect 226777 118961 226811 118989
rect 226839 118961 235625 118989
rect 235653 118961 235687 118989
rect 235715 118961 235749 118989
rect 235777 118961 235811 118989
rect 235839 118961 244625 118989
rect 244653 118961 244687 118989
rect 244715 118961 244749 118989
rect 244777 118961 244811 118989
rect 244839 118961 253625 118989
rect 253653 118961 253687 118989
rect 253715 118961 253749 118989
rect 253777 118961 253811 118989
rect 253839 118961 262625 118989
rect 262653 118961 262687 118989
rect 262715 118961 262749 118989
rect 262777 118961 262811 118989
rect 262839 118961 271625 118989
rect 271653 118961 271687 118989
rect 271715 118961 271749 118989
rect 271777 118961 271811 118989
rect 271839 118961 280625 118989
rect 280653 118961 280687 118989
rect 280715 118961 280749 118989
rect 280777 118961 280811 118989
rect 280839 118961 289625 118989
rect 289653 118961 289687 118989
rect 289715 118961 289749 118989
rect 289777 118961 289811 118989
rect 289839 118961 298248 118989
rect 298276 118961 298310 118989
rect 298338 118961 298372 118989
rect 298400 118961 298434 118989
rect 298462 118961 298990 118989
rect -958 118913 298990 118961
rect -958 113175 298990 113223
rect -958 113147 -910 113175
rect -882 113147 -848 113175
rect -820 113147 -786 113175
rect -758 113147 -724 113175
rect -696 113147 3485 113175
rect 3513 113147 3547 113175
rect 3575 113147 3609 113175
rect 3637 113147 3671 113175
rect 3699 113147 12485 113175
rect 12513 113147 12547 113175
rect 12575 113147 12609 113175
rect 12637 113147 12671 113175
rect 12699 113147 21485 113175
rect 21513 113147 21547 113175
rect 21575 113147 21609 113175
rect 21637 113147 21671 113175
rect 21699 113147 30485 113175
rect 30513 113147 30547 113175
rect 30575 113147 30609 113175
rect 30637 113147 30671 113175
rect 30699 113147 39485 113175
rect 39513 113147 39547 113175
rect 39575 113147 39609 113175
rect 39637 113147 39671 113175
rect 39699 113147 48485 113175
rect 48513 113147 48547 113175
rect 48575 113147 48609 113175
rect 48637 113147 48671 113175
rect 48699 113147 57485 113175
rect 57513 113147 57547 113175
rect 57575 113147 57609 113175
rect 57637 113147 57671 113175
rect 57699 113147 66485 113175
rect 66513 113147 66547 113175
rect 66575 113147 66609 113175
rect 66637 113147 66671 113175
rect 66699 113147 75485 113175
rect 75513 113147 75547 113175
rect 75575 113147 75609 113175
rect 75637 113147 75671 113175
rect 75699 113147 84485 113175
rect 84513 113147 84547 113175
rect 84575 113147 84609 113175
rect 84637 113147 84671 113175
rect 84699 113147 93485 113175
rect 93513 113147 93547 113175
rect 93575 113147 93609 113175
rect 93637 113147 93671 113175
rect 93699 113147 102485 113175
rect 102513 113147 102547 113175
rect 102575 113147 102609 113175
rect 102637 113147 102671 113175
rect 102699 113147 111485 113175
rect 111513 113147 111547 113175
rect 111575 113147 111609 113175
rect 111637 113147 111671 113175
rect 111699 113147 120485 113175
rect 120513 113147 120547 113175
rect 120575 113147 120609 113175
rect 120637 113147 120671 113175
rect 120699 113147 129485 113175
rect 129513 113147 129547 113175
rect 129575 113147 129609 113175
rect 129637 113147 129671 113175
rect 129699 113147 138485 113175
rect 138513 113147 138547 113175
rect 138575 113147 138609 113175
rect 138637 113147 138671 113175
rect 138699 113147 147485 113175
rect 147513 113147 147547 113175
rect 147575 113147 147609 113175
rect 147637 113147 147671 113175
rect 147699 113147 156485 113175
rect 156513 113147 156547 113175
rect 156575 113147 156609 113175
rect 156637 113147 156671 113175
rect 156699 113147 165485 113175
rect 165513 113147 165547 113175
rect 165575 113147 165609 113175
rect 165637 113147 165671 113175
rect 165699 113147 174485 113175
rect 174513 113147 174547 113175
rect 174575 113147 174609 113175
rect 174637 113147 174671 113175
rect 174699 113147 183485 113175
rect 183513 113147 183547 113175
rect 183575 113147 183609 113175
rect 183637 113147 183671 113175
rect 183699 113147 192485 113175
rect 192513 113147 192547 113175
rect 192575 113147 192609 113175
rect 192637 113147 192671 113175
rect 192699 113147 201485 113175
rect 201513 113147 201547 113175
rect 201575 113147 201609 113175
rect 201637 113147 201671 113175
rect 201699 113147 210485 113175
rect 210513 113147 210547 113175
rect 210575 113147 210609 113175
rect 210637 113147 210671 113175
rect 210699 113147 219485 113175
rect 219513 113147 219547 113175
rect 219575 113147 219609 113175
rect 219637 113147 219671 113175
rect 219699 113147 228485 113175
rect 228513 113147 228547 113175
rect 228575 113147 228609 113175
rect 228637 113147 228671 113175
rect 228699 113147 237485 113175
rect 237513 113147 237547 113175
rect 237575 113147 237609 113175
rect 237637 113147 237671 113175
rect 237699 113147 246485 113175
rect 246513 113147 246547 113175
rect 246575 113147 246609 113175
rect 246637 113147 246671 113175
rect 246699 113147 255485 113175
rect 255513 113147 255547 113175
rect 255575 113147 255609 113175
rect 255637 113147 255671 113175
rect 255699 113147 264485 113175
rect 264513 113147 264547 113175
rect 264575 113147 264609 113175
rect 264637 113147 264671 113175
rect 264699 113147 273485 113175
rect 273513 113147 273547 113175
rect 273575 113147 273609 113175
rect 273637 113147 273671 113175
rect 273699 113147 282485 113175
rect 282513 113147 282547 113175
rect 282575 113147 282609 113175
rect 282637 113147 282671 113175
rect 282699 113147 291485 113175
rect 291513 113147 291547 113175
rect 291575 113147 291609 113175
rect 291637 113147 291671 113175
rect 291699 113147 298728 113175
rect 298756 113147 298790 113175
rect 298818 113147 298852 113175
rect 298880 113147 298914 113175
rect 298942 113147 298990 113175
rect -958 113113 298990 113147
rect -958 113085 -910 113113
rect -882 113085 -848 113113
rect -820 113085 -786 113113
rect -758 113085 -724 113113
rect -696 113085 3485 113113
rect 3513 113085 3547 113113
rect 3575 113085 3609 113113
rect 3637 113085 3671 113113
rect 3699 113085 12485 113113
rect 12513 113085 12547 113113
rect 12575 113085 12609 113113
rect 12637 113085 12671 113113
rect 12699 113085 21485 113113
rect 21513 113085 21547 113113
rect 21575 113085 21609 113113
rect 21637 113085 21671 113113
rect 21699 113085 30485 113113
rect 30513 113085 30547 113113
rect 30575 113085 30609 113113
rect 30637 113085 30671 113113
rect 30699 113085 39485 113113
rect 39513 113085 39547 113113
rect 39575 113085 39609 113113
rect 39637 113085 39671 113113
rect 39699 113085 48485 113113
rect 48513 113085 48547 113113
rect 48575 113085 48609 113113
rect 48637 113085 48671 113113
rect 48699 113085 57485 113113
rect 57513 113085 57547 113113
rect 57575 113085 57609 113113
rect 57637 113085 57671 113113
rect 57699 113085 66485 113113
rect 66513 113085 66547 113113
rect 66575 113085 66609 113113
rect 66637 113085 66671 113113
rect 66699 113085 75485 113113
rect 75513 113085 75547 113113
rect 75575 113085 75609 113113
rect 75637 113085 75671 113113
rect 75699 113085 84485 113113
rect 84513 113085 84547 113113
rect 84575 113085 84609 113113
rect 84637 113085 84671 113113
rect 84699 113085 93485 113113
rect 93513 113085 93547 113113
rect 93575 113085 93609 113113
rect 93637 113085 93671 113113
rect 93699 113085 102485 113113
rect 102513 113085 102547 113113
rect 102575 113085 102609 113113
rect 102637 113085 102671 113113
rect 102699 113085 111485 113113
rect 111513 113085 111547 113113
rect 111575 113085 111609 113113
rect 111637 113085 111671 113113
rect 111699 113085 120485 113113
rect 120513 113085 120547 113113
rect 120575 113085 120609 113113
rect 120637 113085 120671 113113
rect 120699 113085 129485 113113
rect 129513 113085 129547 113113
rect 129575 113085 129609 113113
rect 129637 113085 129671 113113
rect 129699 113085 138485 113113
rect 138513 113085 138547 113113
rect 138575 113085 138609 113113
rect 138637 113085 138671 113113
rect 138699 113085 147485 113113
rect 147513 113085 147547 113113
rect 147575 113085 147609 113113
rect 147637 113085 147671 113113
rect 147699 113085 156485 113113
rect 156513 113085 156547 113113
rect 156575 113085 156609 113113
rect 156637 113085 156671 113113
rect 156699 113085 165485 113113
rect 165513 113085 165547 113113
rect 165575 113085 165609 113113
rect 165637 113085 165671 113113
rect 165699 113085 174485 113113
rect 174513 113085 174547 113113
rect 174575 113085 174609 113113
rect 174637 113085 174671 113113
rect 174699 113085 183485 113113
rect 183513 113085 183547 113113
rect 183575 113085 183609 113113
rect 183637 113085 183671 113113
rect 183699 113085 192485 113113
rect 192513 113085 192547 113113
rect 192575 113085 192609 113113
rect 192637 113085 192671 113113
rect 192699 113085 201485 113113
rect 201513 113085 201547 113113
rect 201575 113085 201609 113113
rect 201637 113085 201671 113113
rect 201699 113085 210485 113113
rect 210513 113085 210547 113113
rect 210575 113085 210609 113113
rect 210637 113085 210671 113113
rect 210699 113085 219485 113113
rect 219513 113085 219547 113113
rect 219575 113085 219609 113113
rect 219637 113085 219671 113113
rect 219699 113085 228485 113113
rect 228513 113085 228547 113113
rect 228575 113085 228609 113113
rect 228637 113085 228671 113113
rect 228699 113085 237485 113113
rect 237513 113085 237547 113113
rect 237575 113085 237609 113113
rect 237637 113085 237671 113113
rect 237699 113085 246485 113113
rect 246513 113085 246547 113113
rect 246575 113085 246609 113113
rect 246637 113085 246671 113113
rect 246699 113085 255485 113113
rect 255513 113085 255547 113113
rect 255575 113085 255609 113113
rect 255637 113085 255671 113113
rect 255699 113085 264485 113113
rect 264513 113085 264547 113113
rect 264575 113085 264609 113113
rect 264637 113085 264671 113113
rect 264699 113085 273485 113113
rect 273513 113085 273547 113113
rect 273575 113085 273609 113113
rect 273637 113085 273671 113113
rect 273699 113085 282485 113113
rect 282513 113085 282547 113113
rect 282575 113085 282609 113113
rect 282637 113085 282671 113113
rect 282699 113085 291485 113113
rect 291513 113085 291547 113113
rect 291575 113085 291609 113113
rect 291637 113085 291671 113113
rect 291699 113085 298728 113113
rect 298756 113085 298790 113113
rect 298818 113085 298852 113113
rect 298880 113085 298914 113113
rect 298942 113085 298990 113113
rect -958 113051 298990 113085
rect -958 113023 -910 113051
rect -882 113023 -848 113051
rect -820 113023 -786 113051
rect -758 113023 -724 113051
rect -696 113023 3485 113051
rect 3513 113023 3547 113051
rect 3575 113023 3609 113051
rect 3637 113023 3671 113051
rect 3699 113023 12485 113051
rect 12513 113023 12547 113051
rect 12575 113023 12609 113051
rect 12637 113023 12671 113051
rect 12699 113023 21485 113051
rect 21513 113023 21547 113051
rect 21575 113023 21609 113051
rect 21637 113023 21671 113051
rect 21699 113023 30485 113051
rect 30513 113023 30547 113051
rect 30575 113023 30609 113051
rect 30637 113023 30671 113051
rect 30699 113023 39485 113051
rect 39513 113023 39547 113051
rect 39575 113023 39609 113051
rect 39637 113023 39671 113051
rect 39699 113023 48485 113051
rect 48513 113023 48547 113051
rect 48575 113023 48609 113051
rect 48637 113023 48671 113051
rect 48699 113023 57485 113051
rect 57513 113023 57547 113051
rect 57575 113023 57609 113051
rect 57637 113023 57671 113051
rect 57699 113023 66485 113051
rect 66513 113023 66547 113051
rect 66575 113023 66609 113051
rect 66637 113023 66671 113051
rect 66699 113023 75485 113051
rect 75513 113023 75547 113051
rect 75575 113023 75609 113051
rect 75637 113023 75671 113051
rect 75699 113023 84485 113051
rect 84513 113023 84547 113051
rect 84575 113023 84609 113051
rect 84637 113023 84671 113051
rect 84699 113023 93485 113051
rect 93513 113023 93547 113051
rect 93575 113023 93609 113051
rect 93637 113023 93671 113051
rect 93699 113023 102485 113051
rect 102513 113023 102547 113051
rect 102575 113023 102609 113051
rect 102637 113023 102671 113051
rect 102699 113023 111485 113051
rect 111513 113023 111547 113051
rect 111575 113023 111609 113051
rect 111637 113023 111671 113051
rect 111699 113023 120485 113051
rect 120513 113023 120547 113051
rect 120575 113023 120609 113051
rect 120637 113023 120671 113051
rect 120699 113023 129485 113051
rect 129513 113023 129547 113051
rect 129575 113023 129609 113051
rect 129637 113023 129671 113051
rect 129699 113023 138485 113051
rect 138513 113023 138547 113051
rect 138575 113023 138609 113051
rect 138637 113023 138671 113051
rect 138699 113023 147485 113051
rect 147513 113023 147547 113051
rect 147575 113023 147609 113051
rect 147637 113023 147671 113051
rect 147699 113023 156485 113051
rect 156513 113023 156547 113051
rect 156575 113023 156609 113051
rect 156637 113023 156671 113051
rect 156699 113023 165485 113051
rect 165513 113023 165547 113051
rect 165575 113023 165609 113051
rect 165637 113023 165671 113051
rect 165699 113023 174485 113051
rect 174513 113023 174547 113051
rect 174575 113023 174609 113051
rect 174637 113023 174671 113051
rect 174699 113023 183485 113051
rect 183513 113023 183547 113051
rect 183575 113023 183609 113051
rect 183637 113023 183671 113051
rect 183699 113023 192485 113051
rect 192513 113023 192547 113051
rect 192575 113023 192609 113051
rect 192637 113023 192671 113051
rect 192699 113023 201485 113051
rect 201513 113023 201547 113051
rect 201575 113023 201609 113051
rect 201637 113023 201671 113051
rect 201699 113023 210485 113051
rect 210513 113023 210547 113051
rect 210575 113023 210609 113051
rect 210637 113023 210671 113051
rect 210699 113023 219485 113051
rect 219513 113023 219547 113051
rect 219575 113023 219609 113051
rect 219637 113023 219671 113051
rect 219699 113023 228485 113051
rect 228513 113023 228547 113051
rect 228575 113023 228609 113051
rect 228637 113023 228671 113051
rect 228699 113023 237485 113051
rect 237513 113023 237547 113051
rect 237575 113023 237609 113051
rect 237637 113023 237671 113051
rect 237699 113023 246485 113051
rect 246513 113023 246547 113051
rect 246575 113023 246609 113051
rect 246637 113023 246671 113051
rect 246699 113023 255485 113051
rect 255513 113023 255547 113051
rect 255575 113023 255609 113051
rect 255637 113023 255671 113051
rect 255699 113023 264485 113051
rect 264513 113023 264547 113051
rect 264575 113023 264609 113051
rect 264637 113023 264671 113051
rect 264699 113023 273485 113051
rect 273513 113023 273547 113051
rect 273575 113023 273609 113051
rect 273637 113023 273671 113051
rect 273699 113023 282485 113051
rect 282513 113023 282547 113051
rect 282575 113023 282609 113051
rect 282637 113023 282671 113051
rect 282699 113023 291485 113051
rect 291513 113023 291547 113051
rect 291575 113023 291609 113051
rect 291637 113023 291671 113051
rect 291699 113023 298728 113051
rect 298756 113023 298790 113051
rect 298818 113023 298852 113051
rect 298880 113023 298914 113051
rect 298942 113023 298990 113051
rect -958 112989 298990 113023
rect -958 112961 -910 112989
rect -882 112961 -848 112989
rect -820 112961 -786 112989
rect -758 112961 -724 112989
rect -696 112961 3485 112989
rect 3513 112961 3547 112989
rect 3575 112961 3609 112989
rect 3637 112961 3671 112989
rect 3699 112961 12485 112989
rect 12513 112961 12547 112989
rect 12575 112961 12609 112989
rect 12637 112961 12671 112989
rect 12699 112961 21485 112989
rect 21513 112961 21547 112989
rect 21575 112961 21609 112989
rect 21637 112961 21671 112989
rect 21699 112961 30485 112989
rect 30513 112961 30547 112989
rect 30575 112961 30609 112989
rect 30637 112961 30671 112989
rect 30699 112961 39485 112989
rect 39513 112961 39547 112989
rect 39575 112961 39609 112989
rect 39637 112961 39671 112989
rect 39699 112961 48485 112989
rect 48513 112961 48547 112989
rect 48575 112961 48609 112989
rect 48637 112961 48671 112989
rect 48699 112961 57485 112989
rect 57513 112961 57547 112989
rect 57575 112961 57609 112989
rect 57637 112961 57671 112989
rect 57699 112961 66485 112989
rect 66513 112961 66547 112989
rect 66575 112961 66609 112989
rect 66637 112961 66671 112989
rect 66699 112961 75485 112989
rect 75513 112961 75547 112989
rect 75575 112961 75609 112989
rect 75637 112961 75671 112989
rect 75699 112961 84485 112989
rect 84513 112961 84547 112989
rect 84575 112961 84609 112989
rect 84637 112961 84671 112989
rect 84699 112961 93485 112989
rect 93513 112961 93547 112989
rect 93575 112961 93609 112989
rect 93637 112961 93671 112989
rect 93699 112961 102485 112989
rect 102513 112961 102547 112989
rect 102575 112961 102609 112989
rect 102637 112961 102671 112989
rect 102699 112961 111485 112989
rect 111513 112961 111547 112989
rect 111575 112961 111609 112989
rect 111637 112961 111671 112989
rect 111699 112961 120485 112989
rect 120513 112961 120547 112989
rect 120575 112961 120609 112989
rect 120637 112961 120671 112989
rect 120699 112961 129485 112989
rect 129513 112961 129547 112989
rect 129575 112961 129609 112989
rect 129637 112961 129671 112989
rect 129699 112961 138485 112989
rect 138513 112961 138547 112989
rect 138575 112961 138609 112989
rect 138637 112961 138671 112989
rect 138699 112961 147485 112989
rect 147513 112961 147547 112989
rect 147575 112961 147609 112989
rect 147637 112961 147671 112989
rect 147699 112961 156485 112989
rect 156513 112961 156547 112989
rect 156575 112961 156609 112989
rect 156637 112961 156671 112989
rect 156699 112961 165485 112989
rect 165513 112961 165547 112989
rect 165575 112961 165609 112989
rect 165637 112961 165671 112989
rect 165699 112961 174485 112989
rect 174513 112961 174547 112989
rect 174575 112961 174609 112989
rect 174637 112961 174671 112989
rect 174699 112961 183485 112989
rect 183513 112961 183547 112989
rect 183575 112961 183609 112989
rect 183637 112961 183671 112989
rect 183699 112961 192485 112989
rect 192513 112961 192547 112989
rect 192575 112961 192609 112989
rect 192637 112961 192671 112989
rect 192699 112961 201485 112989
rect 201513 112961 201547 112989
rect 201575 112961 201609 112989
rect 201637 112961 201671 112989
rect 201699 112961 210485 112989
rect 210513 112961 210547 112989
rect 210575 112961 210609 112989
rect 210637 112961 210671 112989
rect 210699 112961 219485 112989
rect 219513 112961 219547 112989
rect 219575 112961 219609 112989
rect 219637 112961 219671 112989
rect 219699 112961 228485 112989
rect 228513 112961 228547 112989
rect 228575 112961 228609 112989
rect 228637 112961 228671 112989
rect 228699 112961 237485 112989
rect 237513 112961 237547 112989
rect 237575 112961 237609 112989
rect 237637 112961 237671 112989
rect 237699 112961 246485 112989
rect 246513 112961 246547 112989
rect 246575 112961 246609 112989
rect 246637 112961 246671 112989
rect 246699 112961 255485 112989
rect 255513 112961 255547 112989
rect 255575 112961 255609 112989
rect 255637 112961 255671 112989
rect 255699 112961 264485 112989
rect 264513 112961 264547 112989
rect 264575 112961 264609 112989
rect 264637 112961 264671 112989
rect 264699 112961 273485 112989
rect 273513 112961 273547 112989
rect 273575 112961 273609 112989
rect 273637 112961 273671 112989
rect 273699 112961 282485 112989
rect 282513 112961 282547 112989
rect 282575 112961 282609 112989
rect 282637 112961 282671 112989
rect 282699 112961 291485 112989
rect 291513 112961 291547 112989
rect 291575 112961 291609 112989
rect 291637 112961 291671 112989
rect 291699 112961 298728 112989
rect 298756 112961 298790 112989
rect 298818 112961 298852 112989
rect 298880 112961 298914 112989
rect 298942 112961 298990 112989
rect -958 112913 298990 112961
rect -958 110175 298990 110223
rect -958 110147 -430 110175
rect -402 110147 -368 110175
rect -340 110147 -306 110175
rect -278 110147 -244 110175
rect -216 110147 1625 110175
rect 1653 110147 1687 110175
rect 1715 110147 1749 110175
rect 1777 110147 1811 110175
rect 1839 110147 10625 110175
rect 10653 110147 10687 110175
rect 10715 110147 10749 110175
rect 10777 110147 10811 110175
rect 10839 110147 19625 110175
rect 19653 110147 19687 110175
rect 19715 110147 19749 110175
rect 19777 110147 19811 110175
rect 19839 110147 28625 110175
rect 28653 110147 28687 110175
rect 28715 110147 28749 110175
rect 28777 110147 28811 110175
rect 28839 110147 37625 110175
rect 37653 110147 37687 110175
rect 37715 110147 37749 110175
rect 37777 110147 37811 110175
rect 37839 110147 46625 110175
rect 46653 110147 46687 110175
rect 46715 110147 46749 110175
rect 46777 110147 46811 110175
rect 46839 110147 55625 110175
rect 55653 110147 55687 110175
rect 55715 110147 55749 110175
rect 55777 110147 55811 110175
rect 55839 110147 64625 110175
rect 64653 110147 64687 110175
rect 64715 110147 64749 110175
rect 64777 110147 64811 110175
rect 64839 110147 73625 110175
rect 73653 110147 73687 110175
rect 73715 110147 73749 110175
rect 73777 110147 73811 110175
rect 73839 110147 82625 110175
rect 82653 110147 82687 110175
rect 82715 110147 82749 110175
rect 82777 110147 82811 110175
rect 82839 110147 91625 110175
rect 91653 110147 91687 110175
rect 91715 110147 91749 110175
rect 91777 110147 91811 110175
rect 91839 110147 100625 110175
rect 100653 110147 100687 110175
rect 100715 110147 100749 110175
rect 100777 110147 100811 110175
rect 100839 110147 109625 110175
rect 109653 110147 109687 110175
rect 109715 110147 109749 110175
rect 109777 110147 109811 110175
rect 109839 110147 118625 110175
rect 118653 110147 118687 110175
rect 118715 110147 118749 110175
rect 118777 110147 118811 110175
rect 118839 110147 127625 110175
rect 127653 110147 127687 110175
rect 127715 110147 127749 110175
rect 127777 110147 127811 110175
rect 127839 110147 136625 110175
rect 136653 110147 136687 110175
rect 136715 110147 136749 110175
rect 136777 110147 136811 110175
rect 136839 110147 145625 110175
rect 145653 110147 145687 110175
rect 145715 110147 145749 110175
rect 145777 110147 145811 110175
rect 145839 110147 154625 110175
rect 154653 110147 154687 110175
rect 154715 110147 154749 110175
rect 154777 110147 154811 110175
rect 154839 110147 163625 110175
rect 163653 110147 163687 110175
rect 163715 110147 163749 110175
rect 163777 110147 163811 110175
rect 163839 110147 172625 110175
rect 172653 110147 172687 110175
rect 172715 110147 172749 110175
rect 172777 110147 172811 110175
rect 172839 110147 181625 110175
rect 181653 110147 181687 110175
rect 181715 110147 181749 110175
rect 181777 110147 181811 110175
rect 181839 110147 190625 110175
rect 190653 110147 190687 110175
rect 190715 110147 190749 110175
rect 190777 110147 190811 110175
rect 190839 110147 199625 110175
rect 199653 110147 199687 110175
rect 199715 110147 199749 110175
rect 199777 110147 199811 110175
rect 199839 110147 208625 110175
rect 208653 110147 208687 110175
rect 208715 110147 208749 110175
rect 208777 110147 208811 110175
rect 208839 110147 217625 110175
rect 217653 110147 217687 110175
rect 217715 110147 217749 110175
rect 217777 110147 217811 110175
rect 217839 110147 226625 110175
rect 226653 110147 226687 110175
rect 226715 110147 226749 110175
rect 226777 110147 226811 110175
rect 226839 110147 235625 110175
rect 235653 110147 235687 110175
rect 235715 110147 235749 110175
rect 235777 110147 235811 110175
rect 235839 110147 244625 110175
rect 244653 110147 244687 110175
rect 244715 110147 244749 110175
rect 244777 110147 244811 110175
rect 244839 110147 253625 110175
rect 253653 110147 253687 110175
rect 253715 110147 253749 110175
rect 253777 110147 253811 110175
rect 253839 110147 262625 110175
rect 262653 110147 262687 110175
rect 262715 110147 262749 110175
rect 262777 110147 262811 110175
rect 262839 110147 271625 110175
rect 271653 110147 271687 110175
rect 271715 110147 271749 110175
rect 271777 110147 271811 110175
rect 271839 110147 280625 110175
rect 280653 110147 280687 110175
rect 280715 110147 280749 110175
rect 280777 110147 280811 110175
rect 280839 110147 289625 110175
rect 289653 110147 289687 110175
rect 289715 110147 289749 110175
rect 289777 110147 289811 110175
rect 289839 110147 298248 110175
rect 298276 110147 298310 110175
rect 298338 110147 298372 110175
rect 298400 110147 298434 110175
rect 298462 110147 298990 110175
rect -958 110113 298990 110147
rect -958 110085 -430 110113
rect -402 110085 -368 110113
rect -340 110085 -306 110113
rect -278 110085 -244 110113
rect -216 110085 1625 110113
rect 1653 110085 1687 110113
rect 1715 110085 1749 110113
rect 1777 110085 1811 110113
rect 1839 110085 10625 110113
rect 10653 110085 10687 110113
rect 10715 110085 10749 110113
rect 10777 110085 10811 110113
rect 10839 110085 19625 110113
rect 19653 110085 19687 110113
rect 19715 110085 19749 110113
rect 19777 110085 19811 110113
rect 19839 110085 28625 110113
rect 28653 110085 28687 110113
rect 28715 110085 28749 110113
rect 28777 110085 28811 110113
rect 28839 110085 37625 110113
rect 37653 110085 37687 110113
rect 37715 110085 37749 110113
rect 37777 110085 37811 110113
rect 37839 110085 46625 110113
rect 46653 110085 46687 110113
rect 46715 110085 46749 110113
rect 46777 110085 46811 110113
rect 46839 110085 55625 110113
rect 55653 110085 55687 110113
rect 55715 110085 55749 110113
rect 55777 110085 55811 110113
rect 55839 110085 64625 110113
rect 64653 110085 64687 110113
rect 64715 110085 64749 110113
rect 64777 110085 64811 110113
rect 64839 110085 73625 110113
rect 73653 110085 73687 110113
rect 73715 110085 73749 110113
rect 73777 110085 73811 110113
rect 73839 110085 82625 110113
rect 82653 110085 82687 110113
rect 82715 110085 82749 110113
rect 82777 110085 82811 110113
rect 82839 110085 91625 110113
rect 91653 110085 91687 110113
rect 91715 110085 91749 110113
rect 91777 110085 91811 110113
rect 91839 110085 100625 110113
rect 100653 110085 100687 110113
rect 100715 110085 100749 110113
rect 100777 110085 100811 110113
rect 100839 110085 109625 110113
rect 109653 110085 109687 110113
rect 109715 110085 109749 110113
rect 109777 110085 109811 110113
rect 109839 110085 118625 110113
rect 118653 110085 118687 110113
rect 118715 110085 118749 110113
rect 118777 110085 118811 110113
rect 118839 110085 127625 110113
rect 127653 110085 127687 110113
rect 127715 110085 127749 110113
rect 127777 110085 127811 110113
rect 127839 110085 136625 110113
rect 136653 110085 136687 110113
rect 136715 110085 136749 110113
rect 136777 110085 136811 110113
rect 136839 110085 145625 110113
rect 145653 110085 145687 110113
rect 145715 110085 145749 110113
rect 145777 110085 145811 110113
rect 145839 110085 154625 110113
rect 154653 110085 154687 110113
rect 154715 110085 154749 110113
rect 154777 110085 154811 110113
rect 154839 110085 163625 110113
rect 163653 110085 163687 110113
rect 163715 110085 163749 110113
rect 163777 110085 163811 110113
rect 163839 110085 172625 110113
rect 172653 110085 172687 110113
rect 172715 110085 172749 110113
rect 172777 110085 172811 110113
rect 172839 110085 181625 110113
rect 181653 110085 181687 110113
rect 181715 110085 181749 110113
rect 181777 110085 181811 110113
rect 181839 110085 190625 110113
rect 190653 110085 190687 110113
rect 190715 110085 190749 110113
rect 190777 110085 190811 110113
rect 190839 110085 199625 110113
rect 199653 110085 199687 110113
rect 199715 110085 199749 110113
rect 199777 110085 199811 110113
rect 199839 110085 208625 110113
rect 208653 110085 208687 110113
rect 208715 110085 208749 110113
rect 208777 110085 208811 110113
rect 208839 110085 217625 110113
rect 217653 110085 217687 110113
rect 217715 110085 217749 110113
rect 217777 110085 217811 110113
rect 217839 110085 226625 110113
rect 226653 110085 226687 110113
rect 226715 110085 226749 110113
rect 226777 110085 226811 110113
rect 226839 110085 235625 110113
rect 235653 110085 235687 110113
rect 235715 110085 235749 110113
rect 235777 110085 235811 110113
rect 235839 110085 244625 110113
rect 244653 110085 244687 110113
rect 244715 110085 244749 110113
rect 244777 110085 244811 110113
rect 244839 110085 253625 110113
rect 253653 110085 253687 110113
rect 253715 110085 253749 110113
rect 253777 110085 253811 110113
rect 253839 110085 262625 110113
rect 262653 110085 262687 110113
rect 262715 110085 262749 110113
rect 262777 110085 262811 110113
rect 262839 110085 271625 110113
rect 271653 110085 271687 110113
rect 271715 110085 271749 110113
rect 271777 110085 271811 110113
rect 271839 110085 280625 110113
rect 280653 110085 280687 110113
rect 280715 110085 280749 110113
rect 280777 110085 280811 110113
rect 280839 110085 289625 110113
rect 289653 110085 289687 110113
rect 289715 110085 289749 110113
rect 289777 110085 289811 110113
rect 289839 110085 298248 110113
rect 298276 110085 298310 110113
rect 298338 110085 298372 110113
rect 298400 110085 298434 110113
rect 298462 110085 298990 110113
rect -958 110051 298990 110085
rect -958 110023 -430 110051
rect -402 110023 -368 110051
rect -340 110023 -306 110051
rect -278 110023 -244 110051
rect -216 110023 1625 110051
rect 1653 110023 1687 110051
rect 1715 110023 1749 110051
rect 1777 110023 1811 110051
rect 1839 110023 10625 110051
rect 10653 110023 10687 110051
rect 10715 110023 10749 110051
rect 10777 110023 10811 110051
rect 10839 110023 19625 110051
rect 19653 110023 19687 110051
rect 19715 110023 19749 110051
rect 19777 110023 19811 110051
rect 19839 110023 28625 110051
rect 28653 110023 28687 110051
rect 28715 110023 28749 110051
rect 28777 110023 28811 110051
rect 28839 110023 37625 110051
rect 37653 110023 37687 110051
rect 37715 110023 37749 110051
rect 37777 110023 37811 110051
rect 37839 110023 46625 110051
rect 46653 110023 46687 110051
rect 46715 110023 46749 110051
rect 46777 110023 46811 110051
rect 46839 110023 55625 110051
rect 55653 110023 55687 110051
rect 55715 110023 55749 110051
rect 55777 110023 55811 110051
rect 55839 110023 64625 110051
rect 64653 110023 64687 110051
rect 64715 110023 64749 110051
rect 64777 110023 64811 110051
rect 64839 110023 73625 110051
rect 73653 110023 73687 110051
rect 73715 110023 73749 110051
rect 73777 110023 73811 110051
rect 73839 110023 82625 110051
rect 82653 110023 82687 110051
rect 82715 110023 82749 110051
rect 82777 110023 82811 110051
rect 82839 110023 91625 110051
rect 91653 110023 91687 110051
rect 91715 110023 91749 110051
rect 91777 110023 91811 110051
rect 91839 110023 100625 110051
rect 100653 110023 100687 110051
rect 100715 110023 100749 110051
rect 100777 110023 100811 110051
rect 100839 110023 109625 110051
rect 109653 110023 109687 110051
rect 109715 110023 109749 110051
rect 109777 110023 109811 110051
rect 109839 110023 118625 110051
rect 118653 110023 118687 110051
rect 118715 110023 118749 110051
rect 118777 110023 118811 110051
rect 118839 110023 127625 110051
rect 127653 110023 127687 110051
rect 127715 110023 127749 110051
rect 127777 110023 127811 110051
rect 127839 110023 136625 110051
rect 136653 110023 136687 110051
rect 136715 110023 136749 110051
rect 136777 110023 136811 110051
rect 136839 110023 145625 110051
rect 145653 110023 145687 110051
rect 145715 110023 145749 110051
rect 145777 110023 145811 110051
rect 145839 110023 154625 110051
rect 154653 110023 154687 110051
rect 154715 110023 154749 110051
rect 154777 110023 154811 110051
rect 154839 110023 163625 110051
rect 163653 110023 163687 110051
rect 163715 110023 163749 110051
rect 163777 110023 163811 110051
rect 163839 110023 172625 110051
rect 172653 110023 172687 110051
rect 172715 110023 172749 110051
rect 172777 110023 172811 110051
rect 172839 110023 181625 110051
rect 181653 110023 181687 110051
rect 181715 110023 181749 110051
rect 181777 110023 181811 110051
rect 181839 110023 190625 110051
rect 190653 110023 190687 110051
rect 190715 110023 190749 110051
rect 190777 110023 190811 110051
rect 190839 110023 199625 110051
rect 199653 110023 199687 110051
rect 199715 110023 199749 110051
rect 199777 110023 199811 110051
rect 199839 110023 208625 110051
rect 208653 110023 208687 110051
rect 208715 110023 208749 110051
rect 208777 110023 208811 110051
rect 208839 110023 217625 110051
rect 217653 110023 217687 110051
rect 217715 110023 217749 110051
rect 217777 110023 217811 110051
rect 217839 110023 226625 110051
rect 226653 110023 226687 110051
rect 226715 110023 226749 110051
rect 226777 110023 226811 110051
rect 226839 110023 235625 110051
rect 235653 110023 235687 110051
rect 235715 110023 235749 110051
rect 235777 110023 235811 110051
rect 235839 110023 244625 110051
rect 244653 110023 244687 110051
rect 244715 110023 244749 110051
rect 244777 110023 244811 110051
rect 244839 110023 253625 110051
rect 253653 110023 253687 110051
rect 253715 110023 253749 110051
rect 253777 110023 253811 110051
rect 253839 110023 262625 110051
rect 262653 110023 262687 110051
rect 262715 110023 262749 110051
rect 262777 110023 262811 110051
rect 262839 110023 271625 110051
rect 271653 110023 271687 110051
rect 271715 110023 271749 110051
rect 271777 110023 271811 110051
rect 271839 110023 280625 110051
rect 280653 110023 280687 110051
rect 280715 110023 280749 110051
rect 280777 110023 280811 110051
rect 280839 110023 289625 110051
rect 289653 110023 289687 110051
rect 289715 110023 289749 110051
rect 289777 110023 289811 110051
rect 289839 110023 298248 110051
rect 298276 110023 298310 110051
rect 298338 110023 298372 110051
rect 298400 110023 298434 110051
rect 298462 110023 298990 110051
rect -958 109989 298990 110023
rect -958 109961 -430 109989
rect -402 109961 -368 109989
rect -340 109961 -306 109989
rect -278 109961 -244 109989
rect -216 109961 1625 109989
rect 1653 109961 1687 109989
rect 1715 109961 1749 109989
rect 1777 109961 1811 109989
rect 1839 109961 10625 109989
rect 10653 109961 10687 109989
rect 10715 109961 10749 109989
rect 10777 109961 10811 109989
rect 10839 109961 19625 109989
rect 19653 109961 19687 109989
rect 19715 109961 19749 109989
rect 19777 109961 19811 109989
rect 19839 109961 28625 109989
rect 28653 109961 28687 109989
rect 28715 109961 28749 109989
rect 28777 109961 28811 109989
rect 28839 109961 37625 109989
rect 37653 109961 37687 109989
rect 37715 109961 37749 109989
rect 37777 109961 37811 109989
rect 37839 109961 46625 109989
rect 46653 109961 46687 109989
rect 46715 109961 46749 109989
rect 46777 109961 46811 109989
rect 46839 109961 55625 109989
rect 55653 109961 55687 109989
rect 55715 109961 55749 109989
rect 55777 109961 55811 109989
rect 55839 109961 64625 109989
rect 64653 109961 64687 109989
rect 64715 109961 64749 109989
rect 64777 109961 64811 109989
rect 64839 109961 73625 109989
rect 73653 109961 73687 109989
rect 73715 109961 73749 109989
rect 73777 109961 73811 109989
rect 73839 109961 82625 109989
rect 82653 109961 82687 109989
rect 82715 109961 82749 109989
rect 82777 109961 82811 109989
rect 82839 109961 91625 109989
rect 91653 109961 91687 109989
rect 91715 109961 91749 109989
rect 91777 109961 91811 109989
rect 91839 109961 100625 109989
rect 100653 109961 100687 109989
rect 100715 109961 100749 109989
rect 100777 109961 100811 109989
rect 100839 109961 109625 109989
rect 109653 109961 109687 109989
rect 109715 109961 109749 109989
rect 109777 109961 109811 109989
rect 109839 109961 118625 109989
rect 118653 109961 118687 109989
rect 118715 109961 118749 109989
rect 118777 109961 118811 109989
rect 118839 109961 127625 109989
rect 127653 109961 127687 109989
rect 127715 109961 127749 109989
rect 127777 109961 127811 109989
rect 127839 109961 136625 109989
rect 136653 109961 136687 109989
rect 136715 109961 136749 109989
rect 136777 109961 136811 109989
rect 136839 109961 145625 109989
rect 145653 109961 145687 109989
rect 145715 109961 145749 109989
rect 145777 109961 145811 109989
rect 145839 109961 154625 109989
rect 154653 109961 154687 109989
rect 154715 109961 154749 109989
rect 154777 109961 154811 109989
rect 154839 109961 163625 109989
rect 163653 109961 163687 109989
rect 163715 109961 163749 109989
rect 163777 109961 163811 109989
rect 163839 109961 172625 109989
rect 172653 109961 172687 109989
rect 172715 109961 172749 109989
rect 172777 109961 172811 109989
rect 172839 109961 181625 109989
rect 181653 109961 181687 109989
rect 181715 109961 181749 109989
rect 181777 109961 181811 109989
rect 181839 109961 190625 109989
rect 190653 109961 190687 109989
rect 190715 109961 190749 109989
rect 190777 109961 190811 109989
rect 190839 109961 199625 109989
rect 199653 109961 199687 109989
rect 199715 109961 199749 109989
rect 199777 109961 199811 109989
rect 199839 109961 208625 109989
rect 208653 109961 208687 109989
rect 208715 109961 208749 109989
rect 208777 109961 208811 109989
rect 208839 109961 217625 109989
rect 217653 109961 217687 109989
rect 217715 109961 217749 109989
rect 217777 109961 217811 109989
rect 217839 109961 226625 109989
rect 226653 109961 226687 109989
rect 226715 109961 226749 109989
rect 226777 109961 226811 109989
rect 226839 109961 235625 109989
rect 235653 109961 235687 109989
rect 235715 109961 235749 109989
rect 235777 109961 235811 109989
rect 235839 109961 244625 109989
rect 244653 109961 244687 109989
rect 244715 109961 244749 109989
rect 244777 109961 244811 109989
rect 244839 109961 253625 109989
rect 253653 109961 253687 109989
rect 253715 109961 253749 109989
rect 253777 109961 253811 109989
rect 253839 109961 262625 109989
rect 262653 109961 262687 109989
rect 262715 109961 262749 109989
rect 262777 109961 262811 109989
rect 262839 109961 271625 109989
rect 271653 109961 271687 109989
rect 271715 109961 271749 109989
rect 271777 109961 271811 109989
rect 271839 109961 280625 109989
rect 280653 109961 280687 109989
rect 280715 109961 280749 109989
rect 280777 109961 280811 109989
rect 280839 109961 289625 109989
rect 289653 109961 289687 109989
rect 289715 109961 289749 109989
rect 289777 109961 289811 109989
rect 289839 109961 298248 109989
rect 298276 109961 298310 109989
rect 298338 109961 298372 109989
rect 298400 109961 298434 109989
rect 298462 109961 298990 109989
rect -958 109913 298990 109961
rect -958 104175 298990 104223
rect -958 104147 -910 104175
rect -882 104147 -848 104175
rect -820 104147 -786 104175
rect -758 104147 -724 104175
rect -696 104147 3485 104175
rect 3513 104147 3547 104175
rect 3575 104147 3609 104175
rect 3637 104147 3671 104175
rect 3699 104147 12485 104175
rect 12513 104147 12547 104175
rect 12575 104147 12609 104175
rect 12637 104147 12671 104175
rect 12699 104147 21485 104175
rect 21513 104147 21547 104175
rect 21575 104147 21609 104175
rect 21637 104147 21671 104175
rect 21699 104147 30485 104175
rect 30513 104147 30547 104175
rect 30575 104147 30609 104175
rect 30637 104147 30671 104175
rect 30699 104147 39485 104175
rect 39513 104147 39547 104175
rect 39575 104147 39609 104175
rect 39637 104147 39671 104175
rect 39699 104147 48485 104175
rect 48513 104147 48547 104175
rect 48575 104147 48609 104175
rect 48637 104147 48671 104175
rect 48699 104147 54509 104175
rect 54537 104147 54571 104175
rect 54599 104147 57485 104175
rect 57513 104147 57547 104175
rect 57575 104147 57609 104175
rect 57637 104147 57671 104175
rect 57699 104147 59009 104175
rect 59037 104147 59071 104175
rect 59099 104147 63509 104175
rect 63537 104147 63571 104175
rect 63599 104147 66485 104175
rect 66513 104147 66547 104175
rect 66575 104147 66609 104175
rect 66637 104147 66671 104175
rect 66699 104147 68009 104175
rect 68037 104147 68071 104175
rect 68099 104147 72509 104175
rect 72537 104147 72571 104175
rect 72599 104147 75485 104175
rect 75513 104147 75547 104175
rect 75575 104147 75609 104175
rect 75637 104147 75671 104175
rect 75699 104147 77009 104175
rect 77037 104147 77071 104175
rect 77099 104147 81509 104175
rect 81537 104147 81571 104175
rect 81599 104147 84485 104175
rect 84513 104147 84547 104175
rect 84575 104147 84609 104175
rect 84637 104147 84671 104175
rect 84699 104147 86009 104175
rect 86037 104147 86071 104175
rect 86099 104147 90509 104175
rect 90537 104147 90571 104175
rect 90599 104147 93485 104175
rect 93513 104147 93547 104175
rect 93575 104147 93609 104175
rect 93637 104147 93671 104175
rect 93699 104147 95009 104175
rect 95037 104147 95071 104175
rect 95099 104147 99509 104175
rect 99537 104147 99571 104175
rect 99599 104147 102485 104175
rect 102513 104147 102547 104175
rect 102575 104147 102609 104175
rect 102637 104147 102671 104175
rect 102699 104147 104009 104175
rect 104037 104147 104071 104175
rect 104099 104147 108509 104175
rect 108537 104147 108571 104175
rect 108599 104147 111485 104175
rect 111513 104147 111547 104175
rect 111575 104147 111609 104175
rect 111637 104147 111671 104175
rect 111699 104147 113009 104175
rect 113037 104147 113071 104175
rect 113099 104147 117509 104175
rect 117537 104147 117571 104175
rect 117599 104147 120485 104175
rect 120513 104147 120547 104175
rect 120575 104147 120609 104175
rect 120637 104147 120671 104175
rect 120699 104147 129485 104175
rect 129513 104147 129547 104175
rect 129575 104147 129609 104175
rect 129637 104147 129671 104175
rect 129699 104147 138485 104175
rect 138513 104147 138547 104175
rect 138575 104147 138609 104175
rect 138637 104147 138671 104175
rect 138699 104147 147485 104175
rect 147513 104147 147547 104175
rect 147575 104147 147609 104175
rect 147637 104147 147671 104175
rect 147699 104147 156485 104175
rect 156513 104147 156547 104175
rect 156575 104147 156609 104175
rect 156637 104147 156671 104175
rect 156699 104147 165485 104175
rect 165513 104147 165547 104175
rect 165575 104147 165609 104175
rect 165637 104147 165671 104175
rect 165699 104147 174485 104175
rect 174513 104147 174547 104175
rect 174575 104147 174609 104175
rect 174637 104147 174671 104175
rect 174699 104147 183485 104175
rect 183513 104147 183547 104175
rect 183575 104147 183609 104175
rect 183637 104147 183671 104175
rect 183699 104147 192485 104175
rect 192513 104147 192547 104175
rect 192575 104147 192609 104175
rect 192637 104147 192671 104175
rect 192699 104147 201485 104175
rect 201513 104147 201547 104175
rect 201575 104147 201609 104175
rect 201637 104147 201671 104175
rect 201699 104147 210485 104175
rect 210513 104147 210547 104175
rect 210575 104147 210609 104175
rect 210637 104147 210671 104175
rect 210699 104147 219485 104175
rect 219513 104147 219547 104175
rect 219575 104147 219609 104175
rect 219637 104147 219671 104175
rect 219699 104147 228485 104175
rect 228513 104147 228547 104175
rect 228575 104147 228609 104175
rect 228637 104147 228671 104175
rect 228699 104147 237485 104175
rect 237513 104147 237547 104175
rect 237575 104147 237609 104175
rect 237637 104147 237671 104175
rect 237699 104147 246485 104175
rect 246513 104147 246547 104175
rect 246575 104147 246609 104175
rect 246637 104147 246671 104175
rect 246699 104147 255485 104175
rect 255513 104147 255547 104175
rect 255575 104147 255609 104175
rect 255637 104147 255671 104175
rect 255699 104147 264485 104175
rect 264513 104147 264547 104175
rect 264575 104147 264609 104175
rect 264637 104147 264671 104175
rect 264699 104147 273485 104175
rect 273513 104147 273547 104175
rect 273575 104147 273609 104175
rect 273637 104147 273671 104175
rect 273699 104147 282485 104175
rect 282513 104147 282547 104175
rect 282575 104147 282609 104175
rect 282637 104147 282671 104175
rect 282699 104147 291485 104175
rect 291513 104147 291547 104175
rect 291575 104147 291609 104175
rect 291637 104147 291671 104175
rect 291699 104147 298728 104175
rect 298756 104147 298790 104175
rect 298818 104147 298852 104175
rect 298880 104147 298914 104175
rect 298942 104147 298990 104175
rect -958 104113 298990 104147
rect -958 104085 -910 104113
rect -882 104085 -848 104113
rect -820 104085 -786 104113
rect -758 104085 -724 104113
rect -696 104085 3485 104113
rect 3513 104085 3547 104113
rect 3575 104085 3609 104113
rect 3637 104085 3671 104113
rect 3699 104085 12485 104113
rect 12513 104085 12547 104113
rect 12575 104085 12609 104113
rect 12637 104085 12671 104113
rect 12699 104085 21485 104113
rect 21513 104085 21547 104113
rect 21575 104085 21609 104113
rect 21637 104085 21671 104113
rect 21699 104085 30485 104113
rect 30513 104085 30547 104113
rect 30575 104085 30609 104113
rect 30637 104085 30671 104113
rect 30699 104085 39485 104113
rect 39513 104085 39547 104113
rect 39575 104085 39609 104113
rect 39637 104085 39671 104113
rect 39699 104085 48485 104113
rect 48513 104085 48547 104113
rect 48575 104085 48609 104113
rect 48637 104085 48671 104113
rect 48699 104085 54509 104113
rect 54537 104085 54571 104113
rect 54599 104085 57485 104113
rect 57513 104085 57547 104113
rect 57575 104085 57609 104113
rect 57637 104085 57671 104113
rect 57699 104085 59009 104113
rect 59037 104085 59071 104113
rect 59099 104085 63509 104113
rect 63537 104085 63571 104113
rect 63599 104085 66485 104113
rect 66513 104085 66547 104113
rect 66575 104085 66609 104113
rect 66637 104085 66671 104113
rect 66699 104085 68009 104113
rect 68037 104085 68071 104113
rect 68099 104085 72509 104113
rect 72537 104085 72571 104113
rect 72599 104085 75485 104113
rect 75513 104085 75547 104113
rect 75575 104085 75609 104113
rect 75637 104085 75671 104113
rect 75699 104085 77009 104113
rect 77037 104085 77071 104113
rect 77099 104085 81509 104113
rect 81537 104085 81571 104113
rect 81599 104085 84485 104113
rect 84513 104085 84547 104113
rect 84575 104085 84609 104113
rect 84637 104085 84671 104113
rect 84699 104085 86009 104113
rect 86037 104085 86071 104113
rect 86099 104085 90509 104113
rect 90537 104085 90571 104113
rect 90599 104085 93485 104113
rect 93513 104085 93547 104113
rect 93575 104085 93609 104113
rect 93637 104085 93671 104113
rect 93699 104085 95009 104113
rect 95037 104085 95071 104113
rect 95099 104085 99509 104113
rect 99537 104085 99571 104113
rect 99599 104085 102485 104113
rect 102513 104085 102547 104113
rect 102575 104085 102609 104113
rect 102637 104085 102671 104113
rect 102699 104085 104009 104113
rect 104037 104085 104071 104113
rect 104099 104085 108509 104113
rect 108537 104085 108571 104113
rect 108599 104085 111485 104113
rect 111513 104085 111547 104113
rect 111575 104085 111609 104113
rect 111637 104085 111671 104113
rect 111699 104085 113009 104113
rect 113037 104085 113071 104113
rect 113099 104085 117509 104113
rect 117537 104085 117571 104113
rect 117599 104085 120485 104113
rect 120513 104085 120547 104113
rect 120575 104085 120609 104113
rect 120637 104085 120671 104113
rect 120699 104085 129485 104113
rect 129513 104085 129547 104113
rect 129575 104085 129609 104113
rect 129637 104085 129671 104113
rect 129699 104085 138485 104113
rect 138513 104085 138547 104113
rect 138575 104085 138609 104113
rect 138637 104085 138671 104113
rect 138699 104085 147485 104113
rect 147513 104085 147547 104113
rect 147575 104085 147609 104113
rect 147637 104085 147671 104113
rect 147699 104085 156485 104113
rect 156513 104085 156547 104113
rect 156575 104085 156609 104113
rect 156637 104085 156671 104113
rect 156699 104085 165485 104113
rect 165513 104085 165547 104113
rect 165575 104085 165609 104113
rect 165637 104085 165671 104113
rect 165699 104085 174485 104113
rect 174513 104085 174547 104113
rect 174575 104085 174609 104113
rect 174637 104085 174671 104113
rect 174699 104085 183485 104113
rect 183513 104085 183547 104113
rect 183575 104085 183609 104113
rect 183637 104085 183671 104113
rect 183699 104085 192485 104113
rect 192513 104085 192547 104113
rect 192575 104085 192609 104113
rect 192637 104085 192671 104113
rect 192699 104085 201485 104113
rect 201513 104085 201547 104113
rect 201575 104085 201609 104113
rect 201637 104085 201671 104113
rect 201699 104085 210485 104113
rect 210513 104085 210547 104113
rect 210575 104085 210609 104113
rect 210637 104085 210671 104113
rect 210699 104085 219485 104113
rect 219513 104085 219547 104113
rect 219575 104085 219609 104113
rect 219637 104085 219671 104113
rect 219699 104085 228485 104113
rect 228513 104085 228547 104113
rect 228575 104085 228609 104113
rect 228637 104085 228671 104113
rect 228699 104085 237485 104113
rect 237513 104085 237547 104113
rect 237575 104085 237609 104113
rect 237637 104085 237671 104113
rect 237699 104085 246485 104113
rect 246513 104085 246547 104113
rect 246575 104085 246609 104113
rect 246637 104085 246671 104113
rect 246699 104085 255485 104113
rect 255513 104085 255547 104113
rect 255575 104085 255609 104113
rect 255637 104085 255671 104113
rect 255699 104085 264485 104113
rect 264513 104085 264547 104113
rect 264575 104085 264609 104113
rect 264637 104085 264671 104113
rect 264699 104085 273485 104113
rect 273513 104085 273547 104113
rect 273575 104085 273609 104113
rect 273637 104085 273671 104113
rect 273699 104085 282485 104113
rect 282513 104085 282547 104113
rect 282575 104085 282609 104113
rect 282637 104085 282671 104113
rect 282699 104085 291485 104113
rect 291513 104085 291547 104113
rect 291575 104085 291609 104113
rect 291637 104085 291671 104113
rect 291699 104085 298728 104113
rect 298756 104085 298790 104113
rect 298818 104085 298852 104113
rect 298880 104085 298914 104113
rect 298942 104085 298990 104113
rect -958 104051 298990 104085
rect -958 104023 -910 104051
rect -882 104023 -848 104051
rect -820 104023 -786 104051
rect -758 104023 -724 104051
rect -696 104023 3485 104051
rect 3513 104023 3547 104051
rect 3575 104023 3609 104051
rect 3637 104023 3671 104051
rect 3699 104023 12485 104051
rect 12513 104023 12547 104051
rect 12575 104023 12609 104051
rect 12637 104023 12671 104051
rect 12699 104023 21485 104051
rect 21513 104023 21547 104051
rect 21575 104023 21609 104051
rect 21637 104023 21671 104051
rect 21699 104023 30485 104051
rect 30513 104023 30547 104051
rect 30575 104023 30609 104051
rect 30637 104023 30671 104051
rect 30699 104023 39485 104051
rect 39513 104023 39547 104051
rect 39575 104023 39609 104051
rect 39637 104023 39671 104051
rect 39699 104023 48485 104051
rect 48513 104023 48547 104051
rect 48575 104023 48609 104051
rect 48637 104023 48671 104051
rect 48699 104023 54509 104051
rect 54537 104023 54571 104051
rect 54599 104023 57485 104051
rect 57513 104023 57547 104051
rect 57575 104023 57609 104051
rect 57637 104023 57671 104051
rect 57699 104023 59009 104051
rect 59037 104023 59071 104051
rect 59099 104023 63509 104051
rect 63537 104023 63571 104051
rect 63599 104023 66485 104051
rect 66513 104023 66547 104051
rect 66575 104023 66609 104051
rect 66637 104023 66671 104051
rect 66699 104023 68009 104051
rect 68037 104023 68071 104051
rect 68099 104023 72509 104051
rect 72537 104023 72571 104051
rect 72599 104023 75485 104051
rect 75513 104023 75547 104051
rect 75575 104023 75609 104051
rect 75637 104023 75671 104051
rect 75699 104023 77009 104051
rect 77037 104023 77071 104051
rect 77099 104023 81509 104051
rect 81537 104023 81571 104051
rect 81599 104023 84485 104051
rect 84513 104023 84547 104051
rect 84575 104023 84609 104051
rect 84637 104023 84671 104051
rect 84699 104023 86009 104051
rect 86037 104023 86071 104051
rect 86099 104023 90509 104051
rect 90537 104023 90571 104051
rect 90599 104023 93485 104051
rect 93513 104023 93547 104051
rect 93575 104023 93609 104051
rect 93637 104023 93671 104051
rect 93699 104023 95009 104051
rect 95037 104023 95071 104051
rect 95099 104023 99509 104051
rect 99537 104023 99571 104051
rect 99599 104023 102485 104051
rect 102513 104023 102547 104051
rect 102575 104023 102609 104051
rect 102637 104023 102671 104051
rect 102699 104023 104009 104051
rect 104037 104023 104071 104051
rect 104099 104023 108509 104051
rect 108537 104023 108571 104051
rect 108599 104023 111485 104051
rect 111513 104023 111547 104051
rect 111575 104023 111609 104051
rect 111637 104023 111671 104051
rect 111699 104023 113009 104051
rect 113037 104023 113071 104051
rect 113099 104023 117509 104051
rect 117537 104023 117571 104051
rect 117599 104023 120485 104051
rect 120513 104023 120547 104051
rect 120575 104023 120609 104051
rect 120637 104023 120671 104051
rect 120699 104023 129485 104051
rect 129513 104023 129547 104051
rect 129575 104023 129609 104051
rect 129637 104023 129671 104051
rect 129699 104023 138485 104051
rect 138513 104023 138547 104051
rect 138575 104023 138609 104051
rect 138637 104023 138671 104051
rect 138699 104023 147485 104051
rect 147513 104023 147547 104051
rect 147575 104023 147609 104051
rect 147637 104023 147671 104051
rect 147699 104023 156485 104051
rect 156513 104023 156547 104051
rect 156575 104023 156609 104051
rect 156637 104023 156671 104051
rect 156699 104023 165485 104051
rect 165513 104023 165547 104051
rect 165575 104023 165609 104051
rect 165637 104023 165671 104051
rect 165699 104023 174485 104051
rect 174513 104023 174547 104051
rect 174575 104023 174609 104051
rect 174637 104023 174671 104051
rect 174699 104023 183485 104051
rect 183513 104023 183547 104051
rect 183575 104023 183609 104051
rect 183637 104023 183671 104051
rect 183699 104023 192485 104051
rect 192513 104023 192547 104051
rect 192575 104023 192609 104051
rect 192637 104023 192671 104051
rect 192699 104023 201485 104051
rect 201513 104023 201547 104051
rect 201575 104023 201609 104051
rect 201637 104023 201671 104051
rect 201699 104023 210485 104051
rect 210513 104023 210547 104051
rect 210575 104023 210609 104051
rect 210637 104023 210671 104051
rect 210699 104023 219485 104051
rect 219513 104023 219547 104051
rect 219575 104023 219609 104051
rect 219637 104023 219671 104051
rect 219699 104023 228485 104051
rect 228513 104023 228547 104051
rect 228575 104023 228609 104051
rect 228637 104023 228671 104051
rect 228699 104023 237485 104051
rect 237513 104023 237547 104051
rect 237575 104023 237609 104051
rect 237637 104023 237671 104051
rect 237699 104023 246485 104051
rect 246513 104023 246547 104051
rect 246575 104023 246609 104051
rect 246637 104023 246671 104051
rect 246699 104023 255485 104051
rect 255513 104023 255547 104051
rect 255575 104023 255609 104051
rect 255637 104023 255671 104051
rect 255699 104023 264485 104051
rect 264513 104023 264547 104051
rect 264575 104023 264609 104051
rect 264637 104023 264671 104051
rect 264699 104023 273485 104051
rect 273513 104023 273547 104051
rect 273575 104023 273609 104051
rect 273637 104023 273671 104051
rect 273699 104023 282485 104051
rect 282513 104023 282547 104051
rect 282575 104023 282609 104051
rect 282637 104023 282671 104051
rect 282699 104023 291485 104051
rect 291513 104023 291547 104051
rect 291575 104023 291609 104051
rect 291637 104023 291671 104051
rect 291699 104023 298728 104051
rect 298756 104023 298790 104051
rect 298818 104023 298852 104051
rect 298880 104023 298914 104051
rect 298942 104023 298990 104051
rect -958 103989 298990 104023
rect -958 103961 -910 103989
rect -882 103961 -848 103989
rect -820 103961 -786 103989
rect -758 103961 -724 103989
rect -696 103961 3485 103989
rect 3513 103961 3547 103989
rect 3575 103961 3609 103989
rect 3637 103961 3671 103989
rect 3699 103961 12485 103989
rect 12513 103961 12547 103989
rect 12575 103961 12609 103989
rect 12637 103961 12671 103989
rect 12699 103961 21485 103989
rect 21513 103961 21547 103989
rect 21575 103961 21609 103989
rect 21637 103961 21671 103989
rect 21699 103961 30485 103989
rect 30513 103961 30547 103989
rect 30575 103961 30609 103989
rect 30637 103961 30671 103989
rect 30699 103961 39485 103989
rect 39513 103961 39547 103989
rect 39575 103961 39609 103989
rect 39637 103961 39671 103989
rect 39699 103961 48485 103989
rect 48513 103961 48547 103989
rect 48575 103961 48609 103989
rect 48637 103961 48671 103989
rect 48699 103961 54509 103989
rect 54537 103961 54571 103989
rect 54599 103961 57485 103989
rect 57513 103961 57547 103989
rect 57575 103961 57609 103989
rect 57637 103961 57671 103989
rect 57699 103961 59009 103989
rect 59037 103961 59071 103989
rect 59099 103961 63509 103989
rect 63537 103961 63571 103989
rect 63599 103961 66485 103989
rect 66513 103961 66547 103989
rect 66575 103961 66609 103989
rect 66637 103961 66671 103989
rect 66699 103961 68009 103989
rect 68037 103961 68071 103989
rect 68099 103961 72509 103989
rect 72537 103961 72571 103989
rect 72599 103961 75485 103989
rect 75513 103961 75547 103989
rect 75575 103961 75609 103989
rect 75637 103961 75671 103989
rect 75699 103961 77009 103989
rect 77037 103961 77071 103989
rect 77099 103961 81509 103989
rect 81537 103961 81571 103989
rect 81599 103961 84485 103989
rect 84513 103961 84547 103989
rect 84575 103961 84609 103989
rect 84637 103961 84671 103989
rect 84699 103961 86009 103989
rect 86037 103961 86071 103989
rect 86099 103961 90509 103989
rect 90537 103961 90571 103989
rect 90599 103961 93485 103989
rect 93513 103961 93547 103989
rect 93575 103961 93609 103989
rect 93637 103961 93671 103989
rect 93699 103961 95009 103989
rect 95037 103961 95071 103989
rect 95099 103961 99509 103989
rect 99537 103961 99571 103989
rect 99599 103961 102485 103989
rect 102513 103961 102547 103989
rect 102575 103961 102609 103989
rect 102637 103961 102671 103989
rect 102699 103961 104009 103989
rect 104037 103961 104071 103989
rect 104099 103961 108509 103989
rect 108537 103961 108571 103989
rect 108599 103961 111485 103989
rect 111513 103961 111547 103989
rect 111575 103961 111609 103989
rect 111637 103961 111671 103989
rect 111699 103961 113009 103989
rect 113037 103961 113071 103989
rect 113099 103961 117509 103989
rect 117537 103961 117571 103989
rect 117599 103961 120485 103989
rect 120513 103961 120547 103989
rect 120575 103961 120609 103989
rect 120637 103961 120671 103989
rect 120699 103961 129485 103989
rect 129513 103961 129547 103989
rect 129575 103961 129609 103989
rect 129637 103961 129671 103989
rect 129699 103961 138485 103989
rect 138513 103961 138547 103989
rect 138575 103961 138609 103989
rect 138637 103961 138671 103989
rect 138699 103961 147485 103989
rect 147513 103961 147547 103989
rect 147575 103961 147609 103989
rect 147637 103961 147671 103989
rect 147699 103961 156485 103989
rect 156513 103961 156547 103989
rect 156575 103961 156609 103989
rect 156637 103961 156671 103989
rect 156699 103961 165485 103989
rect 165513 103961 165547 103989
rect 165575 103961 165609 103989
rect 165637 103961 165671 103989
rect 165699 103961 174485 103989
rect 174513 103961 174547 103989
rect 174575 103961 174609 103989
rect 174637 103961 174671 103989
rect 174699 103961 183485 103989
rect 183513 103961 183547 103989
rect 183575 103961 183609 103989
rect 183637 103961 183671 103989
rect 183699 103961 192485 103989
rect 192513 103961 192547 103989
rect 192575 103961 192609 103989
rect 192637 103961 192671 103989
rect 192699 103961 201485 103989
rect 201513 103961 201547 103989
rect 201575 103961 201609 103989
rect 201637 103961 201671 103989
rect 201699 103961 210485 103989
rect 210513 103961 210547 103989
rect 210575 103961 210609 103989
rect 210637 103961 210671 103989
rect 210699 103961 219485 103989
rect 219513 103961 219547 103989
rect 219575 103961 219609 103989
rect 219637 103961 219671 103989
rect 219699 103961 228485 103989
rect 228513 103961 228547 103989
rect 228575 103961 228609 103989
rect 228637 103961 228671 103989
rect 228699 103961 237485 103989
rect 237513 103961 237547 103989
rect 237575 103961 237609 103989
rect 237637 103961 237671 103989
rect 237699 103961 246485 103989
rect 246513 103961 246547 103989
rect 246575 103961 246609 103989
rect 246637 103961 246671 103989
rect 246699 103961 255485 103989
rect 255513 103961 255547 103989
rect 255575 103961 255609 103989
rect 255637 103961 255671 103989
rect 255699 103961 264485 103989
rect 264513 103961 264547 103989
rect 264575 103961 264609 103989
rect 264637 103961 264671 103989
rect 264699 103961 273485 103989
rect 273513 103961 273547 103989
rect 273575 103961 273609 103989
rect 273637 103961 273671 103989
rect 273699 103961 282485 103989
rect 282513 103961 282547 103989
rect 282575 103961 282609 103989
rect 282637 103961 282671 103989
rect 282699 103961 291485 103989
rect 291513 103961 291547 103989
rect 291575 103961 291609 103989
rect 291637 103961 291671 103989
rect 291699 103961 298728 103989
rect 298756 103961 298790 103989
rect 298818 103961 298852 103989
rect 298880 103961 298914 103989
rect 298942 103961 298990 103989
rect -958 103913 298990 103961
rect -958 101175 298990 101223
rect -958 101147 -430 101175
rect -402 101147 -368 101175
rect -340 101147 -306 101175
rect -278 101147 -244 101175
rect -216 101147 1625 101175
rect 1653 101147 1687 101175
rect 1715 101147 1749 101175
rect 1777 101147 1811 101175
rect 1839 101147 10625 101175
rect 10653 101147 10687 101175
rect 10715 101147 10749 101175
rect 10777 101147 10811 101175
rect 10839 101147 19625 101175
rect 19653 101147 19687 101175
rect 19715 101147 19749 101175
rect 19777 101147 19811 101175
rect 19839 101147 28625 101175
rect 28653 101147 28687 101175
rect 28715 101147 28749 101175
rect 28777 101147 28811 101175
rect 28839 101147 37625 101175
rect 37653 101147 37687 101175
rect 37715 101147 37749 101175
rect 37777 101147 37811 101175
rect 37839 101147 46625 101175
rect 46653 101147 46687 101175
rect 46715 101147 46749 101175
rect 46777 101147 46811 101175
rect 46839 101147 52259 101175
rect 52287 101147 52321 101175
rect 52349 101147 55625 101175
rect 55653 101147 55687 101175
rect 55715 101147 55749 101175
rect 55777 101147 55811 101175
rect 55839 101147 56759 101175
rect 56787 101147 56821 101175
rect 56849 101147 61259 101175
rect 61287 101147 61321 101175
rect 61349 101147 64625 101175
rect 64653 101147 64687 101175
rect 64715 101147 64749 101175
rect 64777 101147 64811 101175
rect 64839 101147 65759 101175
rect 65787 101147 65821 101175
rect 65849 101147 70259 101175
rect 70287 101147 70321 101175
rect 70349 101147 73625 101175
rect 73653 101147 73687 101175
rect 73715 101147 73749 101175
rect 73777 101147 73811 101175
rect 73839 101147 74759 101175
rect 74787 101147 74821 101175
rect 74849 101147 79259 101175
rect 79287 101147 79321 101175
rect 79349 101147 82625 101175
rect 82653 101147 82687 101175
rect 82715 101147 82749 101175
rect 82777 101147 82811 101175
rect 82839 101147 83759 101175
rect 83787 101147 83821 101175
rect 83849 101147 88259 101175
rect 88287 101147 88321 101175
rect 88349 101147 91625 101175
rect 91653 101147 91687 101175
rect 91715 101147 91749 101175
rect 91777 101147 91811 101175
rect 91839 101147 92759 101175
rect 92787 101147 92821 101175
rect 92849 101147 97259 101175
rect 97287 101147 97321 101175
rect 97349 101147 100625 101175
rect 100653 101147 100687 101175
rect 100715 101147 100749 101175
rect 100777 101147 100811 101175
rect 100839 101147 101759 101175
rect 101787 101147 101821 101175
rect 101849 101147 106259 101175
rect 106287 101147 106321 101175
rect 106349 101147 109625 101175
rect 109653 101147 109687 101175
rect 109715 101147 109749 101175
rect 109777 101147 109811 101175
rect 109839 101147 110759 101175
rect 110787 101147 110821 101175
rect 110849 101147 115259 101175
rect 115287 101147 115321 101175
rect 115349 101147 118625 101175
rect 118653 101147 118687 101175
rect 118715 101147 118749 101175
rect 118777 101147 118811 101175
rect 118839 101147 127625 101175
rect 127653 101147 127687 101175
rect 127715 101147 127749 101175
rect 127777 101147 127811 101175
rect 127839 101147 136625 101175
rect 136653 101147 136687 101175
rect 136715 101147 136749 101175
rect 136777 101147 136811 101175
rect 136839 101147 145625 101175
rect 145653 101147 145687 101175
rect 145715 101147 145749 101175
rect 145777 101147 145811 101175
rect 145839 101147 154625 101175
rect 154653 101147 154687 101175
rect 154715 101147 154749 101175
rect 154777 101147 154811 101175
rect 154839 101147 163625 101175
rect 163653 101147 163687 101175
rect 163715 101147 163749 101175
rect 163777 101147 163811 101175
rect 163839 101147 172625 101175
rect 172653 101147 172687 101175
rect 172715 101147 172749 101175
rect 172777 101147 172811 101175
rect 172839 101147 181625 101175
rect 181653 101147 181687 101175
rect 181715 101147 181749 101175
rect 181777 101147 181811 101175
rect 181839 101147 190625 101175
rect 190653 101147 190687 101175
rect 190715 101147 190749 101175
rect 190777 101147 190811 101175
rect 190839 101147 199625 101175
rect 199653 101147 199687 101175
rect 199715 101147 199749 101175
rect 199777 101147 199811 101175
rect 199839 101147 208625 101175
rect 208653 101147 208687 101175
rect 208715 101147 208749 101175
rect 208777 101147 208811 101175
rect 208839 101147 217625 101175
rect 217653 101147 217687 101175
rect 217715 101147 217749 101175
rect 217777 101147 217811 101175
rect 217839 101147 226625 101175
rect 226653 101147 226687 101175
rect 226715 101147 226749 101175
rect 226777 101147 226811 101175
rect 226839 101147 235625 101175
rect 235653 101147 235687 101175
rect 235715 101147 235749 101175
rect 235777 101147 235811 101175
rect 235839 101147 244625 101175
rect 244653 101147 244687 101175
rect 244715 101147 244749 101175
rect 244777 101147 244811 101175
rect 244839 101147 253625 101175
rect 253653 101147 253687 101175
rect 253715 101147 253749 101175
rect 253777 101147 253811 101175
rect 253839 101147 262625 101175
rect 262653 101147 262687 101175
rect 262715 101147 262749 101175
rect 262777 101147 262811 101175
rect 262839 101147 271625 101175
rect 271653 101147 271687 101175
rect 271715 101147 271749 101175
rect 271777 101147 271811 101175
rect 271839 101147 280625 101175
rect 280653 101147 280687 101175
rect 280715 101147 280749 101175
rect 280777 101147 280811 101175
rect 280839 101147 289625 101175
rect 289653 101147 289687 101175
rect 289715 101147 289749 101175
rect 289777 101147 289811 101175
rect 289839 101147 298248 101175
rect 298276 101147 298310 101175
rect 298338 101147 298372 101175
rect 298400 101147 298434 101175
rect 298462 101147 298990 101175
rect -958 101113 298990 101147
rect -958 101085 -430 101113
rect -402 101085 -368 101113
rect -340 101085 -306 101113
rect -278 101085 -244 101113
rect -216 101085 1625 101113
rect 1653 101085 1687 101113
rect 1715 101085 1749 101113
rect 1777 101085 1811 101113
rect 1839 101085 10625 101113
rect 10653 101085 10687 101113
rect 10715 101085 10749 101113
rect 10777 101085 10811 101113
rect 10839 101085 19625 101113
rect 19653 101085 19687 101113
rect 19715 101085 19749 101113
rect 19777 101085 19811 101113
rect 19839 101085 28625 101113
rect 28653 101085 28687 101113
rect 28715 101085 28749 101113
rect 28777 101085 28811 101113
rect 28839 101085 37625 101113
rect 37653 101085 37687 101113
rect 37715 101085 37749 101113
rect 37777 101085 37811 101113
rect 37839 101085 46625 101113
rect 46653 101085 46687 101113
rect 46715 101085 46749 101113
rect 46777 101085 46811 101113
rect 46839 101085 52259 101113
rect 52287 101085 52321 101113
rect 52349 101085 55625 101113
rect 55653 101085 55687 101113
rect 55715 101085 55749 101113
rect 55777 101085 55811 101113
rect 55839 101085 56759 101113
rect 56787 101085 56821 101113
rect 56849 101085 61259 101113
rect 61287 101085 61321 101113
rect 61349 101085 64625 101113
rect 64653 101085 64687 101113
rect 64715 101085 64749 101113
rect 64777 101085 64811 101113
rect 64839 101085 65759 101113
rect 65787 101085 65821 101113
rect 65849 101085 70259 101113
rect 70287 101085 70321 101113
rect 70349 101085 73625 101113
rect 73653 101085 73687 101113
rect 73715 101085 73749 101113
rect 73777 101085 73811 101113
rect 73839 101085 74759 101113
rect 74787 101085 74821 101113
rect 74849 101085 79259 101113
rect 79287 101085 79321 101113
rect 79349 101085 82625 101113
rect 82653 101085 82687 101113
rect 82715 101085 82749 101113
rect 82777 101085 82811 101113
rect 82839 101085 83759 101113
rect 83787 101085 83821 101113
rect 83849 101085 88259 101113
rect 88287 101085 88321 101113
rect 88349 101085 91625 101113
rect 91653 101085 91687 101113
rect 91715 101085 91749 101113
rect 91777 101085 91811 101113
rect 91839 101085 92759 101113
rect 92787 101085 92821 101113
rect 92849 101085 97259 101113
rect 97287 101085 97321 101113
rect 97349 101085 100625 101113
rect 100653 101085 100687 101113
rect 100715 101085 100749 101113
rect 100777 101085 100811 101113
rect 100839 101085 101759 101113
rect 101787 101085 101821 101113
rect 101849 101085 106259 101113
rect 106287 101085 106321 101113
rect 106349 101085 109625 101113
rect 109653 101085 109687 101113
rect 109715 101085 109749 101113
rect 109777 101085 109811 101113
rect 109839 101085 110759 101113
rect 110787 101085 110821 101113
rect 110849 101085 115259 101113
rect 115287 101085 115321 101113
rect 115349 101085 118625 101113
rect 118653 101085 118687 101113
rect 118715 101085 118749 101113
rect 118777 101085 118811 101113
rect 118839 101085 127625 101113
rect 127653 101085 127687 101113
rect 127715 101085 127749 101113
rect 127777 101085 127811 101113
rect 127839 101085 136625 101113
rect 136653 101085 136687 101113
rect 136715 101085 136749 101113
rect 136777 101085 136811 101113
rect 136839 101085 145625 101113
rect 145653 101085 145687 101113
rect 145715 101085 145749 101113
rect 145777 101085 145811 101113
rect 145839 101085 154625 101113
rect 154653 101085 154687 101113
rect 154715 101085 154749 101113
rect 154777 101085 154811 101113
rect 154839 101085 163625 101113
rect 163653 101085 163687 101113
rect 163715 101085 163749 101113
rect 163777 101085 163811 101113
rect 163839 101085 172625 101113
rect 172653 101085 172687 101113
rect 172715 101085 172749 101113
rect 172777 101085 172811 101113
rect 172839 101085 181625 101113
rect 181653 101085 181687 101113
rect 181715 101085 181749 101113
rect 181777 101085 181811 101113
rect 181839 101085 190625 101113
rect 190653 101085 190687 101113
rect 190715 101085 190749 101113
rect 190777 101085 190811 101113
rect 190839 101085 199625 101113
rect 199653 101085 199687 101113
rect 199715 101085 199749 101113
rect 199777 101085 199811 101113
rect 199839 101085 208625 101113
rect 208653 101085 208687 101113
rect 208715 101085 208749 101113
rect 208777 101085 208811 101113
rect 208839 101085 217625 101113
rect 217653 101085 217687 101113
rect 217715 101085 217749 101113
rect 217777 101085 217811 101113
rect 217839 101085 226625 101113
rect 226653 101085 226687 101113
rect 226715 101085 226749 101113
rect 226777 101085 226811 101113
rect 226839 101085 235625 101113
rect 235653 101085 235687 101113
rect 235715 101085 235749 101113
rect 235777 101085 235811 101113
rect 235839 101085 244625 101113
rect 244653 101085 244687 101113
rect 244715 101085 244749 101113
rect 244777 101085 244811 101113
rect 244839 101085 253625 101113
rect 253653 101085 253687 101113
rect 253715 101085 253749 101113
rect 253777 101085 253811 101113
rect 253839 101085 262625 101113
rect 262653 101085 262687 101113
rect 262715 101085 262749 101113
rect 262777 101085 262811 101113
rect 262839 101085 271625 101113
rect 271653 101085 271687 101113
rect 271715 101085 271749 101113
rect 271777 101085 271811 101113
rect 271839 101085 280625 101113
rect 280653 101085 280687 101113
rect 280715 101085 280749 101113
rect 280777 101085 280811 101113
rect 280839 101085 289625 101113
rect 289653 101085 289687 101113
rect 289715 101085 289749 101113
rect 289777 101085 289811 101113
rect 289839 101085 298248 101113
rect 298276 101085 298310 101113
rect 298338 101085 298372 101113
rect 298400 101085 298434 101113
rect 298462 101085 298990 101113
rect -958 101051 298990 101085
rect -958 101023 -430 101051
rect -402 101023 -368 101051
rect -340 101023 -306 101051
rect -278 101023 -244 101051
rect -216 101023 1625 101051
rect 1653 101023 1687 101051
rect 1715 101023 1749 101051
rect 1777 101023 1811 101051
rect 1839 101023 10625 101051
rect 10653 101023 10687 101051
rect 10715 101023 10749 101051
rect 10777 101023 10811 101051
rect 10839 101023 19625 101051
rect 19653 101023 19687 101051
rect 19715 101023 19749 101051
rect 19777 101023 19811 101051
rect 19839 101023 28625 101051
rect 28653 101023 28687 101051
rect 28715 101023 28749 101051
rect 28777 101023 28811 101051
rect 28839 101023 37625 101051
rect 37653 101023 37687 101051
rect 37715 101023 37749 101051
rect 37777 101023 37811 101051
rect 37839 101023 46625 101051
rect 46653 101023 46687 101051
rect 46715 101023 46749 101051
rect 46777 101023 46811 101051
rect 46839 101023 52259 101051
rect 52287 101023 52321 101051
rect 52349 101023 55625 101051
rect 55653 101023 55687 101051
rect 55715 101023 55749 101051
rect 55777 101023 55811 101051
rect 55839 101023 56759 101051
rect 56787 101023 56821 101051
rect 56849 101023 61259 101051
rect 61287 101023 61321 101051
rect 61349 101023 64625 101051
rect 64653 101023 64687 101051
rect 64715 101023 64749 101051
rect 64777 101023 64811 101051
rect 64839 101023 65759 101051
rect 65787 101023 65821 101051
rect 65849 101023 70259 101051
rect 70287 101023 70321 101051
rect 70349 101023 73625 101051
rect 73653 101023 73687 101051
rect 73715 101023 73749 101051
rect 73777 101023 73811 101051
rect 73839 101023 74759 101051
rect 74787 101023 74821 101051
rect 74849 101023 79259 101051
rect 79287 101023 79321 101051
rect 79349 101023 82625 101051
rect 82653 101023 82687 101051
rect 82715 101023 82749 101051
rect 82777 101023 82811 101051
rect 82839 101023 83759 101051
rect 83787 101023 83821 101051
rect 83849 101023 88259 101051
rect 88287 101023 88321 101051
rect 88349 101023 91625 101051
rect 91653 101023 91687 101051
rect 91715 101023 91749 101051
rect 91777 101023 91811 101051
rect 91839 101023 92759 101051
rect 92787 101023 92821 101051
rect 92849 101023 97259 101051
rect 97287 101023 97321 101051
rect 97349 101023 100625 101051
rect 100653 101023 100687 101051
rect 100715 101023 100749 101051
rect 100777 101023 100811 101051
rect 100839 101023 101759 101051
rect 101787 101023 101821 101051
rect 101849 101023 106259 101051
rect 106287 101023 106321 101051
rect 106349 101023 109625 101051
rect 109653 101023 109687 101051
rect 109715 101023 109749 101051
rect 109777 101023 109811 101051
rect 109839 101023 110759 101051
rect 110787 101023 110821 101051
rect 110849 101023 115259 101051
rect 115287 101023 115321 101051
rect 115349 101023 118625 101051
rect 118653 101023 118687 101051
rect 118715 101023 118749 101051
rect 118777 101023 118811 101051
rect 118839 101023 127625 101051
rect 127653 101023 127687 101051
rect 127715 101023 127749 101051
rect 127777 101023 127811 101051
rect 127839 101023 136625 101051
rect 136653 101023 136687 101051
rect 136715 101023 136749 101051
rect 136777 101023 136811 101051
rect 136839 101023 145625 101051
rect 145653 101023 145687 101051
rect 145715 101023 145749 101051
rect 145777 101023 145811 101051
rect 145839 101023 154625 101051
rect 154653 101023 154687 101051
rect 154715 101023 154749 101051
rect 154777 101023 154811 101051
rect 154839 101023 163625 101051
rect 163653 101023 163687 101051
rect 163715 101023 163749 101051
rect 163777 101023 163811 101051
rect 163839 101023 172625 101051
rect 172653 101023 172687 101051
rect 172715 101023 172749 101051
rect 172777 101023 172811 101051
rect 172839 101023 181625 101051
rect 181653 101023 181687 101051
rect 181715 101023 181749 101051
rect 181777 101023 181811 101051
rect 181839 101023 190625 101051
rect 190653 101023 190687 101051
rect 190715 101023 190749 101051
rect 190777 101023 190811 101051
rect 190839 101023 199625 101051
rect 199653 101023 199687 101051
rect 199715 101023 199749 101051
rect 199777 101023 199811 101051
rect 199839 101023 208625 101051
rect 208653 101023 208687 101051
rect 208715 101023 208749 101051
rect 208777 101023 208811 101051
rect 208839 101023 217625 101051
rect 217653 101023 217687 101051
rect 217715 101023 217749 101051
rect 217777 101023 217811 101051
rect 217839 101023 226625 101051
rect 226653 101023 226687 101051
rect 226715 101023 226749 101051
rect 226777 101023 226811 101051
rect 226839 101023 235625 101051
rect 235653 101023 235687 101051
rect 235715 101023 235749 101051
rect 235777 101023 235811 101051
rect 235839 101023 244625 101051
rect 244653 101023 244687 101051
rect 244715 101023 244749 101051
rect 244777 101023 244811 101051
rect 244839 101023 253625 101051
rect 253653 101023 253687 101051
rect 253715 101023 253749 101051
rect 253777 101023 253811 101051
rect 253839 101023 262625 101051
rect 262653 101023 262687 101051
rect 262715 101023 262749 101051
rect 262777 101023 262811 101051
rect 262839 101023 271625 101051
rect 271653 101023 271687 101051
rect 271715 101023 271749 101051
rect 271777 101023 271811 101051
rect 271839 101023 280625 101051
rect 280653 101023 280687 101051
rect 280715 101023 280749 101051
rect 280777 101023 280811 101051
rect 280839 101023 289625 101051
rect 289653 101023 289687 101051
rect 289715 101023 289749 101051
rect 289777 101023 289811 101051
rect 289839 101023 298248 101051
rect 298276 101023 298310 101051
rect 298338 101023 298372 101051
rect 298400 101023 298434 101051
rect 298462 101023 298990 101051
rect -958 100989 298990 101023
rect -958 100961 -430 100989
rect -402 100961 -368 100989
rect -340 100961 -306 100989
rect -278 100961 -244 100989
rect -216 100961 1625 100989
rect 1653 100961 1687 100989
rect 1715 100961 1749 100989
rect 1777 100961 1811 100989
rect 1839 100961 10625 100989
rect 10653 100961 10687 100989
rect 10715 100961 10749 100989
rect 10777 100961 10811 100989
rect 10839 100961 19625 100989
rect 19653 100961 19687 100989
rect 19715 100961 19749 100989
rect 19777 100961 19811 100989
rect 19839 100961 28625 100989
rect 28653 100961 28687 100989
rect 28715 100961 28749 100989
rect 28777 100961 28811 100989
rect 28839 100961 37625 100989
rect 37653 100961 37687 100989
rect 37715 100961 37749 100989
rect 37777 100961 37811 100989
rect 37839 100961 46625 100989
rect 46653 100961 46687 100989
rect 46715 100961 46749 100989
rect 46777 100961 46811 100989
rect 46839 100961 52259 100989
rect 52287 100961 52321 100989
rect 52349 100961 55625 100989
rect 55653 100961 55687 100989
rect 55715 100961 55749 100989
rect 55777 100961 55811 100989
rect 55839 100961 56759 100989
rect 56787 100961 56821 100989
rect 56849 100961 61259 100989
rect 61287 100961 61321 100989
rect 61349 100961 64625 100989
rect 64653 100961 64687 100989
rect 64715 100961 64749 100989
rect 64777 100961 64811 100989
rect 64839 100961 65759 100989
rect 65787 100961 65821 100989
rect 65849 100961 70259 100989
rect 70287 100961 70321 100989
rect 70349 100961 73625 100989
rect 73653 100961 73687 100989
rect 73715 100961 73749 100989
rect 73777 100961 73811 100989
rect 73839 100961 74759 100989
rect 74787 100961 74821 100989
rect 74849 100961 79259 100989
rect 79287 100961 79321 100989
rect 79349 100961 82625 100989
rect 82653 100961 82687 100989
rect 82715 100961 82749 100989
rect 82777 100961 82811 100989
rect 82839 100961 83759 100989
rect 83787 100961 83821 100989
rect 83849 100961 88259 100989
rect 88287 100961 88321 100989
rect 88349 100961 91625 100989
rect 91653 100961 91687 100989
rect 91715 100961 91749 100989
rect 91777 100961 91811 100989
rect 91839 100961 92759 100989
rect 92787 100961 92821 100989
rect 92849 100961 97259 100989
rect 97287 100961 97321 100989
rect 97349 100961 100625 100989
rect 100653 100961 100687 100989
rect 100715 100961 100749 100989
rect 100777 100961 100811 100989
rect 100839 100961 101759 100989
rect 101787 100961 101821 100989
rect 101849 100961 106259 100989
rect 106287 100961 106321 100989
rect 106349 100961 109625 100989
rect 109653 100961 109687 100989
rect 109715 100961 109749 100989
rect 109777 100961 109811 100989
rect 109839 100961 110759 100989
rect 110787 100961 110821 100989
rect 110849 100961 115259 100989
rect 115287 100961 115321 100989
rect 115349 100961 118625 100989
rect 118653 100961 118687 100989
rect 118715 100961 118749 100989
rect 118777 100961 118811 100989
rect 118839 100961 127625 100989
rect 127653 100961 127687 100989
rect 127715 100961 127749 100989
rect 127777 100961 127811 100989
rect 127839 100961 136625 100989
rect 136653 100961 136687 100989
rect 136715 100961 136749 100989
rect 136777 100961 136811 100989
rect 136839 100961 145625 100989
rect 145653 100961 145687 100989
rect 145715 100961 145749 100989
rect 145777 100961 145811 100989
rect 145839 100961 154625 100989
rect 154653 100961 154687 100989
rect 154715 100961 154749 100989
rect 154777 100961 154811 100989
rect 154839 100961 163625 100989
rect 163653 100961 163687 100989
rect 163715 100961 163749 100989
rect 163777 100961 163811 100989
rect 163839 100961 172625 100989
rect 172653 100961 172687 100989
rect 172715 100961 172749 100989
rect 172777 100961 172811 100989
rect 172839 100961 181625 100989
rect 181653 100961 181687 100989
rect 181715 100961 181749 100989
rect 181777 100961 181811 100989
rect 181839 100961 190625 100989
rect 190653 100961 190687 100989
rect 190715 100961 190749 100989
rect 190777 100961 190811 100989
rect 190839 100961 199625 100989
rect 199653 100961 199687 100989
rect 199715 100961 199749 100989
rect 199777 100961 199811 100989
rect 199839 100961 208625 100989
rect 208653 100961 208687 100989
rect 208715 100961 208749 100989
rect 208777 100961 208811 100989
rect 208839 100961 217625 100989
rect 217653 100961 217687 100989
rect 217715 100961 217749 100989
rect 217777 100961 217811 100989
rect 217839 100961 226625 100989
rect 226653 100961 226687 100989
rect 226715 100961 226749 100989
rect 226777 100961 226811 100989
rect 226839 100961 235625 100989
rect 235653 100961 235687 100989
rect 235715 100961 235749 100989
rect 235777 100961 235811 100989
rect 235839 100961 244625 100989
rect 244653 100961 244687 100989
rect 244715 100961 244749 100989
rect 244777 100961 244811 100989
rect 244839 100961 253625 100989
rect 253653 100961 253687 100989
rect 253715 100961 253749 100989
rect 253777 100961 253811 100989
rect 253839 100961 262625 100989
rect 262653 100961 262687 100989
rect 262715 100961 262749 100989
rect 262777 100961 262811 100989
rect 262839 100961 271625 100989
rect 271653 100961 271687 100989
rect 271715 100961 271749 100989
rect 271777 100961 271811 100989
rect 271839 100961 280625 100989
rect 280653 100961 280687 100989
rect 280715 100961 280749 100989
rect 280777 100961 280811 100989
rect 280839 100961 289625 100989
rect 289653 100961 289687 100989
rect 289715 100961 289749 100989
rect 289777 100961 289811 100989
rect 289839 100961 298248 100989
rect 298276 100961 298310 100989
rect 298338 100961 298372 100989
rect 298400 100961 298434 100989
rect 298462 100961 298990 100989
rect -958 100913 298990 100961
rect -958 95175 298990 95223
rect -958 95147 -910 95175
rect -882 95147 -848 95175
rect -820 95147 -786 95175
rect -758 95147 -724 95175
rect -696 95147 3485 95175
rect 3513 95147 3547 95175
rect 3575 95147 3609 95175
rect 3637 95147 3671 95175
rect 3699 95147 12485 95175
rect 12513 95147 12547 95175
rect 12575 95147 12609 95175
rect 12637 95147 12671 95175
rect 12699 95147 21485 95175
rect 21513 95147 21547 95175
rect 21575 95147 21609 95175
rect 21637 95147 21671 95175
rect 21699 95147 30485 95175
rect 30513 95147 30547 95175
rect 30575 95147 30609 95175
rect 30637 95147 30671 95175
rect 30699 95147 39485 95175
rect 39513 95147 39547 95175
rect 39575 95147 39609 95175
rect 39637 95147 39671 95175
rect 39699 95147 48485 95175
rect 48513 95147 48547 95175
rect 48575 95147 48609 95175
rect 48637 95147 48671 95175
rect 48699 95147 54509 95175
rect 54537 95147 54571 95175
rect 54599 95147 57485 95175
rect 57513 95147 57547 95175
rect 57575 95147 57609 95175
rect 57637 95147 57671 95175
rect 57699 95147 59009 95175
rect 59037 95147 59071 95175
rect 59099 95147 63509 95175
rect 63537 95147 63571 95175
rect 63599 95147 66485 95175
rect 66513 95147 66547 95175
rect 66575 95147 66609 95175
rect 66637 95147 66671 95175
rect 66699 95147 68009 95175
rect 68037 95147 68071 95175
rect 68099 95147 72509 95175
rect 72537 95147 72571 95175
rect 72599 95147 75485 95175
rect 75513 95147 75547 95175
rect 75575 95147 75609 95175
rect 75637 95147 75671 95175
rect 75699 95147 77009 95175
rect 77037 95147 77071 95175
rect 77099 95147 81509 95175
rect 81537 95147 81571 95175
rect 81599 95147 84485 95175
rect 84513 95147 84547 95175
rect 84575 95147 84609 95175
rect 84637 95147 84671 95175
rect 84699 95147 86009 95175
rect 86037 95147 86071 95175
rect 86099 95147 90509 95175
rect 90537 95147 90571 95175
rect 90599 95147 95009 95175
rect 95037 95147 95071 95175
rect 95099 95147 99509 95175
rect 99537 95147 99571 95175
rect 99599 95147 104009 95175
rect 104037 95147 104071 95175
rect 104099 95147 108509 95175
rect 108537 95147 108571 95175
rect 108599 95147 113009 95175
rect 113037 95147 113071 95175
rect 113099 95147 117509 95175
rect 117537 95147 117571 95175
rect 117599 95147 120485 95175
rect 120513 95147 120547 95175
rect 120575 95147 120609 95175
rect 120637 95147 120671 95175
rect 120699 95147 129485 95175
rect 129513 95147 129547 95175
rect 129575 95147 129609 95175
rect 129637 95147 129671 95175
rect 129699 95147 138485 95175
rect 138513 95147 138547 95175
rect 138575 95147 138609 95175
rect 138637 95147 138671 95175
rect 138699 95147 147485 95175
rect 147513 95147 147547 95175
rect 147575 95147 147609 95175
rect 147637 95147 147671 95175
rect 147699 95147 156485 95175
rect 156513 95147 156547 95175
rect 156575 95147 156609 95175
rect 156637 95147 156671 95175
rect 156699 95147 165485 95175
rect 165513 95147 165547 95175
rect 165575 95147 165609 95175
rect 165637 95147 165671 95175
rect 165699 95147 174485 95175
rect 174513 95147 174547 95175
rect 174575 95147 174609 95175
rect 174637 95147 174671 95175
rect 174699 95147 183485 95175
rect 183513 95147 183547 95175
rect 183575 95147 183609 95175
rect 183637 95147 183671 95175
rect 183699 95147 192485 95175
rect 192513 95147 192547 95175
rect 192575 95147 192609 95175
rect 192637 95147 192671 95175
rect 192699 95147 201485 95175
rect 201513 95147 201547 95175
rect 201575 95147 201609 95175
rect 201637 95147 201671 95175
rect 201699 95147 210485 95175
rect 210513 95147 210547 95175
rect 210575 95147 210609 95175
rect 210637 95147 210671 95175
rect 210699 95147 219485 95175
rect 219513 95147 219547 95175
rect 219575 95147 219609 95175
rect 219637 95147 219671 95175
rect 219699 95147 228485 95175
rect 228513 95147 228547 95175
rect 228575 95147 228609 95175
rect 228637 95147 228671 95175
rect 228699 95147 237485 95175
rect 237513 95147 237547 95175
rect 237575 95147 237609 95175
rect 237637 95147 237671 95175
rect 237699 95147 246485 95175
rect 246513 95147 246547 95175
rect 246575 95147 246609 95175
rect 246637 95147 246671 95175
rect 246699 95147 255485 95175
rect 255513 95147 255547 95175
rect 255575 95147 255609 95175
rect 255637 95147 255671 95175
rect 255699 95147 264485 95175
rect 264513 95147 264547 95175
rect 264575 95147 264609 95175
rect 264637 95147 264671 95175
rect 264699 95147 273485 95175
rect 273513 95147 273547 95175
rect 273575 95147 273609 95175
rect 273637 95147 273671 95175
rect 273699 95147 282485 95175
rect 282513 95147 282547 95175
rect 282575 95147 282609 95175
rect 282637 95147 282671 95175
rect 282699 95147 291485 95175
rect 291513 95147 291547 95175
rect 291575 95147 291609 95175
rect 291637 95147 291671 95175
rect 291699 95147 298728 95175
rect 298756 95147 298790 95175
rect 298818 95147 298852 95175
rect 298880 95147 298914 95175
rect 298942 95147 298990 95175
rect -958 95113 298990 95147
rect -958 95085 -910 95113
rect -882 95085 -848 95113
rect -820 95085 -786 95113
rect -758 95085 -724 95113
rect -696 95085 3485 95113
rect 3513 95085 3547 95113
rect 3575 95085 3609 95113
rect 3637 95085 3671 95113
rect 3699 95085 12485 95113
rect 12513 95085 12547 95113
rect 12575 95085 12609 95113
rect 12637 95085 12671 95113
rect 12699 95085 21485 95113
rect 21513 95085 21547 95113
rect 21575 95085 21609 95113
rect 21637 95085 21671 95113
rect 21699 95085 30485 95113
rect 30513 95085 30547 95113
rect 30575 95085 30609 95113
rect 30637 95085 30671 95113
rect 30699 95085 39485 95113
rect 39513 95085 39547 95113
rect 39575 95085 39609 95113
rect 39637 95085 39671 95113
rect 39699 95085 48485 95113
rect 48513 95085 48547 95113
rect 48575 95085 48609 95113
rect 48637 95085 48671 95113
rect 48699 95085 54509 95113
rect 54537 95085 54571 95113
rect 54599 95085 57485 95113
rect 57513 95085 57547 95113
rect 57575 95085 57609 95113
rect 57637 95085 57671 95113
rect 57699 95085 59009 95113
rect 59037 95085 59071 95113
rect 59099 95085 63509 95113
rect 63537 95085 63571 95113
rect 63599 95085 66485 95113
rect 66513 95085 66547 95113
rect 66575 95085 66609 95113
rect 66637 95085 66671 95113
rect 66699 95085 68009 95113
rect 68037 95085 68071 95113
rect 68099 95085 72509 95113
rect 72537 95085 72571 95113
rect 72599 95085 75485 95113
rect 75513 95085 75547 95113
rect 75575 95085 75609 95113
rect 75637 95085 75671 95113
rect 75699 95085 77009 95113
rect 77037 95085 77071 95113
rect 77099 95085 81509 95113
rect 81537 95085 81571 95113
rect 81599 95085 84485 95113
rect 84513 95085 84547 95113
rect 84575 95085 84609 95113
rect 84637 95085 84671 95113
rect 84699 95085 86009 95113
rect 86037 95085 86071 95113
rect 86099 95085 90509 95113
rect 90537 95085 90571 95113
rect 90599 95085 95009 95113
rect 95037 95085 95071 95113
rect 95099 95085 99509 95113
rect 99537 95085 99571 95113
rect 99599 95085 104009 95113
rect 104037 95085 104071 95113
rect 104099 95085 108509 95113
rect 108537 95085 108571 95113
rect 108599 95085 113009 95113
rect 113037 95085 113071 95113
rect 113099 95085 117509 95113
rect 117537 95085 117571 95113
rect 117599 95085 120485 95113
rect 120513 95085 120547 95113
rect 120575 95085 120609 95113
rect 120637 95085 120671 95113
rect 120699 95085 129485 95113
rect 129513 95085 129547 95113
rect 129575 95085 129609 95113
rect 129637 95085 129671 95113
rect 129699 95085 138485 95113
rect 138513 95085 138547 95113
rect 138575 95085 138609 95113
rect 138637 95085 138671 95113
rect 138699 95085 147485 95113
rect 147513 95085 147547 95113
rect 147575 95085 147609 95113
rect 147637 95085 147671 95113
rect 147699 95085 156485 95113
rect 156513 95085 156547 95113
rect 156575 95085 156609 95113
rect 156637 95085 156671 95113
rect 156699 95085 165485 95113
rect 165513 95085 165547 95113
rect 165575 95085 165609 95113
rect 165637 95085 165671 95113
rect 165699 95085 174485 95113
rect 174513 95085 174547 95113
rect 174575 95085 174609 95113
rect 174637 95085 174671 95113
rect 174699 95085 183485 95113
rect 183513 95085 183547 95113
rect 183575 95085 183609 95113
rect 183637 95085 183671 95113
rect 183699 95085 192485 95113
rect 192513 95085 192547 95113
rect 192575 95085 192609 95113
rect 192637 95085 192671 95113
rect 192699 95085 201485 95113
rect 201513 95085 201547 95113
rect 201575 95085 201609 95113
rect 201637 95085 201671 95113
rect 201699 95085 210485 95113
rect 210513 95085 210547 95113
rect 210575 95085 210609 95113
rect 210637 95085 210671 95113
rect 210699 95085 219485 95113
rect 219513 95085 219547 95113
rect 219575 95085 219609 95113
rect 219637 95085 219671 95113
rect 219699 95085 228485 95113
rect 228513 95085 228547 95113
rect 228575 95085 228609 95113
rect 228637 95085 228671 95113
rect 228699 95085 237485 95113
rect 237513 95085 237547 95113
rect 237575 95085 237609 95113
rect 237637 95085 237671 95113
rect 237699 95085 246485 95113
rect 246513 95085 246547 95113
rect 246575 95085 246609 95113
rect 246637 95085 246671 95113
rect 246699 95085 255485 95113
rect 255513 95085 255547 95113
rect 255575 95085 255609 95113
rect 255637 95085 255671 95113
rect 255699 95085 264485 95113
rect 264513 95085 264547 95113
rect 264575 95085 264609 95113
rect 264637 95085 264671 95113
rect 264699 95085 273485 95113
rect 273513 95085 273547 95113
rect 273575 95085 273609 95113
rect 273637 95085 273671 95113
rect 273699 95085 282485 95113
rect 282513 95085 282547 95113
rect 282575 95085 282609 95113
rect 282637 95085 282671 95113
rect 282699 95085 291485 95113
rect 291513 95085 291547 95113
rect 291575 95085 291609 95113
rect 291637 95085 291671 95113
rect 291699 95085 298728 95113
rect 298756 95085 298790 95113
rect 298818 95085 298852 95113
rect 298880 95085 298914 95113
rect 298942 95085 298990 95113
rect -958 95051 298990 95085
rect -958 95023 -910 95051
rect -882 95023 -848 95051
rect -820 95023 -786 95051
rect -758 95023 -724 95051
rect -696 95023 3485 95051
rect 3513 95023 3547 95051
rect 3575 95023 3609 95051
rect 3637 95023 3671 95051
rect 3699 95023 12485 95051
rect 12513 95023 12547 95051
rect 12575 95023 12609 95051
rect 12637 95023 12671 95051
rect 12699 95023 21485 95051
rect 21513 95023 21547 95051
rect 21575 95023 21609 95051
rect 21637 95023 21671 95051
rect 21699 95023 30485 95051
rect 30513 95023 30547 95051
rect 30575 95023 30609 95051
rect 30637 95023 30671 95051
rect 30699 95023 39485 95051
rect 39513 95023 39547 95051
rect 39575 95023 39609 95051
rect 39637 95023 39671 95051
rect 39699 95023 48485 95051
rect 48513 95023 48547 95051
rect 48575 95023 48609 95051
rect 48637 95023 48671 95051
rect 48699 95023 54509 95051
rect 54537 95023 54571 95051
rect 54599 95023 57485 95051
rect 57513 95023 57547 95051
rect 57575 95023 57609 95051
rect 57637 95023 57671 95051
rect 57699 95023 59009 95051
rect 59037 95023 59071 95051
rect 59099 95023 63509 95051
rect 63537 95023 63571 95051
rect 63599 95023 66485 95051
rect 66513 95023 66547 95051
rect 66575 95023 66609 95051
rect 66637 95023 66671 95051
rect 66699 95023 68009 95051
rect 68037 95023 68071 95051
rect 68099 95023 72509 95051
rect 72537 95023 72571 95051
rect 72599 95023 75485 95051
rect 75513 95023 75547 95051
rect 75575 95023 75609 95051
rect 75637 95023 75671 95051
rect 75699 95023 77009 95051
rect 77037 95023 77071 95051
rect 77099 95023 81509 95051
rect 81537 95023 81571 95051
rect 81599 95023 84485 95051
rect 84513 95023 84547 95051
rect 84575 95023 84609 95051
rect 84637 95023 84671 95051
rect 84699 95023 86009 95051
rect 86037 95023 86071 95051
rect 86099 95023 90509 95051
rect 90537 95023 90571 95051
rect 90599 95023 95009 95051
rect 95037 95023 95071 95051
rect 95099 95023 99509 95051
rect 99537 95023 99571 95051
rect 99599 95023 104009 95051
rect 104037 95023 104071 95051
rect 104099 95023 108509 95051
rect 108537 95023 108571 95051
rect 108599 95023 113009 95051
rect 113037 95023 113071 95051
rect 113099 95023 117509 95051
rect 117537 95023 117571 95051
rect 117599 95023 120485 95051
rect 120513 95023 120547 95051
rect 120575 95023 120609 95051
rect 120637 95023 120671 95051
rect 120699 95023 129485 95051
rect 129513 95023 129547 95051
rect 129575 95023 129609 95051
rect 129637 95023 129671 95051
rect 129699 95023 138485 95051
rect 138513 95023 138547 95051
rect 138575 95023 138609 95051
rect 138637 95023 138671 95051
rect 138699 95023 147485 95051
rect 147513 95023 147547 95051
rect 147575 95023 147609 95051
rect 147637 95023 147671 95051
rect 147699 95023 156485 95051
rect 156513 95023 156547 95051
rect 156575 95023 156609 95051
rect 156637 95023 156671 95051
rect 156699 95023 165485 95051
rect 165513 95023 165547 95051
rect 165575 95023 165609 95051
rect 165637 95023 165671 95051
rect 165699 95023 174485 95051
rect 174513 95023 174547 95051
rect 174575 95023 174609 95051
rect 174637 95023 174671 95051
rect 174699 95023 183485 95051
rect 183513 95023 183547 95051
rect 183575 95023 183609 95051
rect 183637 95023 183671 95051
rect 183699 95023 192485 95051
rect 192513 95023 192547 95051
rect 192575 95023 192609 95051
rect 192637 95023 192671 95051
rect 192699 95023 201485 95051
rect 201513 95023 201547 95051
rect 201575 95023 201609 95051
rect 201637 95023 201671 95051
rect 201699 95023 210485 95051
rect 210513 95023 210547 95051
rect 210575 95023 210609 95051
rect 210637 95023 210671 95051
rect 210699 95023 219485 95051
rect 219513 95023 219547 95051
rect 219575 95023 219609 95051
rect 219637 95023 219671 95051
rect 219699 95023 228485 95051
rect 228513 95023 228547 95051
rect 228575 95023 228609 95051
rect 228637 95023 228671 95051
rect 228699 95023 237485 95051
rect 237513 95023 237547 95051
rect 237575 95023 237609 95051
rect 237637 95023 237671 95051
rect 237699 95023 246485 95051
rect 246513 95023 246547 95051
rect 246575 95023 246609 95051
rect 246637 95023 246671 95051
rect 246699 95023 255485 95051
rect 255513 95023 255547 95051
rect 255575 95023 255609 95051
rect 255637 95023 255671 95051
rect 255699 95023 264485 95051
rect 264513 95023 264547 95051
rect 264575 95023 264609 95051
rect 264637 95023 264671 95051
rect 264699 95023 273485 95051
rect 273513 95023 273547 95051
rect 273575 95023 273609 95051
rect 273637 95023 273671 95051
rect 273699 95023 282485 95051
rect 282513 95023 282547 95051
rect 282575 95023 282609 95051
rect 282637 95023 282671 95051
rect 282699 95023 291485 95051
rect 291513 95023 291547 95051
rect 291575 95023 291609 95051
rect 291637 95023 291671 95051
rect 291699 95023 298728 95051
rect 298756 95023 298790 95051
rect 298818 95023 298852 95051
rect 298880 95023 298914 95051
rect 298942 95023 298990 95051
rect -958 94989 298990 95023
rect -958 94961 -910 94989
rect -882 94961 -848 94989
rect -820 94961 -786 94989
rect -758 94961 -724 94989
rect -696 94961 3485 94989
rect 3513 94961 3547 94989
rect 3575 94961 3609 94989
rect 3637 94961 3671 94989
rect 3699 94961 12485 94989
rect 12513 94961 12547 94989
rect 12575 94961 12609 94989
rect 12637 94961 12671 94989
rect 12699 94961 21485 94989
rect 21513 94961 21547 94989
rect 21575 94961 21609 94989
rect 21637 94961 21671 94989
rect 21699 94961 30485 94989
rect 30513 94961 30547 94989
rect 30575 94961 30609 94989
rect 30637 94961 30671 94989
rect 30699 94961 39485 94989
rect 39513 94961 39547 94989
rect 39575 94961 39609 94989
rect 39637 94961 39671 94989
rect 39699 94961 48485 94989
rect 48513 94961 48547 94989
rect 48575 94961 48609 94989
rect 48637 94961 48671 94989
rect 48699 94961 54509 94989
rect 54537 94961 54571 94989
rect 54599 94961 57485 94989
rect 57513 94961 57547 94989
rect 57575 94961 57609 94989
rect 57637 94961 57671 94989
rect 57699 94961 59009 94989
rect 59037 94961 59071 94989
rect 59099 94961 63509 94989
rect 63537 94961 63571 94989
rect 63599 94961 66485 94989
rect 66513 94961 66547 94989
rect 66575 94961 66609 94989
rect 66637 94961 66671 94989
rect 66699 94961 68009 94989
rect 68037 94961 68071 94989
rect 68099 94961 72509 94989
rect 72537 94961 72571 94989
rect 72599 94961 75485 94989
rect 75513 94961 75547 94989
rect 75575 94961 75609 94989
rect 75637 94961 75671 94989
rect 75699 94961 77009 94989
rect 77037 94961 77071 94989
rect 77099 94961 81509 94989
rect 81537 94961 81571 94989
rect 81599 94961 84485 94989
rect 84513 94961 84547 94989
rect 84575 94961 84609 94989
rect 84637 94961 84671 94989
rect 84699 94961 86009 94989
rect 86037 94961 86071 94989
rect 86099 94961 90509 94989
rect 90537 94961 90571 94989
rect 90599 94961 95009 94989
rect 95037 94961 95071 94989
rect 95099 94961 99509 94989
rect 99537 94961 99571 94989
rect 99599 94961 104009 94989
rect 104037 94961 104071 94989
rect 104099 94961 108509 94989
rect 108537 94961 108571 94989
rect 108599 94961 113009 94989
rect 113037 94961 113071 94989
rect 113099 94961 117509 94989
rect 117537 94961 117571 94989
rect 117599 94961 120485 94989
rect 120513 94961 120547 94989
rect 120575 94961 120609 94989
rect 120637 94961 120671 94989
rect 120699 94961 129485 94989
rect 129513 94961 129547 94989
rect 129575 94961 129609 94989
rect 129637 94961 129671 94989
rect 129699 94961 138485 94989
rect 138513 94961 138547 94989
rect 138575 94961 138609 94989
rect 138637 94961 138671 94989
rect 138699 94961 147485 94989
rect 147513 94961 147547 94989
rect 147575 94961 147609 94989
rect 147637 94961 147671 94989
rect 147699 94961 156485 94989
rect 156513 94961 156547 94989
rect 156575 94961 156609 94989
rect 156637 94961 156671 94989
rect 156699 94961 165485 94989
rect 165513 94961 165547 94989
rect 165575 94961 165609 94989
rect 165637 94961 165671 94989
rect 165699 94961 174485 94989
rect 174513 94961 174547 94989
rect 174575 94961 174609 94989
rect 174637 94961 174671 94989
rect 174699 94961 183485 94989
rect 183513 94961 183547 94989
rect 183575 94961 183609 94989
rect 183637 94961 183671 94989
rect 183699 94961 192485 94989
rect 192513 94961 192547 94989
rect 192575 94961 192609 94989
rect 192637 94961 192671 94989
rect 192699 94961 201485 94989
rect 201513 94961 201547 94989
rect 201575 94961 201609 94989
rect 201637 94961 201671 94989
rect 201699 94961 210485 94989
rect 210513 94961 210547 94989
rect 210575 94961 210609 94989
rect 210637 94961 210671 94989
rect 210699 94961 219485 94989
rect 219513 94961 219547 94989
rect 219575 94961 219609 94989
rect 219637 94961 219671 94989
rect 219699 94961 228485 94989
rect 228513 94961 228547 94989
rect 228575 94961 228609 94989
rect 228637 94961 228671 94989
rect 228699 94961 237485 94989
rect 237513 94961 237547 94989
rect 237575 94961 237609 94989
rect 237637 94961 237671 94989
rect 237699 94961 246485 94989
rect 246513 94961 246547 94989
rect 246575 94961 246609 94989
rect 246637 94961 246671 94989
rect 246699 94961 255485 94989
rect 255513 94961 255547 94989
rect 255575 94961 255609 94989
rect 255637 94961 255671 94989
rect 255699 94961 264485 94989
rect 264513 94961 264547 94989
rect 264575 94961 264609 94989
rect 264637 94961 264671 94989
rect 264699 94961 273485 94989
rect 273513 94961 273547 94989
rect 273575 94961 273609 94989
rect 273637 94961 273671 94989
rect 273699 94961 282485 94989
rect 282513 94961 282547 94989
rect 282575 94961 282609 94989
rect 282637 94961 282671 94989
rect 282699 94961 291485 94989
rect 291513 94961 291547 94989
rect 291575 94961 291609 94989
rect 291637 94961 291671 94989
rect 291699 94961 298728 94989
rect 298756 94961 298790 94989
rect 298818 94961 298852 94989
rect 298880 94961 298914 94989
rect 298942 94961 298990 94989
rect -958 94913 298990 94961
rect -958 92175 298990 92223
rect -958 92147 -430 92175
rect -402 92147 -368 92175
rect -340 92147 -306 92175
rect -278 92147 -244 92175
rect -216 92147 1625 92175
rect 1653 92147 1687 92175
rect 1715 92147 1749 92175
rect 1777 92147 1811 92175
rect 1839 92147 10625 92175
rect 10653 92147 10687 92175
rect 10715 92147 10749 92175
rect 10777 92147 10811 92175
rect 10839 92147 19625 92175
rect 19653 92147 19687 92175
rect 19715 92147 19749 92175
rect 19777 92147 19811 92175
rect 19839 92147 28625 92175
rect 28653 92147 28687 92175
rect 28715 92147 28749 92175
rect 28777 92147 28811 92175
rect 28839 92147 37625 92175
rect 37653 92147 37687 92175
rect 37715 92147 37749 92175
rect 37777 92147 37811 92175
rect 37839 92147 46625 92175
rect 46653 92147 46687 92175
rect 46715 92147 46749 92175
rect 46777 92147 46811 92175
rect 46839 92147 52259 92175
rect 52287 92147 52321 92175
rect 52349 92147 55625 92175
rect 55653 92147 55687 92175
rect 55715 92147 55749 92175
rect 55777 92147 55811 92175
rect 55839 92147 56759 92175
rect 56787 92147 56821 92175
rect 56849 92147 61259 92175
rect 61287 92147 61321 92175
rect 61349 92147 64625 92175
rect 64653 92147 64687 92175
rect 64715 92147 64749 92175
rect 64777 92147 64811 92175
rect 64839 92147 65759 92175
rect 65787 92147 65821 92175
rect 65849 92147 70259 92175
rect 70287 92147 70321 92175
rect 70349 92147 73625 92175
rect 73653 92147 73687 92175
rect 73715 92147 73749 92175
rect 73777 92147 73811 92175
rect 73839 92147 74759 92175
rect 74787 92147 74821 92175
rect 74849 92147 79259 92175
rect 79287 92147 79321 92175
rect 79349 92147 82625 92175
rect 82653 92147 82687 92175
rect 82715 92147 82749 92175
rect 82777 92147 82811 92175
rect 82839 92147 83759 92175
rect 83787 92147 83821 92175
rect 83849 92147 88259 92175
rect 88287 92147 88321 92175
rect 88349 92147 91625 92175
rect 91653 92147 91687 92175
rect 91715 92147 91749 92175
rect 91777 92147 91811 92175
rect 91839 92147 92759 92175
rect 92787 92147 92821 92175
rect 92849 92147 97259 92175
rect 97287 92147 97321 92175
rect 97349 92147 101759 92175
rect 101787 92147 101821 92175
rect 101849 92147 106259 92175
rect 106287 92147 106321 92175
rect 106349 92147 110759 92175
rect 110787 92147 110821 92175
rect 110849 92147 115259 92175
rect 115287 92147 115321 92175
rect 115349 92147 127625 92175
rect 127653 92147 127687 92175
rect 127715 92147 127749 92175
rect 127777 92147 127811 92175
rect 127839 92147 136625 92175
rect 136653 92147 136687 92175
rect 136715 92147 136749 92175
rect 136777 92147 136811 92175
rect 136839 92147 145625 92175
rect 145653 92147 145687 92175
rect 145715 92147 145749 92175
rect 145777 92147 145811 92175
rect 145839 92147 154625 92175
rect 154653 92147 154687 92175
rect 154715 92147 154749 92175
rect 154777 92147 154811 92175
rect 154839 92147 163625 92175
rect 163653 92147 163687 92175
rect 163715 92147 163749 92175
rect 163777 92147 163811 92175
rect 163839 92147 172625 92175
rect 172653 92147 172687 92175
rect 172715 92147 172749 92175
rect 172777 92147 172811 92175
rect 172839 92147 181625 92175
rect 181653 92147 181687 92175
rect 181715 92147 181749 92175
rect 181777 92147 181811 92175
rect 181839 92147 190625 92175
rect 190653 92147 190687 92175
rect 190715 92147 190749 92175
rect 190777 92147 190811 92175
rect 190839 92147 199625 92175
rect 199653 92147 199687 92175
rect 199715 92147 199749 92175
rect 199777 92147 199811 92175
rect 199839 92147 208625 92175
rect 208653 92147 208687 92175
rect 208715 92147 208749 92175
rect 208777 92147 208811 92175
rect 208839 92147 217625 92175
rect 217653 92147 217687 92175
rect 217715 92147 217749 92175
rect 217777 92147 217811 92175
rect 217839 92147 226625 92175
rect 226653 92147 226687 92175
rect 226715 92147 226749 92175
rect 226777 92147 226811 92175
rect 226839 92147 235625 92175
rect 235653 92147 235687 92175
rect 235715 92147 235749 92175
rect 235777 92147 235811 92175
rect 235839 92147 244625 92175
rect 244653 92147 244687 92175
rect 244715 92147 244749 92175
rect 244777 92147 244811 92175
rect 244839 92147 253625 92175
rect 253653 92147 253687 92175
rect 253715 92147 253749 92175
rect 253777 92147 253811 92175
rect 253839 92147 262625 92175
rect 262653 92147 262687 92175
rect 262715 92147 262749 92175
rect 262777 92147 262811 92175
rect 262839 92147 271625 92175
rect 271653 92147 271687 92175
rect 271715 92147 271749 92175
rect 271777 92147 271811 92175
rect 271839 92147 280625 92175
rect 280653 92147 280687 92175
rect 280715 92147 280749 92175
rect 280777 92147 280811 92175
rect 280839 92147 289625 92175
rect 289653 92147 289687 92175
rect 289715 92147 289749 92175
rect 289777 92147 289811 92175
rect 289839 92147 298248 92175
rect 298276 92147 298310 92175
rect 298338 92147 298372 92175
rect 298400 92147 298434 92175
rect 298462 92147 298990 92175
rect -958 92113 298990 92147
rect -958 92085 -430 92113
rect -402 92085 -368 92113
rect -340 92085 -306 92113
rect -278 92085 -244 92113
rect -216 92085 1625 92113
rect 1653 92085 1687 92113
rect 1715 92085 1749 92113
rect 1777 92085 1811 92113
rect 1839 92085 10625 92113
rect 10653 92085 10687 92113
rect 10715 92085 10749 92113
rect 10777 92085 10811 92113
rect 10839 92085 19625 92113
rect 19653 92085 19687 92113
rect 19715 92085 19749 92113
rect 19777 92085 19811 92113
rect 19839 92085 28625 92113
rect 28653 92085 28687 92113
rect 28715 92085 28749 92113
rect 28777 92085 28811 92113
rect 28839 92085 37625 92113
rect 37653 92085 37687 92113
rect 37715 92085 37749 92113
rect 37777 92085 37811 92113
rect 37839 92085 46625 92113
rect 46653 92085 46687 92113
rect 46715 92085 46749 92113
rect 46777 92085 46811 92113
rect 46839 92085 52259 92113
rect 52287 92085 52321 92113
rect 52349 92085 55625 92113
rect 55653 92085 55687 92113
rect 55715 92085 55749 92113
rect 55777 92085 55811 92113
rect 55839 92085 56759 92113
rect 56787 92085 56821 92113
rect 56849 92085 61259 92113
rect 61287 92085 61321 92113
rect 61349 92085 64625 92113
rect 64653 92085 64687 92113
rect 64715 92085 64749 92113
rect 64777 92085 64811 92113
rect 64839 92085 65759 92113
rect 65787 92085 65821 92113
rect 65849 92085 70259 92113
rect 70287 92085 70321 92113
rect 70349 92085 73625 92113
rect 73653 92085 73687 92113
rect 73715 92085 73749 92113
rect 73777 92085 73811 92113
rect 73839 92085 74759 92113
rect 74787 92085 74821 92113
rect 74849 92085 79259 92113
rect 79287 92085 79321 92113
rect 79349 92085 82625 92113
rect 82653 92085 82687 92113
rect 82715 92085 82749 92113
rect 82777 92085 82811 92113
rect 82839 92085 83759 92113
rect 83787 92085 83821 92113
rect 83849 92085 88259 92113
rect 88287 92085 88321 92113
rect 88349 92085 91625 92113
rect 91653 92085 91687 92113
rect 91715 92085 91749 92113
rect 91777 92085 91811 92113
rect 91839 92085 92759 92113
rect 92787 92085 92821 92113
rect 92849 92085 97259 92113
rect 97287 92085 97321 92113
rect 97349 92085 101759 92113
rect 101787 92085 101821 92113
rect 101849 92085 106259 92113
rect 106287 92085 106321 92113
rect 106349 92085 110759 92113
rect 110787 92085 110821 92113
rect 110849 92085 115259 92113
rect 115287 92085 115321 92113
rect 115349 92085 127625 92113
rect 127653 92085 127687 92113
rect 127715 92085 127749 92113
rect 127777 92085 127811 92113
rect 127839 92085 136625 92113
rect 136653 92085 136687 92113
rect 136715 92085 136749 92113
rect 136777 92085 136811 92113
rect 136839 92085 145625 92113
rect 145653 92085 145687 92113
rect 145715 92085 145749 92113
rect 145777 92085 145811 92113
rect 145839 92085 154625 92113
rect 154653 92085 154687 92113
rect 154715 92085 154749 92113
rect 154777 92085 154811 92113
rect 154839 92085 163625 92113
rect 163653 92085 163687 92113
rect 163715 92085 163749 92113
rect 163777 92085 163811 92113
rect 163839 92085 172625 92113
rect 172653 92085 172687 92113
rect 172715 92085 172749 92113
rect 172777 92085 172811 92113
rect 172839 92085 181625 92113
rect 181653 92085 181687 92113
rect 181715 92085 181749 92113
rect 181777 92085 181811 92113
rect 181839 92085 190625 92113
rect 190653 92085 190687 92113
rect 190715 92085 190749 92113
rect 190777 92085 190811 92113
rect 190839 92085 199625 92113
rect 199653 92085 199687 92113
rect 199715 92085 199749 92113
rect 199777 92085 199811 92113
rect 199839 92085 208625 92113
rect 208653 92085 208687 92113
rect 208715 92085 208749 92113
rect 208777 92085 208811 92113
rect 208839 92085 217625 92113
rect 217653 92085 217687 92113
rect 217715 92085 217749 92113
rect 217777 92085 217811 92113
rect 217839 92085 226625 92113
rect 226653 92085 226687 92113
rect 226715 92085 226749 92113
rect 226777 92085 226811 92113
rect 226839 92085 235625 92113
rect 235653 92085 235687 92113
rect 235715 92085 235749 92113
rect 235777 92085 235811 92113
rect 235839 92085 244625 92113
rect 244653 92085 244687 92113
rect 244715 92085 244749 92113
rect 244777 92085 244811 92113
rect 244839 92085 253625 92113
rect 253653 92085 253687 92113
rect 253715 92085 253749 92113
rect 253777 92085 253811 92113
rect 253839 92085 262625 92113
rect 262653 92085 262687 92113
rect 262715 92085 262749 92113
rect 262777 92085 262811 92113
rect 262839 92085 271625 92113
rect 271653 92085 271687 92113
rect 271715 92085 271749 92113
rect 271777 92085 271811 92113
rect 271839 92085 280625 92113
rect 280653 92085 280687 92113
rect 280715 92085 280749 92113
rect 280777 92085 280811 92113
rect 280839 92085 289625 92113
rect 289653 92085 289687 92113
rect 289715 92085 289749 92113
rect 289777 92085 289811 92113
rect 289839 92085 298248 92113
rect 298276 92085 298310 92113
rect 298338 92085 298372 92113
rect 298400 92085 298434 92113
rect 298462 92085 298990 92113
rect -958 92051 298990 92085
rect -958 92023 -430 92051
rect -402 92023 -368 92051
rect -340 92023 -306 92051
rect -278 92023 -244 92051
rect -216 92023 1625 92051
rect 1653 92023 1687 92051
rect 1715 92023 1749 92051
rect 1777 92023 1811 92051
rect 1839 92023 10625 92051
rect 10653 92023 10687 92051
rect 10715 92023 10749 92051
rect 10777 92023 10811 92051
rect 10839 92023 19625 92051
rect 19653 92023 19687 92051
rect 19715 92023 19749 92051
rect 19777 92023 19811 92051
rect 19839 92023 28625 92051
rect 28653 92023 28687 92051
rect 28715 92023 28749 92051
rect 28777 92023 28811 92051
rect 28839 92023 37625 92051
rect 37653 92023 37687 92051
rect 37715 92023 37749 92051
rect 37777 92023 37811 92051
rect 37839 92023 46625 92051
rect 46653 92023 46687 92051
rect 46715 92023 46749 92051
rect 46777 92023 46811 92051
rect 46839 92023 52259 92051
rect 52287 92023 52321 92051
rect 52349 92023 55625 92051
rect 55653 92023 55687 92051
rect 55715 92023 55749 92051
rect 55777 92023 55811 92051
rect 55839 92023 56759 92051
rect 56787 92023 56821 92051
rect 56849 92023 61259 92051
rect 61287 92023 61321 92051
rect 61349 92023 64625 92051
rect 64653 92023 64687 92051
rect 64715 92023 64749 92051
rect 64777 92023 64811 92051
rect 64839 92023 65759 92051
rect 65787 92023 65821 92051
rect 65849 92023 70259 92051
rect 70287 92023 70321 92051
rect 70349 92023 73625 92051
rect 73653 92023 73687 92051
rect 73715 92023 73749 92051
rect 73777 92023 73811 92051
rect 73839 92023 74759 92051
rect 74787 92023 74821 92051
rect 74849 92023 79259 92051
rect 79287 92023 79321 92051
rect 79349 92023 82625 92051
rect 82653 92023 82687 92051
rect 82715 92023 82749 92051
rect 82777 92023 82811 92051
rect 82839 92023 83759 92051
rect 83787 92023 83821 92051
rect 83849 92023 88259 92051
rect 88287 92023 88321 92051
rect 88349 92023 91625 92051
rect 91653 92023 91687 92051
rect 91715 92023 91749 92051
rect 91777 92023 91811 92051
rect 91839 92023 92759 92051
rect 92787 92023 92821 92051
rect 92849 92023 97259 92051
rect 97287 92023 97321 92051
rect 97349 92023 101759 92051
rect 101787 92023 101821 92051
rect 101849 92023 106259 92051
rect 106287 92023 106321 92051
rect 106349 92023 110759 92051
rect 110787 92023 110821 92051
rect 110849 92023 115259 92051
rect 115287 92023 115321 92051
rect 115349 92023 127625 92051
rect 127653 92023 127687 92051
rect 127715 92023 127749 92051
rect 127777 92023 127811 92051
rect 127839 92023 136625 92051
rect 136653 92023 136687 92051
rect 136715 92023 136749 92051
rect 136777 92023 136811 92051
rect 136839 92023 145625 92051
rect 145653 92023 145687 92051
rect 145715 92023 145749 92051
rect 145777 92023 145811 92051
rect 145839 92023 154625 92051
rect 154653 92023 154687 92051
rect 154715 92023 154749 92051
rect 154777 92023 154811 92051
rect 154839 92023 163625 92051
rect 163653 92023 163687 92051
rect 163715 92023 163749 92051
rect 163777 92023 163811 92051
rect 163839 92023 172625 92051
rect 172653 92023 172687 92051
rect 172715 92023 172749 92051
rect 172777 92023 172811 92051
rect 172839 92023 181625 92051
rect 181653 92023 181687 92051
rect 181715 92023 181749 92051
rect 181777 92023 181811 92051
rect 181839 92023 190625 92051
rect 190653 92023 190687 92051
rect 190715 92023 190749 92051
rect 190777 92023 190811 92051
rect 190839 92023 199625 92051
rect 199653 92023 199687 92051
rect 199715 92023 199749 92051
rect 199777 92023 199811 92051
rect 199839 92023 208625 92051
rect 208653 92023 208687 92051
rect 208715 92023 208749 92051
rect 208777 92023 208811 92051
rect 208839 92023 217625 92051
rect 217653 92023 217687 92051
rect 217715 92023 217749 92051
rect 217777 92023 217811 92051
rect 217839 92023 226625 92051
rect 226653 92023 226687 92051
rect 226715 92023 226749 92051
rect 226777 92023 226811 92051
rect 226839 92023 235625 92051
rect 235653 92023 235687 92051
rect 235715 92023 235749 92051
rect 235777 92023 235811 92051
rect 235839 92023 244625 92051
rect 244653 92023 244687 92051
rect 244715 92023 244749 92051
rect 244777 92023 244811 92051
rect 244839 92023 253625 92051
rect 253653 92023 253687 92051
rect 253715 92023 253749 92051
rect 253777 92023 253811 92051
rect 253839 92023 262625 92051
rect 262653 92023 262687 92051
rect 262715 92023 262749 92051
rect 262777 92023 262811 92051
rect 262839 92023 271625 92051
rect 271653 92023 271687 92051
rect 271715 92023 271749 92051
rect 271777 92023 271811 92051
rect 271839 92023 280625 92051
rect 280653 92023 280687 92051
rect 280715 92023 280749 92051
rect 280777 92023 280811 92051
rect 280839 92023 289625 92051
rect 289653 92023 289687 92051
rect 289715 92023 289749 92051
rect 289777 92023 289811 92051
rect 289839 92023 298248 92051
rect 298276 92023 298310 92051
rect 298338 92023 298372 92051
rect 298400 92023 298434 92051
rect 298462 92023 298990 92051
rect -958 91989 298990 92023
rect -958 91961 -430 91989
rect -402 91961 -368 91989
rect -340 91961 -306 91989
rect -278 91961 -244 91989
rect -216 91961 1625 91989
rect 1653 91961 1687 91989
rect 1715 91961 1749 91989
rect 1777 91961 1811 91989
rect 1839 91961 10625 91989
rect 10653 91961 10687 91989
rect 10715 91961 10749 91989
rect 10777 91961 10811 91989
rect 10839 91961 19625 91989
rect 19653 91961 19687 91989
rect 19715 91961 19749 91989
rect 19777 91961 19811 91989
rect 19839 91961 28625 91989
rect 28653 91961 28687 91989
rect 28715 91961 28749 91989
rect 28777 91961 28811 91989
rect 28839 91961 37625 91989
rect 37653 91961 37687 91989
rect 37715 91961 37749 91989
rect 37777 91961 37811 91989
rect 37839 91961 46625 91989
rect 46653 91961 46687 91989
rect 46715 91961 46749 91989
rect 46777 91961 46811 91989
rect 46839 91961 52259 91989
rect 52287 91961 52321 91989
rect 52349 91961 55625 91989
rect 55653 91961 55687 91989
rect 55715 91961 55749 91989
rect 55777 91961 55811 91989
rect 55839 91961 56759 91989
rect 56787 91961 56821 91989
rect 56849 91961 61259 91989
rect 61287 91961 61321 91989
rect 61349 91961 64625 91989
rect 64653 91961 64687 91989
rect 64715 91961 64749 91989
rect 64777 91961 64811 91989
rect 64839 91961 65759 91989
rect 65787 91961 65821 91989
rect 65849 91961 70259 91989
rect 70287 91961 70321 91989
rect 70349 91961 73625 91989
rect 73653 91961 73687 91989
rect 73715 91961 73749 91989
rect 73777 91961 73811 91989
rect 73839 91961 74759 91989
rect 74787 91961 74821 91989
rect 74849 91961 79259 91989
rect 79287 91961 79321 91989
rect 79349 91961 82625 91989
rect 82653 91961 82687 91989
rect 82715 91961 82749 91989
rect 82777 91961 82811 91989
rect 82839 91961 83759 91989
rect 83787 91961 83821 91989
rect 83849 91961 88259 91989
rect 88287 91961 88321 91989
rect 88349 91961 91625 91989
rect 91653 91961 91687 91989
rect 91715 91961 91749 91989
rect 91777 91961 91811 91989
rect 91839 91961 92759 91989
rect 92787 91961 92821 91989
rect 92849 91961 97259 91989
rect 97287 91961 97321 91989
rect 97349 91961 101759 91989
rect 101787 91961 101821 91989
rect 101849 91961 106259 91989
rect 106287 91961 106321 91989
rect 106349 91961 110759 91989
rect 110787 91961 110821 91989
rect 110849 91961 115259 91989
rect 115287 91961 115321 91989
rect 115349 91961 127625 91989
rect 127653 91961 127687 91989
rect 127715 91961 127749 91989
rect 127777 91961 127811 91989
rect 127839 91961 136625 91989
rect 136653 91961 136687 91989
rect 136715 91961 136749 91989
rect 136777 91961 136811 91989
rect 136839 91961 145625 91989
rect 145653 91961 145687 91989
rect 145715 91961 145749 91989
rect 145777 91961 145811 91989
rect 145839 91961 154625 91989
rect 154653 91961 154687 91989
rect 154715 91961 154749 91989
rect 154777 91961 154811 91989
rect 154839 91961 163625 91989
rect 163653 91961 163687 91989
rect 163715 91961 163749 91989
rect 163777 91961 163811 91989
rect 163839 91961 172625 91989
rect 172653 91961 172687 91989
rect 172715 91961 172749 91989
rect 172777 91961 172811 91989
rect 172839 91961 181625 91989
rect 181653 91961 181687 91989
rect 181715 91961 181749 91989
rect 181777 91961 181811 91989
rect 181839 91961 190625 91989
rect 190653 91961 190687 91989
rect 190715 91961 190749 91989
rect 190777 91961 190811 91989
rect 190839 91961 199625 91989
rect 199653 91961 199687 91989
rect 199715 91961 199749 91989
rect 199777 91961 199811 91989
rect 199839 91961 208625 91989
rect 208653 91961 208687 91989
rect 208715 91961 208749 91989
rect 208777 91961 208811 91989
rect 208839 91961 217625 91989
rect 217653 91961 217687 91989
rect 217715 91961 217749 91989
rect 217777 91961 217811 91989
rect 217839 91961 226625 91989
rect 226653 91961 226687 91989
rect 226715 91961 226749 91989
rect 226777 91961 226811 91989
rect 226839 91961 235625 91989
rect 235653 91961 235687 91989
rect 235715 91961 235749 91989
rect 235777 91961 235811 91989
rect 235839 91961 244625 91989
rect 244653 91961 244687 91989
rect 244715 91961 244749 91989
rect 244777 91961 244811 91989
rect 244839 91961 253625 91989
rect 253653 91961 253687 91989
rect 253715 91961 253749 91989
rect 253777 91961 253811 91989
rect 253839 91961 262625 91989
rect 262653 91961 262687 91989
rect 262715 91961 262749 91989
rect 262777 91961 262811 91989
rect 262839 91961 271625 91989
rect 271653 91961 271687 91989
rect 271715 91961 271749 91989
rect 271777 91961 271811 91989
rect 271839 91961 280625 91989
rect 280653 91961 280687 91989
rect 280715 91961 280749 91989
rect 280777 91961 280811 91989
rect 280839 91961 289625 91989
rect 289653 91961 289687 91989
rect 289715 91961 289749 91989
rect 289777 91961 289811 91989
rect 289839 91961 298248 91989
rect 298276 91961 298310 91989
rect 298338 91961 298372 91989
rect 298400 91961 298434 91989
rect 298462 91961 298990 91989
rect -958 91913 298990 91961
rect -958 86175 298990 86223
rect -958 86147 -910 86175
rect -882 86147 -848 86175
rect -820 86147 -786 86175
rect -758 86147 -724 86175
rect -696 86147 3485 86175
rect 3513 86147 3547 86175
rect 3575 86147 3609 86175
rect 3637 86147 3671 86175
rect 3699 86147 12485 86175
rect 12513 86147 12547 86175
rect 12575 86147 12609 86175
rect 12637 86147 12671 86175
rect 12699 86147 21485 86175
rect 21513 86147 21547 86175
rect 21575 86147 21609 86175
rect 21637 86147 21671 86175
rect 21699 86147 30485 86175
rect 30513 86147 30547 86175
rect 30575 86147 30609 86175
rect 30637 86147 30671 86175
rect 30699 86147 39485 86175
rect 39513 86147 39547 86175
rect 39575 86147 39609 86175
rect 39637 86147 39671 86175
rect 39699 86147 48485 86175
rect 48513 86147 48547 86175
rect 48575 86147 48609 86175
rect 48637 86147 48671 86175
rect 48699 86147 54509 86175
rect 54537 86147 54571 86175
rect 54599 86147 57485 86175
rect 57513 86147 57547 86175
rect 57575 86147 57609 86175
rect 57637 86147 57671 86175
rect 57699 86147 59009 86175
rect 59037 86147 59071 86175
rect 59099 86147 63509 86175
rect 63537 86147 63571 86175
rect 63599 86147 66485 86175
rect 66513 86147 66547 86175
rect 66575 86147 66609 86175
rect 66637 86147 66671 86175
rect 66699 86147 68009 86175
rect 68037 86147 68071 86175
rect 68099 86147 72509 86175
rect 72537 86147 72571 86175
rect 72599 86147 75485 86175
rect 75513 86147 75547 86175
rect 75575 86147 75609 86175
rect 75637 86147 75671 86175
rect 75699 86147 77009 86175
rect 77037 86147 77071 86175
rect 77099 86147 81509 86175
rect 81537 86147 81571 86175
rect 81599 86147 84485 86175
rect 84513 86147 84547 86175
rect 84575 86147 84609 86175
rect 84637 86147 84671 86175
rect 84699 86147 86009 86175
rect 86037 86147 86071 86175
rect 86099 86147 90509 86175
rect 90537 86147 90571 86175
rect 90599 86147 95009 86175
rect 95037 86147 95071 86175
rect 95099 86147 99509 86175
rect 99537 86147 99571 86175
rect 99599 86147 104009 86175
rect 104037 86147 104071 86175
rect 104099 86147 108509 86175
rect 108537 86147 108571 86175
rect 108599 86147 113009 86175
rect 113037 86147 113071 86175
rect 113099 86147 117509 86175
rect 117537 86147 117571 86175
rect 117599 86147 120485 86175
rect 120513 86147 120547 86175
rect 120575 86147 120609 86175
rect 120637 86147 120671 86175
rect 120699 86147 129485 86175
rect 129513 86147 129547 86175
rect 129575 86147 129609 86175
rect 129637 86147 129671 86175
rect 129699 86147 138485 86175
rect 138513 86147 138547 86175
rect 138575 86147 138609 86175
rect 138637 86147 138671 86175
rect 138699 86147 147485 86175
rect 147513 86147 147547 86175
rect 147575 86147 147609 86175
rect 147637 86147 147671 86175
rect 147699 86147 156485 86175
rect 156513 86147 156547 86175
rect 156575 86147 156609 86175
rect 156637 86147 156671 86175
rect 156699 86147 165485 86175
rect 165513 86147 165547 86175
rect 165575 86147 165609 86175
rect 165637 86147 165671 86175
rect 165699 86147 174485 86175
rect 174513 86147 174547 86175
rect 174575 86147 174609 86175
rect 174637 86147 174671 86175
rect 174699 86147 183485 86175
rect 183513 86147 183547 86175
rect 183575 86147 183609 86175
rect 183637 86147 183671 86175
rect 183699 86147 192485 86175
rect 192513 86147 192547 86175
rect 192575 86147 192609 86175
rect 192637 86147 192671 86175
rect 192699 86147 201485 86175
rect 201513 86147 201547 86175
rect 201575 86147 201609 86175
rect 201637 86147 201671 86175
rect 201699 86147 210485 86175
rect 210513 86147 210547 86175
rect 210575 86147 210609 86175
rect 210637 86147 210671 86175
rect 210699 86147 219485 86175
rect 219513 86147 219547 86175
rect 219575 86147 219609 86175
rect 219637 86147 219671 86175
rect 219699 86147 228485 86175
rect 228513 86147 228547 86175
rect 228575 86147 228609 86175
rect 228637 86147 228671 86175
rect 228699 86147 237485 86175
rect 237513 86147 237547 86175
rect 237575 86147 237609 86175
rect 237637 86147 237671 86175
rect 237699 86147 246485 86175
rect 246513 86147 246547 86175
rect 246575 86147 246609 86175
rect 246637 86147 246671 86175
rect 246699 86147 255485 86175
rect 255513 86147 255547 86175
rect 255575 86147 255609 86175
rect 255637 86147 255671 86175
rect 255699 86147 264485 86175
rect 264513 86147 264547 86175
rect 264575 86147 264609 86175
rect 264637 86147 264671 86175
rect 264699 86147 273485 86175
rect 273513 86147 273547 86175
rect 273575 86147 273609 86175
rect 273637 86147 273671 86175
rect 273699 86147 282485 86175
rect 282513 86147 282547 86175
rect 282575 86147 282609 86175
rect 282637 86147 282671 86175
rect 282699 86147 291485 86175
rect 291513 86147 291547 86175
rect 291575 86147 291609 86175
rect 291637 86147 291671 86175
rect 291699 86147 298728 86175
rect 298756 86147 298790 86175
rect 298818 86147 298852 86175
rect 298880 86147 298914 86175
rect 298942 86147 298990 86175
rect -958 86113 298990 86147
rect -958 86085 -910 86113
rect -882 86085 -848 86113
rect -820 86085 -786 86113
rect -758 86085 -724 86113
rect -696 86085 3485 86113
rect 3513 86085 3547 86113
rect 3575 86085 3609 86113
rect 3637 86085 3671 86113
rect 3699 86085 12485 86113
rect 12513 86085 12547 86113
rect 12575 86085 12609 86113
rect 12637 86085 12671 86113
rect 12699 86085 21485 86113
rect 21513 86085 21547 86113
rect 21575 86085 21609 86113
rect 21637 86085 21671 86113
rect 21699 86085 30485 86113
rect 30513 86085 30547 86113
rect 30575 86085 30609 86113
rect 30637 86085 30671 86113
rect 30699 86085 39485 86113
rect 39513 86085 39547 86113
rect 39575 86085 39609 86113
rect 39637 86085 39671 86113
rect 39699 86085 48485 86113
rect 48513 86085 48547 86113
rect 48575 86085 48609 86113
rect 48637 86085 48671 86113
rect 48699 86085 54509 86113
rect 54537 86085 54571 86113
rect 54599 86085 57485 86113
rect 57513 86085 57547 86113
rect 57575 86085 57609 86113
rect 57637 86085 57671 86113
rect 57699 86085 59009 86113
rect 59037 86085 59071 86113
rect 59099 86085 63509 86113
rect 63537 86085 63571 86113
rect 63599 86085 66485 86113
rect 66513 86085 66547 86113
rect 66575 86085 66609 86113
rect 66637 86085 66671 86113
rect 66699 86085 68009 86113
rect 68037 86085 68071 86113
rect 68099 86085 72509 86113
rect 72537 86085 72571 86113
rect 72599 86085 75485 86113
rect 75513 86085 75547 86113
rect 75575 86085 75609 86113
rect 75637 86085 75671 86113
rect 75699 86085 77009 86113
rect 77037 86085 77071 86113
rect 77099 86085 81509 86113
rect 81537 86085 81571 86113
rect 81599 86085 84485 86113
rect 84513 86085 84547 86113
rect 84575 86085 84609 86113
rect 84637 86085 84671 86113
rect 84699 86085 86009 86113
rect 86037 86085 86071 86113
rect 86099 86085 90509 86113
rect 90537 86085 90571 86113
rect 90599 86085 95009 86113
rect 95037 86085 95071 86113
rect 95099 86085 99509 86113
rect 99537 86085 99571 86113
rect 99599 86085 104009 86113
rect 104037 86085 104071 86113
rect 104099 86085 108509 86113
rect 108537 86085 108571 86113
rect 108599 86085 113009 86113
rect 113037 86085 113071 86113
rect 113099 86085 117509 86113
rect 117537 86085 117571 86113
rect 117599 86085 120485 86113
rect 120513 86085 120547 86113
rect 120575 86085 120609 86113
rect 120637 86085 120671 86113
rect 120699 86085 129485 86113
rect 129513 86085 129547 86113
rect 129575 86085 129609 86113
rect 129637 86085 129671 86113
rect 129699 86085 138485 86113
rect 138513 86085 138547 86113
rect 138575 86085 138609 86113
rect 138637 86085 138671 86113
rect 138699 86085 147485 86113
rect 147513 86085 147547 86113
rect 147575 86085 147609 86113
rect 147637 86085 147671 86113
rect 147699 86085 156485 86113
rect 156513 86085 156547 86113
rect 156575 86085 156609 86113
rect 156637 86085 156671 86113
rect 156699 86085 165485 86113
rect 165513 86085 165547 86113
rect 165575 86085 165609 86113
rect 165637 86085 165671 86113
rect 165699 86085 174485 86113
rect 174513 86085 174547 86113
rect 174575 86085 174609 86113
rect 174637 86085 174671 86113
rect 174699 86085 183485 86113
rect 183513 86085 183547 86113
rect 183575 86085 183609 86113
rect 183637 86085 183671 86113
rect 183699 86085 192485 86113
rect 192513 86085 192547 86113
rect 192575 86085 192609 86113
rect 192637 86085 192671 86113
rect 192699 86085 201485 86113
rect 201513 86085 201547 86113
rect 201575 86085 201609 86113
rect 201637 86085 201671 86113
rect 201699 86085 210485 86113
rect 210513 86085 210547 86113
rect 210575 86085 210609 86113
rect 210637 86085 210671 86113
rect 210699 86085 219485 86113
rect 219513 86085 219547 86113
rect 219575 86085 219609 86113
rect 219637 86085 219671 86113
rect 219699 86085 228485 86113
rect 228513 86085 228547 86113
rect 228575 86085 228609 86113
rect 228637 86085 228671 86113
rect 228699 86085 237485 86113
rect 237513 86085 237547 86113
rect 237575 86085 237609 86113
rect 237637 86085 237671 86113
rect 237699 86085 246485 86113
rect 246513 86085 246547 86113
rect 246575 86085 246609 86113
rect 246637 86085 246671 86113
rect 246699 86085 255485 86113
rect 255513 86085 255547 86113
rect 255575 86085 255609 86113
rect 255637 86085 255671 86113
rect 255699 86085 264485 86113
rect 264513 86085 264547 86113
rect 264575 86085 264609 86113
rect 264637 86085 264671 86113
rect 264699 86085 273485 86113
rect 273513 86085 273547 86113
rect 273575 86085 273609 86113
rect 273637 86085 273671 86113
rect 273699 86085 282485 86113
rect 282513 86085 282547 86113
rect 282575 86085 282609 86113
rect 282637 86085 282671 86113
rect 282699 86085 291485 86113
rect 291513 86085 291547 86113
rect 291575 86085 291609 86113
rect 291637 86085 291671 86113
rect 291699 86085 298728 86113
rect 298756 86085 298790 86113
rect 298818 86085 298852 86113
rect 298880 86085 298914 86113
rect 298942 86085 298990 86113
rect -958 86051 298990 86085
rect -958 86023 -910 86051
rect -882 86023 -848 86051
rect -820 86023 -786 86051
rect -758 86023 -724 86051
rect -696 86023 3485 86051
rect 3513 86023 3547 86051
rect 3575 86023 3609 86051
rect 3637 86023 3671 86051
rect 3699 86023 12485 86051
rect 12513 86023 12547 86051
rect 12575 86023 12609 86051
rect 12637 86023 12671 86051
rect 12699 86023 21485 86051
rect 21513 86023 21547 86051
rect 21575 86023 21609 86051
rect 21637 86023 21671 86051
rect 21699 86023 30485 86051
rect 30513 86023 30547 86051
rect 30575 86023 30609 86051
rect 30637 86023 30671 86051
rect 30699 86023 39485 86051
rect 39513 86023 39547 86051
rect 39575 86023 39609 86051
rect 39637 86023 39671 86051
rect 39699 86023 48485 86051
rect 48513 86023 48547 86051
rect 48575 86023 48609 86051
rect 48637 86023 48671 86051
rect 48699 86023 54509 86051
rect 54537 86023 54571 86051
rect 54599 86023 57485 86051
rect 57513 86023 57547 86051
rect 57575 86023 57609 86051
rect 57637 86023 57671 86051
rect 57699 86023 59009 86051
rect 59037 86023 59071 86051
rect 59099 86023 63509 86051
rect 63537 86023 63571 86051
rect 63599 86023 66485 86051
rect 66513 86023 66547 86051
rect 66575 86023 66609 86051
rect 66637 86023 66671 86051
rect 66699 86023 68009 86051
rect 68037 86023 68071 86051
rect 68099 86023 72509 86051
rect 72537 86023 72571 86051
rect 72599 86023 75485 86051
rect 75513 86023 75547 86051
rect 75575 86023 75609 86051
rect 75637 86023 75671 86051
rect 75699 86023 77009 86051
rect 77037 86023 77071 86051
rect 77099 86023 81509 86051
rect 81537 86023 81571 86051
rect 81599 86023 84485 86051
rect 84513 86023 84547 86051
rect 84575 86023 84609 86051
rect 84637 86023 84671 86051
rect 84699 86023 86009 86051
rect 86037 86023 86071 86051
rect 86099 86023 90509 86051
rect 90537 86023 90571 86051
rect 90599 86023 95009 86051
rect 95037 86023 95071 86051
rect 95099 86023 99509 86051
rect 99537 86023 99571 86051
rect 99599 86023 104009 86051
rect 104037 86023 104071 86051
rect 104099 86023 108509 86051
rect 108537 86023 108571 86051
rect 108599 86023 113009 86051
rect 113037 86023 113071 86051
rect 113099 86023 117509 86051
rect 117537 86023 117571 86051
rect 117599 86023 120485 86051
rect 120513 86023 120547 86051
rect 120575 86023 120609 86051
rect 120637 86023 120671 86051
rect 120699 86023 129485 86051
rect 129513 86023 129547 86051
rect 129575 86023 129609 86051
rect 129637 86023 129671 86051
rect 129699 86023 138485 86051
rect 138513 86023 138547 86051
rect 138575 86023 138609 86051
rect 138637 86023 138671 86051
rect 138699 86023 147485 86051
rect 147513 86023 147547 86051
rect 147575 86023 147609 86051
rect 147637 86023 147671 86051
rect 147699 86023 156485 86051
rect 156513 86023 156547 86051
rect 156575 86023 156609 86051
rect 156637 86023 156671 86051
rect 156699 86023 165485 86051
rect 165513 86023 165547 86051
rect 165575 86023 165609 86051
rect 165637 86023 165671 86051
rect 165699 86023 174485 86051
rect 174513 86023 174547 86051
rect 174575 86023 174609 86051
rect 174637 86023 174671 86051
rect 174699 86023 183485 86051
rect 183513 86023 183547 86051
rect 183575 86023 183609 86051
rect 183637 86023 183671 86051
rect 183699 86023 192485 86051
rect 192513 86023 192547 86051
rect 192575 86023 192609 86051
rect 192637 86023 192671 86051
rect 192699 86023 201485 86051
rect 201513 86023 201547 86051
rect 201575 86023 201609 86051
rect 201637 86023 201671 86051
rect 201699 86023 210485 86051
rect 210513 86023 210547 86051
rect 210575 86023 210609 86051
rect 210637 86023 210671 86051
rect 210699 86023 219485 86051
rect 219513 86023 219547 86051
rect 219575 86023 219609 86051
rect 219637 86023 219671 86051
rect 219699 86023 228485 86051
rect 228513 86023 228547 86051
rect 228575 86023 228609 86051
rect 228637 86023 228671 86051
rect 228699 86023 237485 86051
rect 237513 86023 237547 86051
rect 237575 86023 237609 86051
rect 237637 86023 237671 86051
rect 237699 86023 246485 86051
rect 246513 86023 246547 86051
rect 246575 86023 246609 86051
rect 246637 86023 246671 86051
rect 246699 86023 255485 86051
rect 255513 86023 255547 86051
rect 255575 86023 255609 86051
rect 255637 86023 255671 86051
rect 255699 86023 264485 86051
rect 264513 86023 264547 86051
rect 264575 86023 264609 86051
rect 264637 86023 264671 86051
rect 264699 86023 273485 86051
rect 273513 86023 273547 86051
rect 273575 86023 273609 86051
rect 273637 86023 273671 86051
rect 273699 86023 282485 86051
rect 282513 86023 282547 86051
rect 282575 86023 282609 86051
rect 282637 86023 282671 86051
rect 282699 86023 291485 86051
rect 291513 86023 291547 86051
rect 291575 86023 291609 86051
rect 291637 86023 291671 86051
rect 291699 86023 298728 86051
rect 298756 86023 298790 86051
rect 298818 86023 298852 86051
rect 298880 86023 298914 86051
rect 298942 86023 298990 86051
rect -958 85989 298990 86023
rect -958 85961 -910 85989
rect -882 85961 -848 85989
rect -820 85961 -786 85989
rect -758 85961 -724 85989
rect -696 85961 3485 85989
rect 3513 85961 3547 85989
rect 3575 85961 3609 85989
rect 3637 85961 3671 85989
rect 3699 85961 12485 85989
rect 12513 85961 12547 85989
rect 12575 85961 12609 85989
rect 12637 85961 12671 85989
rect 12699 85961 21485 85989
rect 21513 85961 21547 85989
rect 21575 85961 21609 85989
rect 21637 85961 21671 85989
rect 21699 85961 30485 85989
rect 30513 85961 30547 85989
rect 30575 85961 30609 85989
rect 30637 85961 30671 85989
rect 30699 85961 39485 85989
rect 39513 85961 39547 85989
rect 39575 85961 39609 85989
rect 39637 85961 39671 85989
rect 39699 85961 48485 85989
rect 48513 85961 48547 85989
rect 48575 85961 48609 85989
rect 48637 85961 48671 85989
rect 48699 85961 54509 85989
rect 54537 85961 54571 85989
rect 54599 85961 57485 85989
rect 57513 85961 57547 85989
rect 57575 85961 57609 85989
rect 57637 85961 57671 85989
rect 57699 85961 59009 85989
rect 59037 85961 59071 85989
rect 59099 85961 63509 85989
rect 63537 85961 63571 85989
rect 63599 85961 66485 85989
rect 66513 85961 66547 85989
rect 66575 85961 66609 85989
rect 66637 85961 66671 85989
rect 66699 85961 68009 85989
rect 68037 85961 68071 85989
rect 68099 85961 72509 85989
rect 72537 85961 72571 85989
rect 72599 85961 75485 85989
rect 75513 85961 75547 85989
rect 75575 85961 75609 85989
rect 75637 85961 75671 85989
rect 75699 85961 77009 85989
rect 77037 85961 77071 85989
rect 77099 85961 81509 85989
rect 81537 85961 81571 85989
rect 81599 85961 84485 85989
rect 84513 85961 84547 85989
rect 84575 85961 84609 85989
rect 84637 85961 84671 85989
rect 84699 85961 86009 85989
rect 86037 85961 86071 85989
rect 86099 85961 90509 85989
rect 90537 85961 90571 85989
rect 90599 85961 95009 85989
rect 95037 85961 95071 85989
rect 95099 85961 99509 85989
rect 99537 85961 99571 85989
rect 99599 85961 104009 85989
rect 104037 85961 104071 85989
rect 104099 85961 108509 85989
rect 108537 85961 108571 85989
rect 108599 85961 113009 85989
rect 113037 85961 113071 85989
rect 113099 85961 117509 85989
rect 117537 85961 117571 85989
rect 117599 85961 120485 85989
rect 120513 85961 120547 85989
rect 120575 85961 120609 85989
rect 120637 85961 120671 85989
rect 120699 85961 129485 85989
rect 129513 85961 129547 85989
rect 129575 85961 129609 85989
rect 129637 85961 129671 85989
rect 129699 85961 138485 85989
rect 138513 85961 138547 85989
rect 138575 85961 138609 85989
rect 138637 85961 138671 85989
rect 138699 85961 147485 85989
rect 147513 85961 147547 85989
rect 147575 85961 147609 85989
rect 147637 85961 147671 85989
rect 147699 85961 156485 85989
rect 156513 85961 156547 85989
rect 156575 85961 156609 85989
rect 156637 85961 156671 85989
rect 156699 85961 165485 85989
rect 165513 85961 165547 85989
rect 165575 85961 165609 85989
rect 165637 85961 165671 85989
rect 165699 85961 174485 85989
rect 174513 85961 174547 85989
rect 174575 85961 174609 85989
rect 174637 85961 174671 85989
rect 174699 85961 183485 85989
rect 183513 85961 183547 85989
rect 183575 85961 183609 85989
rect 183637 85961 183671 85989
rect 183699 85961 192485 85989
rect 192513 85961 192547 85989
rect 192575 85961 192609 85989
rect 192637 85961 192671 85989
rect 192699 85961 201485 85989
rect 201513 85961 201547 85989
rect 201575 85961 201609 85989
rect 201637 85961 201671 85989
rect 201699 85961 210485 85989
rect 210513 85961 210547 85989
rect 210575 85961 210609 85989
rect 210637 85961 210671 85989
rect 210699 85961 219485 85989
rect 219513 85961 219547 85989
rect 219575 85961 219609 85989
rect 219637 85961 219671 85989
rect 219699 85961 228485 85989
rect 228513 85961 228547 85989
rect 228575 85961 228609 85989
rect 228637 85961 228671 85989
rect 228699 85961 237485 85989
rect 237513 85961 237547 85989
rect 237575 85961 237609 85989
rect 237637 85961 237671 85989
rect 237699 85961 246485 85989
rect 246513 85961 246547 85989
rect 246575 85961 246609 85989
rect 246637 85961 246671 85989
rect 246699 85961 255485 85989
rect 255513 85961 255547 85989
rect 255575 85961 255609 85989
rect 255637 85961 255671 85989
rect 255699 85961 264485 85989
rect 264513 85961 264547 85989
rect 264575 85961 264609 85989
rect 264637 85961 264671 85989
rect 264699 85961 273485 85989
rect 273513 85961 273547 85989
rect 273575 85961 273609 85989
rect 273637 85961 273671 85989
rect 273699 85961 282485 85989
rect 282513 85961 282547 85989
rect 282575 85961 282609 85989
rect 282637 85961 282671 85989
rect 282699 85961 291485 85989
rect 291513 85961 291547 85989
rect 291575 85961 291609 85989
rect 291637 85961 291671 85989
rect 291699 85961 298728 85989
rect 298756 85961 298790 85989
rect 298818 85961 298852 85989
rect 298880 85961 298914 85989
rect 298942 85961 298990 85989
rect -958 85913 298990 85961
rect -958 83175 298990 83223
rect -958 83147 -430 83175
rect -402 83147 -368 83175
rect -340 83147 -306 83175
rect -278 83147 -244 83175
rect -216 83147 1625 83175
rect 1653 83147 1687 83175
rect 1715 83147 1749 83175
rect 1777 83147 1811 83175
rect 1839 83147 10625 83175
rect 10653 83147 10687 83175
rect 10715 83147 10749 83175
rect 10777 83147 10811 83175
rect 10839 83147 19625 83175
rect 19653 83147 19687 83175
rect 19715 83147 19749 83175
rect 19777 83147 19811 83175
rect 19839 83147 28625 83175
rect 28653 83147 28687 83175
rect 28715 83147 28749 83175
rect 28777 83147 28811 83175
rect 28839 83147 37625 83175
rect 37653 83147 37687 83175
rect 37715 83147 37749 83175
rect 37777 83147 37811 83175
rect 37839 83147 46625 83175
rect 46653 83147 46687 83175
rect 46715 83147 46749 83175
rect 46777 83147 46811 83175
rect 46839 83147 52259 83175
rect 52287 83147 52321 83175
rect 52349 83147 55625 83175
rect 55653 83147 55687 83175
rect 55715 83147 55749 83175
rect 55777 83147 55811 83175
rect 55839 83147 56759 83175
rect 56787 83147 56821 83175
rect 56849 83147 61259 83175
rect 61287 83147 61321 83175
rect 61349 83147 64625 83175
rect 64653 83147 64687 83175
rect 64715 83147 64749 83175
rect 64777 83147 64811 83175
rect 64839 83147 65759 83175
rect 65787 83147 65821 83175
rect 65849 83147 70259 83175
rect 70287 83147 70321 83175
rect 70349 83147 73625 83175
rect 73653 83147 73687 83175
rect 73715 83147 73749 83175
rect 73777 83147 73811 83175
rect 73839 83147 74759 83175
rect 74787 83147 74821 83175
rect 74849 83147 79259 83175
rect 79287 83147 79321 83175
rect 79349 83147 82625 83175
rect 82653 83147 82687 83175
rect 82715 83147 82749 83175
rect 82777 83147 82811 83175
rect 82839 83147 83759 83175
rect 83787 83147 83821 83175
rect 83849 83147 88259 83175
rect 88287 83147 88321 83175
rect 88349 83147 91625 83175
rect 91653 83147 91687 83175
rect 91715 83147 91749 83175
rect 91777 83147 91811 83175
rect 91839 83147 92759 83175
rect 92787 83147 92821 83175
rect 92849 83147 97259 83175
rect 97287 83147 97321 83175
rect 97349 83147 101759 83175
rect 101787 83147 101821 83175
rect 101849 83147 106259 83175
rect 106287 83147 106321 83175
rect 106349 83147 110759 83175
rect 110787 83147 110821 83175
rect 110849 83147 115259 83175
rect 115287 83147 115321 83175
rect 115349 83147 127625 83175
rect 127653 83147 127687 83175
rect 127715 83147 127749 83175
rect 127777 83147 127811 83175
rect 127839 83147 136625 83175
rect 136653 83147 136687 83175
rect 136715 83147 136749 83175
rect 136777 83147 136811 83175
rect 136839 83147 145625 83175
rect 145653 83147 145687 83175
rect 145715 83147 145749 83175
rect 145777 83147 145811 83175
rect 145839 83147 154625 83175
rect 154653 83147 154687 83175
rect 154715 83147 154749 83175
rect 154777 83147 154811 83175
rect 154839 83147 163625 83175
rect 163653 83147 163687 83175
rect 163715 83147 163749 83175
rect 163777 83147 163811 83175
rect 163839 83147 172625 83175
rect 172653 83147 172687 83175
rect 172715 83147 172749 83175
rect 172777 83147 172811 83175
rect 172839 83147 181625 83175
rect 181653 83147 181687 83175
rect 181715 83147 181749 83175
rect 181777 83147 181811 83175
rect 181839 83147 190625 83175
rect 190653 83147 190687 83175
rect 190715 83147 190749 83175
rect 190777 83147 190811 83175
rect 190839 83147 199625 83175
rect 199653 83147 199687 83175
rect 199715 83147 199749 83175
rect 199777 83147 199811 83175
rect 199839 83147 208625 83175
rect 208653 83147 208687 83175
rect 208715 83147 208749 83175
rect 208777 83147 208811 83175
rect 208839 83147 217625 83175
rect 217653 83147 217687 83175
rect 217715 83147 217749 83175
rect 217777 83147 217811 83175
rect 217839 83147 226625 83175
rect 226653 83147 226687 83175
rect 226715 83147 226749 83175
rect 226777 83147 226811 83175
rect 226839 83147 235625 83175
rect 235653 83147 235687 83175
rect 235715 83147 235749 83175
rect 235777 83147 235811 83175
rect 235839 83147 244625 83175
rect 244653 83147 244687 83175
rect 244715 83147 244749 83175
rect 244777 83147 244811 83175
rect 244839 83147 253625 83175
rect 253653 83147 253687 83175
rect 253715 83147 253749 83175
rect 253777 83147 253811 83175
rect 253839 83147 262625 83175
rect 262653 83147 262687 83175
rect 262715 83147 262749 83175
rect 262777 83147 262811 83175
rect 262839 83147 271625 83175
rect 271653 83147 271687 83175
rect 271715 83147 271749 83175
rect 271777 83147 271811 83175
rect 271839 83147 280625 83175
rect 280653 83147 280687 83175
rect 280715 83147 280749 83175
rect 280777 83147 280811 83175
rect 280839 83147 289625 83175
rect 289653 83147 289687 83175
rect 289715 83147 289749 83175
rect 289777 83147 289811 83175
rect 289839 83147 298248 83175
rect 298276 83147 298310 83175
rect 298338 83147 298372 83175
rect 298400 83147 298434 83175
rect 298462 83147 298990 83175
rect -958 83113 298990 83147
rect -958 83085 -430 83113
rect -402 83085 -368 83113
rect -340 83085 -306 83113
rect -278 83085 -244 83113
rect -216 83085 1625 83113
rect 1653 83085 1687 83113
rect 1715 83085 1749 83113
rect 1777 83085 1811 83113
rect 1839 83085 10625 83113
rect 10653 83085 10687 83113
rect 10715 83085 10749 83113
rect 10777 83085 10811 83113
rect 10839 83085 19625 83113
rect 19653 83085 19687 83113
rect 19715 83085 19749 83113
rect 19777 83085 19811 83113
rect 19839 83085 28625 83113
rect 28653 83085 28687 83113
rect 28715 83085 28749 83113
rect 28777 83085 28811 83113
rect 28839 83085 37625 83113
rect 37653 83085 37687 83113
rect 37715 83085 37749 83113
rect 37777 83085 37811 83113
rect 37839 83085 46625 83113
rect 46653 83085 46687 83113
rect 46715 83085 46749 83113
rect 46777 83085 46811 83113
rect 46839 83085 52259 83113
rect 52287 83085 52321 83113
rect 52349 83085 55625 83113
rect 55653 83085 55687 83113
rect 55715 83085 55749 83113
rect 55777 83085 55811 83113
rect 55839 83085 56759 83113
rect 56787 83085 56821 83113
rect 56849 83085 61259 83113
rect 61287 83085 61321 83113
rect 61349 83085 64625 83113
rect 64653 83085 64687 83113
rect 64715 83085 64749 83113
rect 64777 83085 64811 83113
rect 64839 83085 65759 83113
rect 65787 83085 65821 83113
rect 65849 83085 70259 83113
rect 70287 83085 70321 83113
rect 70349 83085 73625 83113
rect 73653 83085 73687 83113
rect 73715 83085 73749 83113
rect 73777 83085 73811 83113
rect 73839 83085 74759 83113
rect 74787 83085 74821 83113
rect 74849 83085 79259 83113
rect 79287 83085 79321 83113
rect 79349 83085 82625 83113
rect 82653 83085 82687 83113
rect 82715 83085 82749 83113
rect 82777 83085 82811 83113
rect 82839 83085 83759 83113
rect 83787 83085 83821 83113
rect 83849 83085 88259 83113
rect 88287 83085 88321 83113
rect 88349 83085 91625 83113
rect 91653 83085 91687 83113
rect 91715 83085 91749 83113
rect 91777 83085 91811 83113
rect 91839 83085 92759 83113
rect 92787 83085 92821 83113
rect 92849 83085 97259 83113
rect 97287 83085 97321 83113
rect 97349 83085 101759 83113
rect 101787 83085 101821 83113
rect 101849 83085 106259 83113
rect 106287 83085 106321 83113
rect 106349 83085 110759 83113
rect 110787 83085 110821 83113
rect 110849 83085 115259 83113
rect 115287 83085 115321 83113
rect 115349 83085 127625 83113
rect 127653 83085 127687 83113
rect 127715 83085 127749 83113
rect 127777 83085 127811 83113
rect 127839 83085 136625 83113
rect 136653 83085 136687 83113
rect 136715 83085 136749 83113
rect 136777 83085 136811 83113
rect 136839 83085 145625 83113
rect 145653 83085 145687 83113
rect 145715 83085 145749 83113
rect 145777 83085 145811 83113
rect 145839 83085 154625 83113
rect 154653 83085 154687 83113
rect 154715 83085 154749 83113
rect 154777 83085 154811 83113
rect 154839 83085 163625 83113
rect 163653 83085 163687 83113
rect 163715 83085 163749 83113
rect 163777 83085 163811 83113
rect 163839 83085 172625 83113
rect 172653 83085 172687 83113
rect 172715 83085 172749 83113
rect 172777 83085 172811 83113
rect 172839 83085 181625 83113
rect 181653 83085 181687 83113
rect 181715 83085 181749 83113
rect 181777 83085 181811 83113
rect 181839 83085 190625 83113
rect 190653 83085 190687 83113
rect 190715 83085 190749 83113
rect 190777 83085 190811 83113
rect 190839 83085 199625 83113
rect 199653 83085 199687 83113
rect 199715 83085 199749 83113
rect 199777 83085 199811 83113
rect 199839 83085 208625 83113
rect 208653 83085 208687 83113
rect 208715 83085 208749 83113
rect 208777 83085 208811 83113
rect 208839 83085 217625 83113
rect 217653 83085 217687 83113
rect 217715 83085 217749 83113
rect 217777 83085 217811 83113
rect 217839 83085 226625 83113
rect 226653 83085 226687 83113
rect 226715 83085 226749 83113
rect 226777 83085 226811 83113
rect 226839 83085 235625 83113
rect 235653 83085 235687 83113
rect 235715 83085 235749 83113
rect 235777 83085 235811 83113
rect 235839 83085 244625 83113
rect 244653 83085 244687 83113
rect 244715 83085 244749 83113
rect 244777 83085 244811 83113
rect 244839 83085 253625 83113
rect 253653 83085 253687 83113
rect 253715 83085 253749 83113
rect 253777 83085 253811 83113
rect 253839 83085 262625 83113
rect 262653 83085 262687 83113
rect 262715 83085 262749 83113
rect 262777 83085 262811 83113
rect 262839 83085 271625 83113
rect 271653 83085 271687 83113
rect 271715 83085 271749 83113
rect 271777 83085 271811 83113
rect 271839 83085 280625 83113
rect 280653 83085 280687 83113
rect 280715 83085 280749 83113
rect 280777 83085 280811 83113
rect 280839 83085 289625 83113
rect 289653 83085 289687 83113
rect 289715 83085 289749 83113
rect 289777 83085 289811 83113
rect 289839 83085 298248 83113
rect 298276 83085 298310 83113
rect 298338 83085 298372 83113
rect 298400 83085 298434 83113
rect 298462 83085 298990 83113
rect -958 83051 298990 83085
rect -958 83023 -430 83051
rect -402 83023 -368 83051
rect -340 83023 -306 83051
rect -278 83023 -244 83051
rect -216 83023 1625 83051
rect 1653 83023 1687 83051
rect 1715 83023 1749 83051
rect 1777 83023 1811 83051
rect 1839 83023 10625 83051
rect 10653 83023 10687 83051
rect 10715 83023 10749 83051
rect 10777 83023 10811 83051
rect 10839 83023 19625 83051
rect 19653 83023 19687 83051
rect 19715 83023 19749 83051
rect 19777 83023 19811 83051
rect 19839 83023 28625 83051
rect 28653 83023 28687 83051
rect 28715 83023 28749 83051
rect 28777 83023 28811 83051
rect 28839 83023 37625 83051
rect 37653 83023 37687 83051
rect 37715 83023 37749 83051
rect 37777 83023 37811 83051
rect 37839 83023 46625 83051
rect 46653 83023 46687 83051
rect 46715 83023 46749 83051
rect 46777 83023 46811 83051
rect 46839 83023 52259 83051
rect 52287 83023 52321 83051
rect 52349 83023 55625 83051
rect 55653 83023 55687 83051
rect 55715 83023 55749 83051
rect 55777 83023 55811 83051
rect 55839 83023 56759 83051
rect 56787 83023 56821 83051
rect 56849 83023 61259 83051
rect 61287 83023 61321 83051
rect 61349 83023 64625 83051
rect 64653 83023 64687 83051
rect 64715 83023 64749 83051
rect 64777 83023 64811 83051
rect 64839 83023 65759 83051
rect 65787 83023 65821 83051
rect 65849 83023 70259 83051
rect 70287 83023 70321 83051
rect 70349 83023 73625 83051
rect 73653 83023 73687 83051
rect 73715 83023 73749 83051
rect 73777 83023 73811 83051
rect 73839 83023 74759 83051
rect 74787 83023 74821 83051
rect 74849 83023 79259 83051
rect 79287 83023 79321 83051
rect 79349 83023 82625 83051
rect 82653 83023 82687 83051
rect 82715 83023 82749 83051
rect 82777 83023 82811 83051
rect 82839 83023 83759 83051
rect 83787 83023 83821 83051
rect 83849 83023 88259 83051
rect 88287 83023 88321 83051
rect 88349 83023 91625 83051
rect 91653 83023 91687 83051
rect 91715 83023 91749 83051
rect 91777 83023 91811 83051
rect 91839 83023 92759 83051
rect 92787 83023 92821 83051
rect 92849 83023 97259 83051
rect 97287 83023 97321 83051
rect 97349 83023 101759 83051
rect 101787 83023 101821 83051
rect 101849 83023 106259 83051
rect 106287 83023 106321 83051
rect 106349 83023 110759 83051
rect 110787 83023 110821 83051
rect 110849 83023 115259 83051
rect 115287 83023 115321 83051
rect 115349 83023 127625 83051
rect 127653 83023 127687 83051
rect 127715 83023 127749 83051
rect 127777 83023 127811 83051
rect 127839 83023 136625 83051
rect 136653 83023 136687 83051
rect 136715 83023 136749 83051
rect 136777 83023 136811 83051
rect 136839 83023 145625 83051
rect 145653 83023 145687 83051
rect 145715 83023 145749 83051
rect 145777 83023 145811 83051
rect 145839 83023 154625 83051
rect 154653 83023 154687 83051
rect 154715 83023 154749 83051
rect 154777 83023 154811 83051
rect 154839 83023 163625 83051
rect 163653 83023 163687 83051
rect 163715 83023 163749 83051
rect 163777 83023 163811 83051
rect 163839 83023 172625 83051
rect 172653 83023 172687 83051
rect 172715 83023 172749 83051
rect 172777 83023 172811 83051
rect 172839 83023 181625 83051
rect 181653 83023 181687 83051
rect 181715 83023 181749 83051
rect 181777 83023 181811 83051
rect 181839 83023 190625 83051
rect 190653 83023 190687 83051
rect 190715 83023 190749 83051
rect 190777 83023 190811 83051
rect 190839 83023 199625 83051
rect 199653 83023 199687 83051
rect 199715 83023 199749 83051
rect 199777 83023 199811 83051
rect 199839 83023 208625 83051
rect 208653 83023 208687 83051
rect 208715 83023 208749 83051
rect 208777 83023 208811 83051
rect 208839 83023 217625 83051
rect 217653 83023 217687 83051
rect 217715 83023 217749 83051
rect 217777 83023 217811 83051
rect 217839 83023 226625 83051
rect 226653 83023 226687 83051
rect 226715 83023 226749 83051
rect 226777 83023 226811 83051
rect 226839 83023 235625 83051
rect 235653 83023 235687 83051
rect 235715 83023 235749 83051
rect 235777 83023 235811 83051
rect 235839 83023 244625 83051
rect 244653 83023 244687 83051
rect 244715 83023 244749 83051
rect 244777 83023 244811 83051
rect 244839 83023 253625 83051
rect 253653 83023 253687 83051
rect 253715 83023 253749 83051
rect 253777 83023 253811 83051
rect 253839 83023 262625 83051
rect 262653 83023 262687 83051
rect 262715 83023 262749 83051
rect 262777 83023 262811 83051
rect 262839 83023 271625 83051
rect 271653 83023 271687 83051
rect 271715 83023 271749 83051
rect 271777 83023 271811 83051
rect 271839 83023 280625 83051
rect 280653 83023 280687 83051
rect 280715 83023 280749 83051
rect 280777 83023 280811 83051
rect 280839 83023 289625 83051
rect 289653 83023 289687 83051
rect 289715 83023 289749 83051
rect 289777 83023 289811 83051
rect 289839 83023 298248 83051
rect 298276 83023 298310 83051
rect 298338 83023 298372 83051
rect 298400 83023 298434 83051
rect 298462 83023 298990 83051
rect -958 82989 298990 83023
rect -958 82961 -430 82989
rect -402 82961 -368 82989
rect -340 82961 -306 82989
rect -278 82961 -244 82989
rect -216 82961 1625 82989
rect 1653 82961 1687 82989
rect 1715 82961 1749 82989
rect 1777 82961 1811 82989
rect 1839 82961 10625 82989
rect 10653 82961 10687 82989
rect 10715 82961 10749 82989
rect 10777 82961 10811 82989
rect 10839 82961 19625 82989
rect 19653 82961 19687 82989
rect 19715 82961 19749 82989
rect 19777 82961 19811 82989
rect 19839 82961 28625 82989
rect 28653 82961 28687 82989
rect 28715 82961 28749 82989
rect 28777 82961 28811 82989
rect 28839 82961 37625 82989
rect 37653 82961 37687 82989
rect 37715 82961 37749 82989
rect 37777 82961 37811 82989
rect 37839 82961 46625 82989
rect 46653 82961 46687 82989
rect 46715 82961 46749 82989
rect 46777 82961 46811 82989
rect 46839 82961 52259 82989
rect 52287 82961 52321 82989
rect 52349 82961 55625 82989
rect 55653 82961 55687 82989
rect 55715 82961 55749 82989
rect 55777 82961 55811 82989
rect 55839 82961 56759 82989
rect 56787 82961 56821 82989
rect 56849 82961 61259 82989
rect 61287 82961 61321 82989
rect 61349 82961 64625 82989
rect 64653 82961 64687 82989
rect 64715 82961 64749 82989
rect 64777 82961 64811 82989
rect 64839 82961 65759 82989
rect 65787 82961 65821 82989
rect 65849 82961 70259 82989
rect 70287 82961 70321 82989
rect 70349 82961 73625 82989
rect 73653 82961 73687 82989
rect 73715 82961 73749 82989
rect 73777 82961 73811 82989
rect 73839 82961 74759 82989
rect 74787 82961 74821 82989
rect 74849 82961 79259 82989
rect 79287 82961 79321 82989
rect 79349 82961 82625 82989
rect 82653 82961 82687 82989
rect 82715 82961 82749 82989
rect 82777 82961 82811 82989
rect 82839 82961 83759 82989
rect 83787 82961 83821 82989
rect 83849 82961 88259 82989
rect 88287 82961 88321 82989
rect 88349 82961 91625 82989
rect 91653 82961 91687 82989
rect 91715 82961 91749 82989
rect 91777 82961 91811 82989
rect 91839 82961 92759 82989
rect 92787 82961 92821 82989
rect 92849 82961 97259 82989
rect 97287 82961 97321 82989
rect 97349 82961 101759 82989
rect 101787 82961 101821 82989
rect 101849 82961 106259 82989
rect 106287 82961 106321 82989
rect 106349 82961 110759 82989
rect 110787 82961 110821 82989
rect 110849 82961 115259 82989
rect 115287 82961 115321 82989
rect 115349 82961 127625 82989
rect 127653 82961 127687 82989
rect 127715 82961 127749 82989
rect 127777 82961 127811 82989
rect 127839 82961 136625 82989
rect 136653 82961 136687 82989
rect 136715 82961 136749 82989
rect 136777 82961 136811 82989
rect 136839 82961 145625 82989
rect 145653 82961 145687 82989
rect 145715 82961 145749 82989
rect 145777 82961 145811 82989
rect 145839 82961 154625 82989
rect 154653 82961 154687 82989
rect 154715 82961 154749 82989
rect 154777 82961 154811 82989
rect 154839 82961 163625 82989
rect 163653 82961 163687 82989
rect 163715 82961 163749 82989
rect 163777 82961 163811 82989
rect 163839 82961 172625 82989
rect 172653 82961 172687 82989
rect 172715 82961 172749 82989
rect 172777 82961 172811 82989
rect 172839 82961 181625 82989
rect 181653 82961 181687 82989
rect 181715 82961 181749 82989
rect 181777 82961 181811 82989
rect 181839 82961 190625 82989
rect 190653 82961 190687 82989
rect 190715 82961 190749 82989
rect 190777 82961 190811 82989
rect 190839 82961 199625 82989
rect 199653 82961 199687 82989
rect 199715 82961 199749 82989
rect 199777 82961 199811 82989
rect 199839 82961 208625 82989
rect 208653 82961 208687 82989
rect 208715 82961 208749 82989
rect 208777 82961 208811 82989
rect 208839 82961 217625 82989
rect 217653 82961 217687 82989
rect 217715 82961 217749 82989
rect 217777 82961 217811 82989
rect 217839 82961 226625 82989
rect 226653 82961 226687 82989
rect 226715 82961 226749 82989
rect 226777 82961 226811 82989
rect 226839 82961 235625 82989
rect 235653 82961 235687 82989
rect 235715 82961 235749 82989
rect 235777 82961 235811 82989
rect 235839 82961 244625 82989
rect 244653 82961 244687 82989
rect 244715 82961 244749 82989
rect 244777 82961 244811 82989
rect 244839 82961 253625 82989
rect 253653 82961 253687 82989
rect 253715 82961 253749 82989
rect 253777 82961 253811 82989
rect 253839 82961 262625 82989
rect 262653 82961 262687 82989
rect 262715 82961 262749 82989
rect 262777 82961 262811 82989
rect 262839 82961 271625 82989
rect 271653 82961 271687 82989
rect 271715 82961 271749 82989
rect 271777 82961 271811 82989
rect 271839 82961 280625 82989
rect 280653 82961 280687 82989
rect 280715 82961 280749 82989
rect 280777 82961 280811 82989
rect 280839 82961 289625 82989
rect 289653 82961 289687 82989
rect 289715 82961 289749 82989
rect 289777 82961 289811 82989
rect 289839 82961 298248 82989
rect 298276 82961 298310 82989
rect 298338 82961 298372 82989
rect 298400 82961 298434 82989
rect 298462 82961 298990 82989
rect -958 82913 298990 82961
rect -958 77175 298990 77223
rect -958 77147 -910 77175
rect -882 77147 -848 77175
rect -820 77147 -786 77175
rect -758 77147 -724 77175
rect -696 77147 3485 77175
rect 3513 77147 3547 77175
rect 3575 77147 3609 77175
rect 3637 77147 3671 77175
rect 3699 77147 12485 77175
rect 12513 77147 12547 77175
rect 12575 77147 12609 77175
rect 12637 77147 12671 77175
rect 12699 77147 21485 77175
rect 21513 77147 21547 77175
rect 21575 77147 21609 77175
rect 21637 77147 21671 77175
rect 21699 77147 30485 77175
rect 30513 77147 30547 77175
rect 30575 77147 30609 77175
rect 30637 77147 30671 77175
rect 30699 77147 39485 77175
rect 39513 77147 39547 77175
rect 39575 77147 39609 77175
rect 39637 77147 39671 77175
rect 39699 77147 48485 77175
rect 48513 77147 48547 77175
rect 48575 77147 48609 77175
rect 48637 77147 48671 77175
rect 48699 77147 54509 77175
rect 54537 77147 54571 77175
rect 54599 77147 57485 77175
rect 57513 77147 57547 77175
rect 57575 77147 57609 77175
rect 57637 77147 57671 77175
rect 57699 77147 59009 77175
rect 59037 77147 59071 77175
rect 59099 77147 63509 77175
rect 63537 77147 63571 77175
rect 63599 77147 66485 77175
rect 66513 77147 66547 77175
rect 66575 77147 66609 77175
rect 66637 77147 66671 77175
rect 66699 77147 68009 77175
rect 68037 77147 68071 77175
rect 68099 77147 72509 77175
rect 72537 77147 72571 77175
rect 72599 77147 75485 77175
rect 75513 77147 75547 77175
rect 75575 77147 75609 77175
rect 75637 77147 75671 77175
rect 75699 77147 77009 77175
rect 77037 77147 77071 77175
rect 77099 77147 81509 77175
rect 81537 77147 81571 77175
rect 81599 77147 84485 77175
rect 84513 77147 84547 77175
rect 84575 77147 84609 77175
rect 84637 77147 84671 77175
rect 84699 77147 86009 77175
rect 86037 77147 86071 77175
rect 86099 77147 90509 77175
rect 90537 77147 90571 77175
rect 90599 77147 95009 77175
rect 95037 77147 95071 77175
rect 95099 77147 99509 77175
rect 99537 77147 99571 77175
rect 99599 77147 104009 77175
rect 104037 77147 104071 77175
rect 104099 77147 108509 77175
rect 108537 77147 108571 77175
rect 108599 77147 113009 77175
rect 113037 77147 113071 77175
rect 113099 77147 117509 77175
rect 117537 77147 117571 77175
rect 117599 77147 120485 77175
rect 120513 77147 120547 77175
rect 120575 77147 120609 77175
rect 120637 77147 120671 77175
rect 120699 77147 129485 77175
rect 129513 77147 129547 77175
rect 129575 77147 129609 77175
rect 129637 77147 129671 77175
rect 129699 77147 138485 77175
rect 138513 77147 138547 77175
rect 138575 77147 138609 77175
rect 138637 77147 138671 77175
rect 138699 77147 147485 77175
rect 147513 77147 147547 77175
rect 147575 77147 147609 77175
rect 147637 77147 147671 77175
rect 147699 77147 156485 77175
rect 156513 77147 156547 77175
rect 156575 77147 156609 77175
rect 156637 77147 156671 77175
rect 156699 77147 165485 77175
rect 165513 77147 165547 77175
rect 165575 77147 165609 77175
rect 165637 77147 165671 77175
rect 165699 77147 174485 77175
rect 174513 77147 174547 77175
rect 174575 77147 174609 77175
rect 174637 77147 174671 77175
rect 174699 77147 183485 77175
rect 183513 77147 183547 77175
rect 183575 77147 183609 77175
rect 183637 77147 183671 77175
rect 183699 77147 192485 77175
rect 192513 77147 192547 77175
rect 192575 77147 192609 77175
rect 192637 77147 192671 77175
rect 192699 77147 201485 77175
rect 201513 77147 201547 77175
rect 201575 77147 201609 77175
rect 201637 77147 201671 77175
rect 201699 77147 210485 77175
rect 210513 77147 210547 77175
rect 210575 77147 210609 77175
rect 210637 77147 210671 77175
rect 210699 77147 219485 77175
rect 219513 77147 219547 77175
rect 219575 77147 219609 77175
rect 219637 77147 219671 77175
rect 219699 77147 228485 77175
rect 228513 77147 228547 77175
rect 228575 77147 228609 77175
rect 228637 77147 228671 77175
rect 228699 77147 237485 77175
rect 237513 77147 237547 77175
rect 237575 77147 237609 77175
rect 237637 77147 237671 77175
rect 237699 77147 246485 77175
rect 246513 77147 246547 77175
rect 246575 77147 246609 77175
rect 246637 77147 246671 77175
rect 246699 77147 255485 77175
rect 255513 77147 255547 77175
rect 255575 77147 255609 77175
rect 255637 77147 255671 77175
rect 255699 77147 264485 77175
rect 264513 77147 264547 77175
rect 264575 77147 264609 77175
rect 264637 77147 264671 77175
rect 264699 77147 273485 77175
rect 273513 77147 273547 77175
rect 273575 77147 273609 77175
rect 273637 77147 273671 77175
rect 273699 77147 282485 77175
rect 282513 77147 282547 77175
rect 282575 77147 282609 77175
rect 282637 77147 282671 77175
rect 282699 77147 291485 77175
rect 291513 77147 291547 77175
rect 291575 77147 291609 77175
rect 291637 77147 291671 77175
rect 291699 77147 298728 77175
rect 298756 77147 298790 77175
rect 298818 77147 298852 77175
rect 298880 77147 298914 77175
rect 298942 77147 298990 77175
rect -958 77113 298990 77147
rect -958 77085 -910 77113
rect -882 77085 -848 77113
rect -820 77085 -786 77113
rect -758 77085 -724 77113
rect -696 77085 3485 77113
rect 3513 77085 3547 77113
rect 3575 77085 3609 77113
rect 3637 77085 3671 77113
rect 3699 77085 12485 77113
rect 12513 77085 12547 77113
rect 12575 77085 12609 77113
rect 12637 77085 12671 77113
rect 12699 77085 21485 77113
rect 21513 77085 21547 77113
rect 21575 77085 21609 77113
rect 21637 77085 21671 77113
rect 21699 77085 30485 77113
rect 30513 77085 30547 77113
rect 30575 77085 30609 77113
rect 30637 77085 30671 77113
rect 30699 77085 39485 77113
rect 39513 77085 39547 77113
rect 39575 77085 39609 77113
rect 39637 77085 39671 77113
rect 39699 77085 48485 77113
rect 48513 77085 48547 77113
rect 48575 77085 48609 77113
rect 48637 77085 48671 77113
rect 48699 77085 54509 77113
rect 54537 77085 54571 77113
rect 54599 77085 57485 77113
rect 57513 77085 57547 77113
rect 57575 77085 57609 77113
rect 57637 77085 57671 77113
rect 57699 77085 59009 77113
rect 59037 77085 59071 77113
rect 59099 77085 63509 77113
rect 63537 77085 63571 77113
rect 63599 77085 66485 77113
rect 66513 77085 66547 77113
rect 66575 77085 66609 77113
rect 66637 77085 66671 77113
rect 66699 77085 68009 77113
rect 68037 77085 68071 77113
rect 68099 77085 72509 77113
rect 72537 77085 72571 77113
rect 72599 77085 75485 77113
rect 75513 77085 75547 77113
rect 75575 77085 75609 77113
rect 75637 77085 75671 77113
rect 75699 77085 77009 77113
rect 77037 77085 77071 77113
rect 77099 77085 81509 77113
rect 81537 77085 81571 77113
rect 81599 77085 84485 77113
rect 84513 77085 84547 77113
rect 84575 77085 84609 77113
rect 84637 77085 84671 77113
rect 84699 77085 86009 77113
rect 86037 77085 86071 77113
rect 86099 77085 90509 77113
rect 90537 77085 90571 77113
rect 90599 77085 95009 77113
rect 95037 77085 95071 77113
rect 95099 77085 99509 77113
rect 99537 77085 99571 77113
rect 99599 77085 104009 77113
rect 104037 77085 104071 77113
rect 104099 77085 108509 77113
rect 108537 77085 108571 77113
rect 108599 77085 113009 77113
rect 113037 77085 113071 77113
rect 113099 77085 117509 77113
rect 117537 77085 117571 77113
rect 117599 77085 120485 77113
rect 120513 77085 120547 77113
rect 120575 77085 120609 77113
rect 120637 77085 120671 77113
rect 120699 77085 129485 77113
rect 129513 77085 129547 77113
rect 129575 77085 129609 77113
rect 129637 77085 129671 77113
rect 129699 77085 138485 77113
rect 138513 77085 138547 77113
rect 138575 77085 138609 77113
rect 138637 77085 138671 77113
rect 138699 77085 147485 77113
rect 147513 77085 147547 77113
rect 147575 77085 147609 77113
rect 147637 77085 147671 77113
rect 147699 77085 156485 77113
rect 156513 77085 156547 77113
rect 156575 77085 156609 77113
rect 156637 77085 156671 77113
rect 156699 77085 165485 77113
rect 165513 77085 165547 77113
rect 165575 77085 165609 77113
rect 165637 77085 165671 77113
rect 165699 77085 174485 77113
rect 174513 77085 174547 77113
rect 174575 77085 174609 77113
rect 174637 77085 174671 77113
rect 174699 77085 183485 77113
rect 183513 77085 183547 77113
rect 183575 77085 183609 77113
rect 183637 77085 183671 77113
rect 183699 77085 192485 77113
rect 192513 77085 192547 77113
rect 192575 77085 192609 77113
rect 192637 77085 192671 77113
rect 192699 77085 201485 77113
rect 201513 77085 201547 77113
rect 201575 77085 201609 77113
rect 201637 77085 201671 77113
rect 201699 77085 210485 77113
rect 210513 77085 210547 77113
rect 210575 77085 210609 77113
rect 210637 77085 210671 77113
rect 210699 77085 219485 77113
rect 219513 77085 219547 77113
rect 219575 77085 219609 77113
rect 219637 77085 219671 77113
rect 219699 77085 228485 77113
rect 228513 77085 228547 77113
rect 228575 77085 228609 77113
rect 228637 77085 228671 77113
rect 228699 77085 237485 77113
rect 237513 77085 237547 77113
rect 237575 77085 237609 77113
rect 237637 77085 237671 77113
rect 237699 77085 246485 77113
rect 246513 77085 246547 77113
rect 246575 77085 246609 77113
rect 246637 77085 246671 77113
rect 246699 77085 255485 77113
rect 255513 77085 255547 77113
rect 255575 77085 255609 77113
rect 255637 77085 255671 77113
rect 255699 77085 264485 77113
rect 264513 77085 264547 77113
rect 264575 77085 264609 77113
rect 264637 77085 264671 77113
rect 264699 77085 273485 77113
rect 273513 77085 273547 77113
rect 273575 77085 273609 77113
rect 273637 77085 273671 77113
rect 273699 77085 282485 77113
rect 282513 77085 282547 77113
rect 282575 77085 282609 77113
rect 282637 77085 282671 77113
rect 282699 77085 291485 77113
rect 291513 77085 291547 77113
rect 291575 77085 291609 77113
rect 291637 77085 291671 77113
rect 291699 77085 298728 77113
rect 298756 77085 298790 77113
rect 298818 77085 298852 77113
rect 298880 77085 298914 77113
rect 298942 77085 298990 77113
rect -958 77051 298990 77085
rect -958 77023 -910 77051
rect -882 77023 -848 77051
rect -820 77023 -786 77051
rect -758 77023 -724 77051
rect -696 77023 3485 77051
rect 3513 77023 3547 77051
rect 3575 77023 3609 77051
rect 3637 77023 3671 77051
rect 3699 77023 12485 77051
rect 12513 77023 12547 77051
rect 12575 77023 12609 77051
rect 12637 77023 12671 77051
rect 12699 77023 21485 77051
rect 21513 77023 21547 77051
rect 21575 77023 21609 77051
rect 21637 77023 21671 77051
rect 21699 77023 30485 77051
rect 30513 77023 30547 77051
rect 30575 77023 30609 77051
rect 30637 77023 30671 77051
rect 30699 77023 39485 77051
rect 39513 77023 39547 77051
rect 39575 77023 39609 77051
rect 39637 77023 39671 77051
rect 39699 77023 48485 77051
rect 48513 77023 48547 77051
rect 48575 77023 48609 77051
rect 48637 77023 48671 77051
rect 48699 77023 54509 77051
rect 54537 77023 54571 77051
rect 54599 77023 57485 77051
rect 57513 77023 57547 77051
rect 57575 77023 57609 77051
rect 57637 77023 57671 77051
rect 57699 77023 59009 77051
rect 59037 77023 59071 77051
rect 59099 77023 63509 77051
rect 63537 77023 63571 77051
rect 63599 77023 66485 77051
rect 66513 77023 66547 77051
rect 66575 77023 66609 77051
rect 66637 77023 66671 77051
rect 66699 77023 68009 77051
rect 68037 77023 68071 77051
rect 68099 77023 72509 77051
rect 72537 77023 72571 77051
rect 72599 77023 75485 77051
rect 75513 77023 75547 77051
rect 75575 77023 75609 77051
rect 75637 77023 75671 77051
rect 75699 77023 77009 77051
rect 77037 77023 77071 77051
rect 77099 77023 81509 77051
rect 81537 77023 81571 77051
rect 81599 77023 84485 77051
rect 84513 77023 84547 77051
rect 84575 77023 84609 77051
rect 84637 77023 84671 77051
rect 84699 77023 86009 77051
rect 86037 77023 86071 77051
rect 86099 77023 90509 77051
rect 90537 77023 90571 77051
rect 90599 77023 95009 77051
rect 95037 77023 95071 77051
rect 95099 77023 99509 77051
rect 99537 77023 99571 77051
rect 99599 77023 104009 77051
rect 104037 77023 104071 77051
rect 104099 77023 108509 77051
rect 108537 77023 108571 77051
rect 108599 77023 113009 77051
rect 113037 77023 113071 77051
rect 113099 77023 117509 77051
rect 117537 77023 117571 77051
rect 117599 77023 120485 77051
rect 120513 77023 120547 77051
rect 120575 77023 120609 77051
rect 120637 77023 120671 77051
rect 120699 77023 129485 77051
rect 129513 77023 129547 77051
rect 129575 77023 129609 77051
rect 129637 77023 129671 77051
rect 129699 77023 138485 77051
rect 138513 77023 138547 77051
rect 138575 77023 138609 77051
rect 138637 77023 138671 77051
rect 138699 77023 147485 77051
rect 147513 77023 147547 77051
rect 147575 77023 147609 77051
rect 147637 77023 147671 77051
rect 147699 77023 156485 77051
rect 156513 77023 156547 77051
rect 156575 77023 156609 77051
rect 156637 77023 156671 77051
rect 156699 77023 165485 77051
rect 165513 77023 165547 77051
rect 165575 77023 165609 77051
rect 165637 77023 165671 77051
rect 165699 77023 174485 77051
rect 174513 77023 174547 77051
rect 174575 77023 174609 77051
rect 174637 77023 174671 77051
rect 174699 77023 183485 77051
rect 183513 77023 183547 77051
rect 183575 77023 183609 77051
rect 183637 77023 183671 77051
rect 183699 77023 192485 77051
rect 192513 77023 192547 77051
rect 192575 77023 192609 77051
rect 192637 77023 192671 77051
rect 192699 77023 201485 77051
rect 201513 77023 201547 77051
rect 201575 77023 201609 77051
rect 201637 77023 201671 77051
rect 201699 77023 210485 77051
rect 210513 77023 210547 77051
rect 210575 77023 210609 77051
rect 210637 77023 210671 77051
rect 210699 77023 219485 77051
rect 219513 77023 219547 77051
rect 219575 77023 219609 77051
rect 219637 77023 219671 77051
rect 219699 77023 228485 77051
rect 228513 77023 228547 77051
rect 228575 77023 228609 77051
rect 228637 77023 228671 77051
rect 228699 77023 237485 77051
rect 237513 77023 237547 77051
rect 237575 77023 237609 77051
rect 237637 77023 237671 77051
rect 237699 77023 246485 77051
rect 246513 77023 246547 77051
rect 246575 77023 246609 77051
rect 246637 77023 246671 77051
rect 246699 77023 255485 77051
rect 255513 77023 255547 77051
rect 255575 77023 255609 77051
rect 255637 77023 255671 77051
rect 255699 77023 264485 77051
rect 264513 77023 264547 77051
rect 264575 77023 264609 77051
rect 264637 77023 264671 77051
rect 264699 77023 273485 77051
rect 273513 77023 273547 77051
rect 273575 77023 273609 77051
rect 273637 77023 273671 77051
rect 273699 77023 282485 77051
rect 282513 77023 282547 77051
rect 282575 77023 282609 77051
rect 282637 77023 282671 77051
rect 282699 77023 291485 77051
rect 291513 77023 291547 77051
rect 291575 77023 291609 77051
rect 291637 77023 291671 77051
rect 291699 77023 298728 77051
rect 298756 77023 298790 77051
rect 298818 77023 298852 77051
rect 298880 77023 298914 77051
rect 298942 77023 298990 77051
rect -958 76989 298990 77023
rect -958 76961 -910 76989
rect -882 76961 -848 76989
rect -820 76961 -786 76989
rect -758 76961 -724 76989
rect -696 76961 3485 76989
rect 3513 76961 3547 76989
rect 3575 76961 3609 76989
rect 3637 76961 3671 76989
rect 3699 76961 12485 76989
rect 12513 76961 12547 76989
rect 12575 76961 12609 76989
rect 12637 76961 12671 76989
rect 12699 76961 21485 76989
rect 21513 76961 21547 76989
rect 21575 76961 21609 76989
rect 21637 76961 21671 76989
rect 21699 76961 30485 76989
rect 30513 76961 30547 76989
rect 30575 76961 30609 76989
rect 30637 76961 30671 76989
rect 30699 76961 39485 76989
rect 39513 76961 39547 76989
rect 39575 76961 39609 76989
rect 39637 76961 39671 76989
rect 39699 76961 48485 76989
rect 48513 76961 48547 76989
rect 48575 76961 48609 76989
rect 48637 76961 48671 76989
rect 48699 76961 54509 76989
rect 54537 76961 54571 76989
rect 54599 76961 57485 76989
rect 57513 76961 57547 76989
rect 57575 76961 57609 76989
rect 57637 76961 57671 76989
rect 57699 76961 59009 76989
rect 59037 76961 59071 76989
rect 59099 76961 63509 76989
rect 63537 76961 63571 76989
rect 63599 76961 66485 76989
rect 66513 76961 66547 76989
rect 66575 76961 66609 76989
rect 66637 76961 66671 76989
rect 66699 76961 68009 76989
rect 68037 76961 68071 76989
rect 68099 76961 72509 76989
rect 72537 76961 72571 76989
rect 72599 76961 75485 76989
rect 75513 76961 75547 76989
rect 75575 76961 75609 76989
rect 75637 76961 75671 76989
rect 75699 76961 77009 76989
rect 77037 76961 77071 76989
rect 77099 76961 81509 76989
rect 81537 76961 81571 76989
rect 81599 76961 84485 76989
rect 84513 76961 84547 76989
rect 84575 76961 84609 76989
rect 84637 76961 84671 76989
rect 84699 76961 86009 76989
rect 86037 76961 86071 76989
rect 86099 76961 90509 76989
rect 90537 76961 90571 76989
rect 90599 76961 95009 76989
rect 95037 76961 95071 76989
rect 95099 76961 99509 76989
rect 99537 76961 99571 76989
rect 99599 76961 104009 76989
rect 104037 76961 104071 76989
rect 104099 76961 108509 76989
rect 108537 76961 108571 76989
rect 108599 76961 113009 76989
rect 113037 76961 113071 76989
rect 113099 76961 117509 76989
rect 117537 76961 117571 76989
rect 117599 76961 120485 76989
rect 120513 76961 120547 76989
rect 120575 76961 120609 76989
rect 120637 76961 120671 76989
rect 120699 76961 129485 76989
rect 129513 76961 129547 76989
rect 129575 76961 129609 76989
rect 129637 76961 129671 76989
rect 129699 76961 138485 76989
rect 138513 76961 138547 76989
rect 138575 76961 138609 76989
rect 138637 76961 138671 76989
rect 138699 76961 147485 76989
rect 147513 76961 147547 76989
rect 147575 76961 147609 76989
rect 147637 76961 147671 76989
rect 147699 76961 156485 76989
rect 156513 76961 156547 76989
rect 156575 76961 156609 76989
rect 156637 76961 156671 76989
rect 156699 76961 165485 76989
rect 165513 76961 165547 76989
rect 165575 76961 165609 76989
rect 165637 76961 165671 76989
rect 165699 76961 174485 76989
rect 174513 76961 174547 76989
rect 174575 76961 174609 76989
rect 174637 76961 174671 76989
rect 174699 76961 183485 76989
rect 183513 76961 183547 76989
rect 183575 76961 183609 76989
rect 183637 76961 183671 76989
rect 183699 76961 192485 76989
rect 192513 76961 192547 76989
rect 192575 76961 192609 76989
rect 192637 76961 192671 76989
rect 192699 76961 201485 76989
rect 201513 76961 201547 76989
rect 201575 76961 201609 76989
rect 201637 76961 201671 76989
rect 201699 76961 210485 76989
rect 210513 76961 210547 76989
rect 210575 76961 210609 76989
rect 210637 76961 210671 76989
rect 210699 76961 219485 76989
rect 219513 76961 219547 76989
rect 219575 76961 219609 76989
rect 219637 76961 219671 76989
rect 219699 76961 228485 76989
rect 228513 76961 228547 76989
rect 228575 76961 228609 76989
rect 228637 76961 228671 76989
rect 228699 76961 237485 76989
rect 237513 76961 237547 76989
rect 237575 76961 237609 76989
rect 237637 76961 237671 76989
rect 237699 76961 246485 76989
rect 246513 76961 246547 76989
rect 246575 76961 246609 76989
rect 246637 76961 246671 76989
rect 246699 76961 255485 76989
rect 255513 76961 255547 76989
rect 255575 76961 255609 76989
rect 255637 76961 255671 76989
rect 255699 76961 264485 76989
rect 264513 76961 264547 76989
rect 264575 76961 264609 76989
rect 264637 76961 264671 76989
rect 264699 76961 273485 76989
rect 273513 76961 273547 76989
rect 273575 76961 273609 76989
rect 273637 76961 273671 76989
rect 273699 76961 282485 76989
rect 282513 76961 282547 76989
rect 282575 76961 282609 76989
rect 282637 76961 282671 76989
rect 282699 76961 291485 76989
rect 291513 76961 291547 76989
rect 291575 76961 291609 76989
rect 291637 76961 291671 76989
rect 291699 76961 298728 76989
rect 298756 76961 298790 76989
rect 298818 76961 298852 76989
rect 298880 76961 298914 76989
rect 298942 76961 298990 76989
rect -958 76913 298990 76961
rect -958 74175 298990 74223
rect -958 74147 -430 74175
rect -402 74147 -368 74175
rect -340 74147 -306 74175
rect -278 74147 -244 74175
rect -216 74147 1625 74175
rect 1653 74147 1687 74175
rect 1715 74147 1749 74175
rect 1777 74147 1811 74175
rect 1839 74147 10625 74175
rect 10653 74147 10687 74175
rect 10715 74147 10749 74175
rect 10777 74147 10811 74175
rect 10839 74147 19625 74175
rect 19653 74147 19687 74175
rect 19715 74147 19749 74175
rect 19777 74147 19811 74175
rect 19839 74147 28625 74175
rect 28653 74147 28687 74175
rect 28715 74147 28749 74175
rect 28777 74147 28811 74175
rect 28839 74147 37625 74175
rect 37653 74147 37687 74175
rect 37715 74147 37749 74175
rect 37777 74147 37811 74175
rect 37839 74147 46625 74175
rect 46653 74147 46687 74175
rect 46715 74147 46749 74175
rect 46777 74147 46811 74175
rect 46839 74147 52259 74175
rect 52287 74147 52321 74175
rect 52349 74147 55625 74175
rect 55653 74147 55687 74175
rect 55715 74147 55749 74175
rect 55777 74147 55811 74175
rect 55839 74147 56759 74175
rect 56787 74147 56821 74175
rect 56849 74147 61259 74175
rect 61287 74147 61321 74175
rect 61349 74147 64625 74175
rect 64653 74147 64687 74175
rect 64715 74147 64749 74175
rect 64777 74147 64811 74175
rect 64839 74147 65759 74175
rect 65787 74147 65821 74175
rect 65849 74147 70259 74175
rect 70287 74147 70321 74175
rect 70349 74147 73625 74175
rect 73653 74147 73687 74175
rect 73715 74147 73749 74175
rect 73777 74147 73811 74175
rect 73839 74147 74759 74175
rect 74787 74147 74821 74175
rect 74849 74147 79259 74175
rect 79287 74147 79321 74175
rect 79349 74147 82625 74175
rect 82653 74147 82687 74175
rect 82715 74147 82749 74175
rect 82777 74147 82811 74175
rect 82839 74147 83759 74175
rect 83787 74147 83821 74175
rect 83849 74147 88259 74175
rect 88287 74147 88321 74175
rect 88349 74147 91625 74175
rect 91653 74147 91687 74175
rect 91715 74147 91749 74175
rect 91777 74147 91811 74175
rect 91839 74147 92759 74175
rect 92787 74147 92821 74175
rect 92849 74147 97259 74175
rect 97287 74147 97321 74175
rect 97349 74147 101759 74175
rect 101787 74147 101821 74175
rect 101849 74147 106259 74175
rect 106287 74147 106321 74175
rect 106349 74147 110759 74175
rect 110787 74147 110821 74175
rect 110849 74147 115259 74175
rect 115287 74147 115321 74175
rect 115349 74147 127625 74175
rect 127653 74147 127687 74175
rect 127715 74147 127749 74175
rect 127777 74147 127811 74175
rect 127839 74147 136625 74175
rect 136653 74147 136687 74175
rect 136715 74147 136749 74175
rect 136777 74147 136811 74175
rect 136839 74147 145625 74175
rect 145653 74147 145687 74175
rect 145715 74147 145749 74175
rect 145777 74147 145811 74175
rect 145839 74147 154625 74175
rect 154653 74147 154687 74175
rect 154715 74147 154749 74175
rect 154777 74147 154811 74175
rect 154839 74147 163625 74175
rect 163653 74147 163687 74175
rect 163715 74147 163749 74175
rect 163777 74147 163811 74175
rect 163839 74147 172625 74175
rect 172653 74147 172687 74175
rect 172715 74147 172749 74175
rect 172777 74147 172811 74175
rect 172839 74147 181625 74175
rect 181653 74147 181687 74175
rect 181715 74147 181749 74175
rect 181777 74147 181811 74175
rect 181839 74147 190625 74175
rect 190653 74147 190687 74175
rect 190715 74147 190749 74175
rect 190777 74147 190811 74175
rect 190839 74147 199625 74175
rect 199653 74147 199687 74175
rect 199715 74147 199749 74175
rect 199777 74147 199811 74175
rect 199839 74147 208625 74175
rect 208653 74147 208687 74175
rect 208715 74147 208749 74175
rect 208777 74147 208811 74175
rect 208839 74147 217625 74175
rect 217653 74147 217687 74175
rect 217715 74147 217749 74175
rect 217777 74147 217811 74175
rect 217839 74147 226625 74175
rect 226653 74147 226687 74175
rect 226715 74147 226749 74175
rect 226777 74147 226811 74175
rect 226839 74147 235625 74175
rect 235653 74147 235687 74175
rect 235715 74147 235749 74175
rect 235777 74147 235811 74175
rect 235839 74147 244625 74175
rect 244653 74147 244687 74175
rect 244715 74147 244749 74175
rect 244777 74147 244811 74175
rect 244839 74147 253625 74175
rect 253653 74147 253687 74175
rect 253715 74147 253749 74175
rect 253777 74147 253811 74175
rect 253839 74147 262625 74175
rect 262653 74147 262687 74175
rect 262715 74147 262749 74175
rect 262777 74147 262811 74175
rect 262839 74147 271625 74175
rect 271653 74147 271687 74175
rect 271715 74147 271749 74175
rect 271777 74147 271811 74175
rect 271839 74147 280625 74175
rect 280653 74147 280687 74175
rect 280715 74147 280749 74175
rect 280777 74147 280811 74175
rect 280839 74147 289625 74175
rect 289653 74147 289687 74175
rect 289715 74147 289749 74175
rect 289777 74147 289811 74175
rect 289839 74147 298248 74175
rect 298276 74147 298310 74175
rect 298338 74147 298372 74175
rect 298400 74147 298434 74175
rect 298462 74147 298990 74175
rect -958 74113 298990 74147
rect -958 74085 -430 74113
rect -402 74085 -368 74113
rect -340 74085 -306 74113
rect -278 74085 -244 74113
rect -216 74085 1625 74113
rect 1653 74085 1687 74113
rect 1715 74085 1749 74113
rect 1777 74085 1811 74113
rect 1839 74085 10625 74113
rect 10653 74085 10687 74113
rect 10715 74085 10749 74113
rect 10777 74085 10811 74113
rect 10839 74085 19625 74113
rect 19653 74085 19687 74113
rect 19715 74085 19749 74113
rect 19777 74085 19811 74113
rect 19839 74085 28625 74113
rect 28653 74085 28687 74113
rect 28715 74085 28749 74113
rect 28777 74085 28811 74113
rect 28839 74085 37625 74113
rect 37653 74085 37687 74113
rect 37715 74085 37749 74113
rect 37777 74085 37811 74113
rect 37839 74085 46625 74113
rect 46653 74085 46687 74113
rect 46715 74085 46749 74113
rect 46777 74085 46811 74113
rect 46839 74085 52259 74113
rect 52287 74085 52321 74113
rect 52349 74085 55625 74113
rect 55653 74085 55687 74113
rect 55715 74085 55749 74113
rect 55777 74085 55811 74113
rect 55839 74085 56759 74113
rect 56787 74085 56821 74113
rect 56849 74085 61259 74113
rect 61287 74085 61321 74113
rect 61349 74085 64625 74113
rect 64653 74085 64687 74113
rect 64715 74085 64749 74113
rect 64777 74085 64811 74113
rect 64839 74085 65759 74113
rect 65787 74085 65821 74113
rect 65849 74085 70259 74113
rect 70287 74085 70321 74113
rect 70349 74085 73625 74113
rect 73653 74085 73687 74113
rect 73715 74085 73749 74113
rect 73777 74085 73811 74113
rect 73839 74085 74759 74113
rect 74787 74085 74821 74113
rect 74849 74085 79259 74113
rect 79287 74085 79321 74113
rect 79349 74085 82625 74113
rect 82653 74085 82687 74113
rect 82715 74085 82749 74113
rect 82777 74085 82811 74113
rect 82839 74085 83759 74113
rect 83787 74085 83821 74113
rect 83849 74085 88259 74113
rect 88287 74085 88321 74113
rect 88349 74085 91625 74113
rect 91653 74085 91687 74113
rect 91715 74085 91749 74113
rect 91777 74085 91811 74113
rect 91839 74085 92759 74113
rect 92787 74085 92821 74113
rect 92849 74085 97259 74113
rect 97287 74085 97321 74113
rect 97349 74085 101759 74113
rect 101787 74085 101821 74113
rect 101849 74085 106259 74113
rect 106287 74085 106321 74113
rect 106349 74085 110759 74113
rect 110787 74085 110821 74113
rect 110849 74085 115259 74113
rect 115287 74085 115321 74113
rect 115349 74085 127625 74113
rect 127653 74085 127687 74113
rect 127715 74085 127749 74113
rect 127777 74085 127811 74113
rect 127839 74085 136625 74113
rect 136653 74085 136687 74113
rect 136715 74085 136749 74113
rect 136777 74085 136811 74113
rect 136839 74085 145625 74113
rect 145653 74085 145687 74113
rect 145715 74085 145749 74113
rect 145777 74085 145811 74113
rect 145839 74085 154625 74113
rect 154653 74085 154687 74113
rect 154715 74085 154749 74113
rect 154777 74085 154811 74113
rect 154839 74085 163625 74113
rect 163653 74085 163687 74113
rect 163715 74085 163749 74113
rect 163777 74085 163811 74113
rect 163839 74085 172625 74113
rect 172653 74085 172687 74113
rect 172715 74085 172749 74113
rect 172777 74085 172811 74113
rect 172839 74085 181625 74113
rect 181653 74085 181687 74113
rect 181715 74085 181749 74113
rect 181777 74085 181811 74113
rect 181839 74085 190625 74113
rect 190653 74085 190687 74113
rect 190715 74085 190749 74113
rect 190777 74085 190811 74113
rect 190839 74085 199625 74113
rect 199653 74085 199687 74113
rect 199715 74085 199749 74113
rect 199777 74085 199811 74113
rect 199839 74085 208625 74113
rect 208653 74085 208687 74113
rect 208715 74085 208749 74113
rect 208777 74085 208811 74113
rect 208839 74085 217625 74113
rect 217653 74085 217687 74113
rect 217715 74085 217749 74113
rect 217777 74085 217811 74113
rect 217839 74085 226625 74113
rect 226653 74085 226687 74113
rect 226715 74085 226749 74113
rect 226777 74085 226811 74113
rect 226839 74085 235625 74113
rect 235653 74085 235687 74113
rect 235715 74085 235749 74113
rect 235777 74085 235811 74113
rect 235839 74085 244625 74113
rect 244653 74085 244687 74113
rect 244715 74085 244749 74113
rect 244777 74085 244811 74113
rect 244839 74085 253625 74113
rect 253653 74085 253687 74113
rect 253715 74085 253749 74113
rect 253777 74085 253811 74113
rect 253839 74085 262625 74113
rect 262653 74085 262687 74113
rect 262715 74085 262749 74113
rect 262777 74085 262811 74113
rect 262839 74085 271625 74113
rect 271653 74085 271687 74113
rect 271715 74085 271749 74113
rect 271777 74085 271811 74113
rect 271839 74085 280625 74113
rect 280653 74085 280687 74113
rect 280715 74085 280749 74113
rect 280777 74085 280811 74113
rect 280839 74085 289625 74113
rect 289653 74085 289687 74113
rect 289715 74085 289749 74113
rect 289777 74085 289811 74113
rect 289839 74085 298248 74113
rect 298276 74085 298310 74113
rect 298338 74085 298372 74113
rect 298400 74085 298434 74113
rect 298462 74085 298990 74113
rect -958 74051 298990 74085
rect -958 74023 -430 74051
rect -402 74023 -368 74051
rect -340 74023 -306 74051
rect -278 74023 -244 74051
rect -216 74023 1625 74051
rect 1653 74023 1687 74051
rect 1715 74023 1749 74051
rect 1777 74023 1811 74051
rect 1839 74023 10625 74051
rect 10653 74023 10687 74051
rect 10715 74023 10749 74051
rect 10777 74023 10811 74051
rect 10839 74023 19625 74051
rect 19653 74023 19687 74051
rect 19715 74023 19749 74051
rect 19777 74023 19811 74051
rect 19839 74023 28625 74051
rect 28653 74023 28687 74051
rect 28715 74023 28749 74051
rect 28777 74023 28811 74051
rect 28839 74023 37625 74051
rect 37653 74023 37687 74051
rect 37715 74023 37749 74051
rect 37777 74023 37811 74051
rect 37839 74023 46625 74051
rect 46653 74023 46687 74051
rect 46715 74023 46749 74051
rect 46777 74023 46811 74051
rect 46839 74023 52259 74051
rect 52287 74023 52321 74051
rect 52349 74023 55625 74051
rect 55653 74023 55687 74051
rect 55715 74023 55749 74051
rect 55777 74023 55811 74051
rect 55839 74023 56759 74051
rect 56787 74023 56821 74051
rect 56849 74023 61259 74051
rect 61287 74023 61321 74051
rect 61349 74023 64625 74051
rect 64653 74023 64687 74051
rect 64715 74023 64749 74051
rect 64777 74023 64811 74051
rect 64839 74023 65759 74051
rect 65787 74023 65821 74051
rect 65849 74023 70259 74051
rect 70287 74023 70321 74051
rect 70349 74023 73625 74051
rect 73653 74023 73687 74051
rect 73715 74023 73749 74051
rect 73777 74023 73811 74051
rect 73839 74023 74759 74051
rect 74787 74023 74821 74051
rect 74849 74023 79259 74051
rect 79287 74023 79321 74051
rect 79349 74023 82625 74051
rect 82653 74023 82687 74051
rect 82715 74023 82749 74051
rect 82777 74023 82811 74051
rect 82839 74023 83759 74051
rect 83787 74023 83821 74051
rect 83849 74023 88259 74051
rect 88287 74023 88321 74051
rect 88349 74023 91625 74051
rect 91653 74023 91687 74051
rect 91715 74023 91749 74051
rect 91777 74023 91811 74051
rect 91839 74023 92759 74051
rect 92787 74023 92821 74051
rect 92849 74023 97259 74051
rect 97287 74023 97321 74051
rect 97349 74023 101759 74051
rect 101787 74023 101821 74051
rect 101849 74023 106259 74051
rect 106287 74023 106321 74051
rect 106349 74023 110759 74051
rect 110787 74023 110821 74051
rect 110849 74023 115259 74051
rect 115287 74023 115321 74051
rect 115349 74023 127625 74051
rect 127653 74023 127687 74051
rect 127715 74023 127749 74051
rect 127777 74023 127811 74051
rect 127839 74023 136625 74051
rect 136653 74023 136687 74051
rect 136715 74023 136749 74051
rect 136777 74023 136811 74051
rect 136839 74023 145625 74051
rect 145653 74023 145687 74051
rect 145715 74023 145749 74051
rect 145777 74023 145811 74051
rect 145839 74023 154625 74051
rect 154653 74023 154687 74051
rect 154715 74023 154749 74051
rect 154777 74023 154811 74051
rect 154839 74023 163625 74051
rect 163653 74023 163687 74051
rect 163715 74023 163749 74051
rect 163777 74023 163811 74051
rect 163839 74023 172625 74051
rect 172653 74023 172687 74051
rect 172715 74023 172749 74051
rect 172777 74023 172811 74051
rect 172839 74023 181625 74051
rect 181653 74023 181687 74051
rect 181715 74023 181749 74051
rect 181777 74023 181811 74051
rect 181839 74023 190625 74051
rect 190653 74023 190687 74051
rect 190715 74023 190749 74051
rect 190777 74023 190811 74051
rect 190839 74023 199625 74051
rect 199653 74023 199687 74051
rect 199715 74023 199749 74051
rect 199777 74023 199811 74051
rect 199839 74023 208625 74051
rect 208653 74023 208687 74051
rect 208715 74023 208749 74051
rect 208777 74023 208811 74051
rect 208839 74023 217625 74051
rect 217653 74023 217687 74051
rect 217715 74023 217749 74051
rect 217777 74023 217811 74051
rect 217839 74023 226625 74051
rect 226653 74023 226687 74051
rect 226715 74023 226749 74051
rect 226777 74023 226811 74051
rect 226839 74023 235625 74051
rect 235653 74023 235687 74051
rect 235715 74023 235749 74051
rect 235777 74023 235811 74051
rect 235839 74023 244625 74051
rect 244653 74023 244687 74051
rect 244715 74023 244749 74051
rect 244777 74023 244811 74051
rect 244839 74023 253625 74051
rect 253653 74023 253687 74051
rect 253715 74023 253749 74051
rect 253777 74023 253811 74051
rect 253839 74023 262625 74051
rect 262653 74023 262687 74051
rect 262715 74023 262749 74051
rect 262777 74023 262811 74051
rect 262839 74023 271625 74051
rect 271653 74023 271687 74051
rect 271715 74023 271749 74051
rect 271777 74023 271811 74051
rect 271839 74023 280625 74051
rect 280653 74023 280687 74051
rect 280715 74023 280749 74051
rect 280777 74023 280811 74051
rect 280839 74023 289625 74051
rect 289653 74023 289687 74051
rect 289715 74023 289749 74051
rect 289777 74023 289811 74051
rect 289839 74023 298248 74051
rect 298276 74023 298310 74051
rect 298338 74023 298372 74051
rect 298400 74023 298434 74051
rect 298462 74023 298990 74051
rect -958 73989 298990 74023
rect -958 73961 -430 73989
rect -402 73961 -368 73989
rect -340 73961 -306 73989
rect -278 73961 -244 73989
rect -216 73961 1625 73989
rect 1653 73961 1687 73989
rect 1715 73961 1749 73989
rect 1777 73961 1811 73989
rect 1839 73961 10625 73989
rect 10653 73961 10687 73989
rect 10715 73961 10749 73989
rect 10777 73961 10811 73989
rect 10839 73961 19625 73989
rect 19653 73961 19687 73989
rect 19715 73961 19749 73989
rect 19777 73961 19811 73989
rect 19839 73961 28625 73989
rect 28653 73961 28687 73989
rect 28715 73961 28749 73989
rect 28777 73961 28811 73989
rect 28839 73961 37625 73989
rect 37653 73961 37687 73989
rect 37715 73961 37749 73989
rect 37777 73961 37811 73989
rect 37839 73961 46625 73989
rect 46653 73961 46687 73989
rect 46715 73961 46749 73989
rect 46777 73961 46811 73989
rect 46839 73961 52259 73989
rect 52287 73961 52321 73989
rect 52349 73961 55625 73989
rect 55653 73961 55687 73989
rect 55715 73961 55749 73989
rect 55777 73961 55811 73989
rect 55839 73961 56759 73989
rect 56787 73961 56821 73989
rect 56849 73961 61259 73989
rect 61287 73961 61321 73989
rect 61349 73961 64625 73989
rect 64653 73961 64687 73989
rect 64715 73961 64749 73989
rect 64777 73961 64811 73989
rect 64839 73961 65759 73989
rect 65787 73961 65821 73989
rect 65849 73961 70259 73989
rect 70287 73961 70321 73989
rect 70349 73961 73625 73989
rect 73653 73961 73687 73989
rect 73715 73961 73749 73989
rect 73777 73961 73811 73989
rect 73839 73961 74759 73989
rect 74787 73961 74821 73989
rect 74849 73961 79259 73989
rect 79287 73961 79321 73989
rect 79349 73961 82625 73989
rect 82653 73961 82687 73989
rect 82715 73961 82749 73989
rect 82777 73961 82811 73989
rect 82839 73961 83759 73989
rect 83787 73961 83821 73989
rect 83849 73961 88259 73989
rect 88287 73961 88321 73989
rect 88349 73961 91625 73989
rect 91653 73961 91687 73989
rect 91715 73961 91749 73989
rect 91777 73961 91811 73989
rect 91839 73961 92759 73989
rect 92787 73961 92821 73989
rect 92849 73961 97259 73989
rect 97287 73961 97321 73989
rect 97349 73961 101759 73989
rect 101787 73961 101821 73989
rect 101849 73961 106259 73989
rect 106287 73961 106321 73989
rect 106349 73961 110759 73989
rect 110787 73961 110821 73989
rect 110849 73961 115259 73989
rect 115287 73961 115321 73989
rect 115349 73961 127625 73989
rect 127653 73961 127687 73989
rect 127715 73961 127749 73989
rect 127777 73961 127811 73989
rect 127839 73961 136625 73989
rect 136653 73961 136687 73989
rect 136715 73961 136749 73989
rect 136777 73961 136811 73989
rect 136839 73961 145625 73989
rect 145653 73961 145687 73989
rect 145715 73961 145749 73989
rect 145777 73961 145811 73989
rect 145839 73961 154625 73989
rect 154653 73961 154687 73989
rect 154715 73961 154749 73989
rect 154777 73961 154811 73989
rect 154839 73961 163625 73989
rect 163653 73961 163687 73989
rect 163715 73961 163749 73989
rect 163777 73961 163811 73989
rect 163839 73961 172625 73989
rect 172653 73961 172687 73989
rect 172715 73961 172749 73989
rect 172777 73961 172811 73989
rect 172839 73961 181625 73989
rect 181653 73961 181687 73989
rect 181715 73961 181749 73989
rect 181777 73961 181811 73989
rect 181839 73961 190625 73989
rect 190653 73961 190687 73989
rect 190715 73961 190749 73989
rect 190777 73961 190811 73989
rect 190839 73961 199625 73989
rect 199653 73961 199687 73989
rect 199715 73961 199749 73989
rect 199777 73961 199811 73989
rect 199839 73961 208625 73989
rect 208653 73961 208687 73989
rect 208715 73961 208749 73989
rect 208777 73961 208811 73989
rect 208839 73961 217625 73989
rect 217653 73961 217687 73989
rect 217715 73961 217749 73989
rect 217777 73961 217811 73989
rect 217839 73961 226625 73989
rect 226653 73961 226687 73989
rect 226715 73961 226749 73989
rect 226777 73961 226811 73989
rect 226839 73961 235625 73989
rect 235653 73961 235687 73989
rect 235715 73961 235749 73989
rect 235777 73961 235811 73989
rect 235839 73961 244625 73989
rect 244653 73961 244687 73989
rect 244715 73961 244749 73989
rect 244777 73961 244811 73989
rect 244839 73961 253625 73989
rect 253653 73961 253687 73989
rect 253715 73961 253749 73989
rect 253777 73961 253811 73989
rect 253839 73961 262625 73989
rect 262653 73961 262687 73989
rect 262715 73961 262749 73989
rect 262777 73961 262811 73989
rect 262839 73961 271625 73989
rect 271653 73961 271687 73989
rect 271715 73961 271749 73989
rect 271777 73961 271811 73989
rect 271839 73961 280625 73989
rect 280653 73961 280687 73989
rect 280715 73961 280749 73989
rect 280777 73961 280811 73989
rect 280839 73961 289625 73989
rect 289653 73961 289687 73989
rect 289715 73961 289749 73989
rect 289777 73961 289811 73989
rect 289839 73961 298248 73989
rect 298276 73961 298310 73989
rect 298338 73961 298372 73989
rect 298400 73961 298434 73989
rect 298462 73961 298990 73989
rect -958 73913 298990 73961
rect -958 68175 298990 68223
rect -958 68147 -910 68175
rect -882 68147 -848 68175
rect -820 68147 -786 68175
rect -758 68147 -724 68175
rect -696 68147 3485 68175
rect 3513 68147 3547 68175
rect 3575 68147 3609 68175
rect 3637 68147 3671 68175
rect 3699 68147 12485 68175
rect 12513 68147 12547 68175
rect 12575 68147 12609 68175
rect 12637 68147 12671 68175
rect 12699 68147 21485 68175
rect 21513 68147 21547 68175
rect 21575 68147 21609 68175
rect 21637 68147 21671 68175
rect 21699 68147 30485 68175
rect 30513 68147 30547 68175
rect 30575 68147 30609 68175
rect 30637 68147 30671 68175
rect 30699 68147 39485 68175
rect 39513 68147 39547 68175
rect 39575 68147 39609 68175
rect 39637 68147 39671 68175
rect 39699 68147 48485 68175
rect 48513 68147 48547 68175
rect 48575 68147 48609 68175
rect 48637 68147 48671 68175
rect 48699 68147 54509 68175
rect 54537 68147 54571 68175
rect 54599 68147 57485 68175
rect 57513 68147 57547 68175
rect 57575 68147 57609 68175
rect 57637 68147 57671 68175
rect 57699 68147 59009 68175
rect 59037 68147 59071 68175
rect 59099 68147 63509 68175
rect 63537 68147 63571 68175
rect 63599 68147 66485 68175
rect 66513 68147 66547 68175
rect 66575 68147 66609 68175
rect 66637 68147 66671 68175
rect 66699 68147 68009 68175
rect 68037 68147 68071 68175
rect 68099 68147 72509 68175
rect 72537 68147 72571 68175
rect 72599 68147 75485 68175
rect 75513 68147 75547 68175
rect 75575 68147 75609 68175
rect 75637 68147 75671 68175
rect 75699 68147 77009 68175
rect 77037 68147 77071 68175
rect 77099 68147 81509 68175
rect 81537 68147 81571 68175
rect 81599 68147 84485 68175
rect 84513 68147 84547 68175
rect 84575 68147 84609 68175
rect 84637 68147 84671 68175
rect 84699 68147 86009 68175
rect 86037 68147 86071 68175
rect 86099 68147 90509 68175
rect 90537 68147 90571 68175
rect 90599 68147 95009 68175
rect 95037 68147 95071 68175
rect 95099 68147 99509 68175
rect 99537 68147 99571 68175
rect 99599 68147 104009 68175
rect 104037 68147 104071 68175
rect 104099 68147 108509 68175
rect 108537 68147 108571 68175
rect 108599 68147 113009 68175
rect 113037 68147 113071 68175
rect 113099 68147 117509 68175
rect 117537 68147 117571 68175
rect 117599 68147 120485 68175
rect 120513 68147 120547 68175
rect 120575 68147 120609 68175
rect 120637 68147 120671 68175
rect 120699 68147 129485 68175
rect 129513 68147 129547 68175
rect 129575 68147 129609 68175
rect 129637 68147 129671 68175
rect 129699 68147 138485 68175
rect 138513 68147 138547 68175
rect 138575 68147 138609 68175
rect 138637 68147 138671 68175
rect 138699 68147 147485 68175
rect 147513 68147 147547 68175
rect 147575 68147 147609 68175
rect 147637 68147 147671 68175
rect 147699 68147 156485 68175
rect 156513 68147 156547 68175
rect 156575 68147 156609 68175
rect 156637 68147 156671 68175
rect 156699 68147 165485 68175
rect 165513 68147 165547 68175
rect 165575 68147 165609 68175
rect 165637 68147 165671 68175
rect 165699 68147 174485 68175
rect 174513 68147 174547 68175
rect 174575 68147 174609 68175
rect 174637 68147 174671 68175
rect 174699 68147 183485 68175
rect 183513 68147 183547 68175
rect 183575 68147 183609 68175
rect 183637 68147 183671 68175
rect 183699 68147 192485 68175
rect 192513 68147 192547 68175
rect 192575 68147 192609 68175
rect 192637 68147 192671 68175
rect 192699 68147 201485 68175
rect 201513 68147 201547 68175
rect 201575 68147 201609 68175
rect 201637 68147 201671 68175
rect 201699 68147 210485 68175
rect 210513 68147 210547 68175
rect 210575 68147 210609 68175
rect 210637 68147 210671 68175
rect 210699 68147 219485 68175
rect 219513 68147 219547 68175
rect 219575 68147 219609 68175
rect 219637 68147 219671 68175
rect 219699 68147 228485 68175
rect 228513 68147 228547 68175
rect 228575 68147 228609 68175
rect 228637 68147 228671 68175
rect 228699 68147 237485 68175
rect 237513 68147 237547 68175
rect 237575 68147 237609 68175
rect 237637 68147 237671 68175
rect 237699 68147 246485 68175
rect 246513 68147 246547 68175
rect 246575 68147 246609 68175
rect 246637 68147 246671 68175
rect 246699 68147 255485 68175
rect 255513 68147 255547 68175
rect 255575 68147 255609 68175
rect 255637 68147 255671 68175
rect 255699 68147 264485 68175
rect 264513 68147 264547 68175
rect 264575 68147 264609 68175
rect 264637 68147 264671 68175
rect 264699 68147 273485 68175
rect 273513 68147 273547 68175
rect 273575 68147 273609 68175
rect 273637 68147 273671 68175
rect 273699 68147 282485 68175
rect 282513 68147 282547 68175
rect 282575 68147 282609 68175
rect 282637 68147 282671 68175
rect 282699 68147 291485 68175
rect 291513 68147 291547 68175
rect 291575 68147 291609 68175
rect 291637 68147 291671 68175
rect 291699 68147 298728 68175
rect 298756 68147 298790 68175
rect 298818 68147 298852 68175
rect 298880 68147 298914 68175
rect 298942 68147 298990 68175
rect -958 68113 298990 68147
rect -958 68085 -910 68113
rect -882 68085 -848 68113
rect -820 68085 -786 68113
rect -758 68085 -724 68113
rect -696 68085 3485 68113
rect 3513 68085 3547 68113
rect 3575 68085 3609 68113
rect 3637 68085 3671 68113
rect 3699 68085 12485 68113
rect 12513 68085 12547 68113
rect 12575 68085 12609 68113
rect 12637 68085 12671 68113
rect 12699 68085 21485 68113
rect 21513 68085 21547 68113
rect 21575 68085 21609 68113
rect 21637 68085 21671 68113
rect 21699 68085 30485 68113
rect 30513 68085 30547 68113
rect 30575 68085 30609 68113
rect 30637 68085 30671 68113
rect 30699 68085 39485 68113
rect 39513 68085 39547 68113
rect 39575 68085 39609 68113
rect 39637 68085 39671 68113
rect 39699 68085 48485 68113
rect 48513 68085 48547 68113
rect 48575 68085 48609 68113
rect 48637 68085 48671 68113
rect 48699 68085 54509 68113
rect 54537 68085 54571 68113
rect 54599 68085 57485 68113
rect 57513 68085 57547 68113
rect 57575 68085 57609 68113
rect 57637 68085 57671 68113
rect 57699 68085 59009 68113
rect 59037 68085 59071 68113
rect 59099 68085 63509 68113
rect 63537 68085 63571 68113
rect 63599 68085 66485 68113
rect 66513 68085 66547 68113
rect 66575 68085 66609 68113
rect 66637 68085 66671 68113
rect 66699 68085 68009 68113
rect 68037 68085 68071 68113
rect 68099 68085 72509 68113
rect 72537 68085 72571 68113
rect 72599 68085 75485 68113
rect 75513 68085 75547 68113
rect 75575 68085 75609 68113
rect 75637 68085 75671 68113
rect 75699 68085 77009 68113
rect 77037 68085 77071 68113
rect 77099 68085 81509 68113
rect 81537 68085 81571 68113
rect 81599 68085 84485 68113
rect 84513 68085 84547 68113
rect 84575 68085 84609 68113
rect 84637 68085 84671 68113
rect 84699 68085 86009 68113
rect 86037 68085 86071 68113
rect 86099 68085 90509 68113
rect 90537 68085 90571 68113
rect 90599 68085 95009 68113
rect 95037 68085 95071 68113
rect 95099 68085 99509 68113
rect 99537 68085 99571 68113
rect 99599 68085 104009 68113
rect 104037 68085 104071 68113
rect 104099 68085 108509 68113
rect 108537 68085 108571 68113
rect 108599 68085 113009 68113
rect 113037 68085 113071 68113
rect 113099 68085 117509 68113
rect 117537 68085 117571 68113
rect 117599 68085 120485 68113
rect 120513 68085 120547 68113
rect 120575 68085 120609 68113
rect 120637 68085 120671 68113
rect 120699 68085 129485 68113
rect 129513 68085 129547 68113
rect 129575 68085 129609 68113
rect 129637 68085 129671 68113
rect 129699 68085 138485 68113
rect 138513 68085 138547 68113
rect 138575 68085 138609 68113
rect 138637 68085 138671 68113
rect 138699 68085 147485 68113
rect 147513 68085 147547 68113
rect 147575 68085 147609 68113
rect 147637 68085 147671 68113
rect 147699 68085 156485 68113
rect 156513 68085 156547 68113
rect 156575 68085 156609 68113
rect 156637 68085 156671 68113
rect 156699 68085 165485 68113
rect 165513 68085 165547 68113
rect 165575 68085 165609 68113
rect 165637 68085 165671 68113
rect 165699 68085 174485 68113
rect 174513 68085 174547 68113
rect 174575 68085 174609 68113
rect 174637 68085 174671 68113
rect 174699 68085 183485 68113
rect 183513 68085 183547 68113
rect 183575 68085 183609 68113
rect 183637 68085 183671 68113
rect 183699 68085 192485 68113
rect 192513 68085 192547 68113
rect 192575 68085 192609 68113
rect 192637 68085 192671 68113
rect 192699 68085 201485 68113
rect 201513 68085 201547 68113
rect 201575 68085 201609 68113
rect 201637 68085 201671 68113
rect 201699 68085 210485 68113
rect 210513 68085 210547 68113
rect 210575 68085 210609 68113
rect 210637 68085 210671 68113
rect 210699 68085 219485 68113
rect 219513 68085 219547 68113
rect 219575 68085 219609 68113
rect 219637 68085 219671 68113
rect 219699 68085 228485 68113
rect 228513 68085 228547 68113
rect 228575 68085 228609 68113
rect 228637 68085 228671 68113
rect 228699 68085 237485 68113
rect 237513 68085 237547 68113
rect 237575 68085 237609 68113
rect 237637 68085 237671 68113
rect 237699 68085 246485 68113
rect 246513 68085 246547 68113
rect 246575 68085 246609 68113
rect 246637 68085 246671 68113
rect 246699 68085 255485 68113
rect 255513 68085 255547 68113
rect 255575 68085 255609 68113
rect 255637 68085 255671 68113
rect 255699 68085 264485 68113
rect 264513 68085 264547 68113
rect 264575 68085 264609 68113
rect 264637 68085 264671 68113
rect 264699 68085 273485 68113
rect 273513 68085 273547 68113
rect 273575 68085 273609 68113
rect 273637 68085 273671 68113
rect 273699 68085 282485 68113
rect 282513 68085 282547 68113
rect 282575 68085 282609 68113
rect 282637 68085 282671 68113
rect 282699 68085 291485 68113
rect 291513 68085 291547 68113
rect 291575 68085 291609 68113
rect 291637 68085 291671 68113
rect 291699 68085 298728 68113
rect 298756 68085 298790 68113
rect 298818 68085 298852 68113
rect 298880 68085 298914 68113
rect 298942 68085 298990 68113
rect -958 68051 298990 68085
rect -958 68023 -910 68051
rect -882 68023 -848 68051
rect -820 68023 -786 68051
rect -758 68023 -724 68051
rect -696 68023 3485 68051
rect 3513 68023 3547 68051
rect 3575 68023 3609 68051
rect 3637 68023 3671 68051
rect 3699 68023 12485 68051
rect 12513 68023 12547 68051
rect 12575 68023 12609 68051
rect 12637 68023 12671 68051
rect 12699 68023 21485 68051
rect 21513 68023 21547 68051
rect 21575 68023 21609 68051
rect 21637 68023 21671 68051
rect 21699 68023 30485 68051
rect 30513 68023 30547 68051
rect 30575 68023 30609 68051
rect 30637 68023 30671 68051
rect 30699 68023 39485 68051
rect 39513 68023 39547 68051
rect 39575 68023 39609 68051
rect 39637 68023 39671 68051
rect 39699 68023 48485 68051
rect 48513 68023 48547 68051
rect 48575 68023 48609 68051
rect 48637 68023 48671 68051
rect 48699 68023 54509 68051
rect 54537 68023 54571 68051
rect 54599 68023 57485 68051
rect 57513 68023 57547 68051
rect 57575 68023 57609 68051
rect 57637 68023 57671 68051
rect 57699 68023 59009 68051
rect 59037 68023 59071 68051
rect 59099 68023 63509 68051
rect 63537 68023 63571 68051
rect 63599 68023 66485 68051
rect 66513 68023 66547 68051
rect 66575 68023 66609 68051
rect 66637 68023 66671 68051
rect 66699 68023 68009 68051
rect 68037 68023 68071 68051
rect 68099 68023 72509 68051
rect 72537 68023 72571 68051
rect 72599 68023 75485 68051
rect 75513 68023 75547 68051
rect 75575 68023 75609 68051
rect 75637 68023 75671 68051
rect 75699 68023 77009 68051
rect 77037 68023 77071 68051
rect 77099 68023 81509 68051
rect 81537 68023 81571 68051
rect 81599 68023 84485 68051
rect 84513 68023 84547 68051
rect 84575 68023 84609 68051
rect 84637 68023 84671 68051
rect 84699 68023 86009 68051
rect 86037 68023 86071 68051
rect 86099 68023 90509 68051
rect 90537 68023 90571 68051
rect 90599 68023 95009 68051
rect 95037 68023 95071 68051
rect 95099 68023 99509 68051
rect 99537 68023 99571 68051
rect 99599 68023 104009 68051
rect 104037 68023 104071 68051
rect 104099 68023 108509 68051
rect 108537 68023 108571 68051
rect 108599 68023 113009 68051
rect 113037 68023 113071 68051
rect 113099 68023 117509 68051
rect 117537 68023 117571 68051
rect 117599 68023 120485 68051
rect 120513 68023 120547 68051
rect 120575 68023 120609 68051
rect 120637 68023 120671 68051
rect 120699 68023 129485 68051
rect 129513 68023 129547 68051
rect 129575 68023 129609 68051
rect 129637 68023 129671 68051
rect 129699 68023 138485 68051
rect 138513 68023 138547 68051
rect 138575 68023 138609 68051
rect 138637 68023 138671 68051
rect 138699 68023 147485 68051
rect 147513 68023 147547 68051
rect 147575 68023 147609 68051
rect 147637 68023 147671 68051
rect 147699 68023 156485 68051
rect 156513 68023 156547 68051
rect 156575 68023 156609 68051
rect 156637 68023 156671 68051
rect 156699 68023 165485 68051
rect 165513 68023 165547 68051
rect 165575 68023 165609 68051
rect 165637 68023 165671 68051
rect 165699 68023 174485 68051
rect 174513 68023 174547 68051
rect 174575 68023 174609 68051
rect 174637 68023 174671 68051
rect 174699 68023 183485 68051
rect 183513 68023 183547 68051
rect 183575 68023 183609 68051
rect 183637 68023 183671 68051
rect 183699 68023 192485 68051
rect 192513 68023 192547 68051
rect 192575 68023 192609 68051
rect 192637 68023 192671 68051
rect 192699 68023 201485 68051
rect 201513 68023 201547 68051
rect 201575 68023 201609 68051
rect 201637 68023 201671 68051
rect 201699 68023 210485 68051
rect 210513 68023 210547 68051
rect 210575 68023 210609 68051
rect 210637 68023 210671 68051
rect 210699 68023 219485 68051
rect 219513 68023 219547 68051
rect 219575 68023 219609 68051
rect 219637 68023 219671 68051
rect 219699 68023 228485 68051
rect 228513 68023 228547 68051
rect 228575 68023 228609 68051
rect 228637 68023 228671 68051
rect 228699 68023 237485 68051
rect 237513 68023 237547 68051
rect 237575 68023 237609 68051
rect 237637 68023 237671 68051
rect 237699 68023 246485 68051
rect 246513 68023 246547 68051
rect 246575 68023 246609 68051
rect 246637 68023 246671 68051
rect 246699 68023 255485 68051
rect 255513 68023 255547 68051
rect 255575 68023 255609 68051
rect 255637 68023 255671 68051
rect 255699 68023 264485 68051
rect 264513 68023 264547 68051
rect 264575 68023 264609 68051
rect 264637 68023 264671 68051
rect 264699 68023 273485 68051
rect 273513 68023 273547 68051
rect 273575 68023 273609 68051
rect 273637 68023 273671 68051
rect 273699 68023 282485 68051
rect 282513 68023 282547 68051
rect 282575 68023 282609 68051
rect 282637 68023 282671 68051
rect 282699 68023 291485 68051
rect 291513 68023 291547 68051
rect 291575 68023 291609 68051
rect 291637 68023 291671 68051
rect 291699 68023 298728 68051
rect 298756 68023 298790 68051
rect 298818 68023 298852 68051
rect 298880 68023 298914 68051
rect 298942 68023 298990 68051
rect -958 67989 298990 68023
rect -958 67961 -910 67989
rect -882 67961 -848 67989
rect -820 67961 -786 67989
rect -758 67961 -724 67989
rect -696 67961 3485 67989
rect 3513 67961 3547 67989
rect 3575 67961 3609 67989
rect 3637 67961 3671 67989
rect 3699 67961 12485 67989
rect 12513 67961 12547 67989
rect 12575 67961 12609 67989
rect 12637 67961 12671 67989
rect 12699 67961 21485 67989
rect 21513 67961 21547 67989
rect 21575 67961 21609 67989
rect 21637 67961 21671 67989
rect 21699 67961 30485 67989
rect 30513 67961 30547 67989
rect 30575 67961 30609 67989
rect 30637 67961 30671 67989
rect 30699 67961 39485 67989
rect 39513 67961 39547 67989
rect 39575 67961 39609 67989
rect 39637 67961 39671 67989
rect 39699 67961 48485 67989
rect 48513 67961 48547 67989
rect 48575 67961 48609 67989
rect 48637 67961 48671 67989
rect 48699 67961 54509 67989
rect 54537 67961 54571 67989
rect 54599 67961 57485 67989
rect 57513 67961 57547 67989
rect 57575 67961 57609 67989
rect 57637 67961 57671 67989
rect 57699 67961 59009 67989
rect 59037 67961 59071 67989
rect 59099 67961 63509 67989
rect 63537 67961 63571 67989
rect 63599 67961 66485 67989
rect 66513 67961 66547 67989
rect 66575 67961 66609 67989
rect 66637 67961 66671 67989
rect 66699 67961 68009 67989
rect 68037 67961 68071 67989
rect 68099 67961 72509 67989
rect 72537 67961 72571 67989
rect 72599 67961 75485 67989
rect 75513 67961 75547 67989
rect 75575 67961 75609 67989
rect 75637 67961 75671 67989
rect 75699 67961 77009 67989
rect 77037 67961 77071 67989
rect 77099 67961 81509 67989
rect 81537 67961 81571 67989
rect 81599 67961 84485 67989
rect 84513 67961 84547 67989
rect 84575 67961 84609 67989
rect 84637 67961 84671 67989
rect 84699 67961 86009 67989
rect 86037 67961 86071 67989
rect 86099 67961 90509 67989
rect 90537 67961 90571 67989
rect 90599 67961 95009 67989
rect 95037 67961 95071 67989
rect 95099 67961 99509 67989
rect 99537 67961 99571 67989
rect 99599 67961 104009 67989
rect 104037 67961 104071 67989
rect 104099 67961 108509 67989
rect 108537 67961 108571 67989
rect 108599 67961 113009 67989
rect 113037 67961 113071 67989
rect 113099 67961 117509 67989
rect 117537 67961 117571 67989
rect 117599 67961 120485 67989
rect 120513 67961 120547 67989
rect 120575 67961 120609 67989
rect 120637 67961 120671 67989
rect 120699 67961 129485 67989
rect 129513 67961 129547 67989
rect 129575 67961 129609 67989
rect 129637 67961 129671 67989
rect 129699 67961 138485 67989
rect 138513 67961 138547 67989
rect 138575 67961 138609 67989
rect 138637 67961 138671 67989
rect 138699 67961 147485 67989
rect 147513 67961 147547 67989
rect 147575 67961 147609 67989
rect 147637 67961 147671 67989
rect 147699 67961 156485 67989
rect 156513 67961 156547 67989
rect 156575 67961 156609 67989
rect 156637 67961 156671 67989
rect 156699 67961 165485 67989
rect 165513 67961 165547 67989
rect 165575 67961 165609 67989
rect 165637 67961 165671 67989
rect 165699 67961 174485 67989
rect 174513 67961 174547 67989
rect 174575 67961 174609 67989
rect 174637 67961 174671 67989
rect 174699 67961 183485 67989
rect 183513 67961 183547 67989
rect 183575 67961 183609 67989
rect 183637 67961 183671 67989
rect 183699 67961 192485 67989
rect 192513 67961 192547 67989
rect 192575 67961 192609 67989
rect 192637 67961 192671 67989
rect 192699 67961 201485 67989
rect 201513 67961 201547 67989
rect 201575 67961 201609 67989
rect 201637 67961 201671 67989
rect 201699 67961 210485 67989
rect 210513 67961 210547 67989
rect 210575 67961 210609 67989
rect 210637 67961 210671 67989
rect 210699 67961 219485 67989
rect 219513 67961 219547 67989
rect 219575 67961 219609 67989
rect 219637 67961 219671 67989
rect 219699 67961 228485 67989
rect 228513 67961 228547 67989
rect 228575 67961 228609 67989
rect 228637 67961 228671 67989
rect 228699 67961 237485 67989
rect 237513 67961 237547 67989
rect 237575 67961 237609 67989
rect 237637 67961 237671 67989
rect 237699 67961 246485 67989
rect 246513 67961 246547 67989
rect 246575 67961 246609 67989
rect 246637 67961 246671 67989
rect 246699 67961 255485 67989
rect 255513 67961 255547 67989
rect 255575 67961 255609 67989
rect 255637 67961 255671 67989
rect 255699 67961 264485 67989
rect 264513 67961 264547 67989
rect 264575 67961 264609 67989
rect 264637 67961 264671 67989
rect 264699 67961 273485 67989
rect 273513 67961 273547 67989
rect 273575 67961 273609 67989
rect 273637 67961 273671 67989
rect 273699 67961 282485 67989
rect 282513 67961 282547 67989
rect 282575 67961 282609 67989
rect 282637 67961 282671 67989
rect 282699 67961 291485 67989
rect 291513 67961 291547 67989
rect 291575 67961 291609 67989
rect 291637 67961 291671 67989
rect 291699 67961 298728 67989
rect 298756 67961 298790 67989
rect 298818 67961 298852 67989
rect 298880 67961 298914 67989
rect 298942 67961 298990 67989
rect -958 67913 298990 67961
rect -958 65175 298990 65223
rect -958 65147 -430 65175
rect -402 65147 -368 65175
rect -340 65147 -306 65175
rect -278 65147 -244 65175
rect -216 65147 1625 65175
rect 1653 65147 1687 65175
rect 1715 65147 1749 65175
rect 1777 65147 1811 65175
rect 1839 65147 10625 65175
rect 10653 65147 10687 65175
rect 10715 65147 10749 65175
rect 10777 65147 10811 65175
rect 10839 65147 19625 65175
rect 19653 65147 19687 65175
rect 19715 65147 19749 65175
rect 19777 65147 19811 65175
rect 19839 65147 28625 65175
rect 28653 65147 28687 65175
rect 28715 65147 28749 65175
rect 28777 65147 28811 65175
rect 28839 65147 37625 65175
rect 37653 65147 37687 65175
rect 37715 65147 37749 65175
rect 37777 65147 37811 65175
rect 37839 65147 46625 65175
rect 46653 65147 46687 65175
rect 46715 65147 46749 65175
rect 46777 65147 46811 65175
rect 46839 65147 52259 65175
rect 52287 65147 52321 65175
rect 52349 65147 55625 65175
rect 55653 65147 55687 65175
rect 55715 65147 55749 65175
rect 55777 65147 55811 65175
rect 55839 65147 56759 65175
rect 56787 65147 56821 65175
rect 56849 65147 61259 65175
rect 61287 65147 61321 65175
rect 61349 65147 64625 65175
rect 64653 65147 64687 65175
rect 64715 65147 64749 65175
rect 64777 65147 64811 65175
rect 64839 65147 65759 65175
rect 65787 65147 65821 65175
rect 65849 65147 70259 65175
rect 70287 65147 70321 65175
rect 70349 65147 73625 65175
rect 73653 65147 73687 65175
rect 73715 65147 73749 65175
rect 73777 65147 73811 65175
rect 73839 65147 74759 65175
rect 74787 65147 74821 65175
rect 74849 65147 79259 65175
rect 79287 65147 79321 65175
rect 79349 65147 82625 65175
rect 82653 65147 82687 65175
rect 82715 65147 82749 65175
rect 82777 65147 82811 65175
rect 82839 65147 83759 65175
rect 83787 65147 83821 65175
rect 83849 65147 88259 65175
rect 88287 65147 88321 65175
rect 88349 65147 91625 65175
rect 91653 65147 91687 65175
rect 91715 65147 91749 65175
rect 91777 65147 91811 65175
rect 91839 65147 92759 65175
rect 92787 65147 92821 65175
rect 92849 65147 97259 65175
rect 97287 65147 97321 65175
rect 97349 65147 101759 65175
rect 101787 65147 101821 65175
rect 101849 65147 106259 65175
rect 106287 65147 106321 65175
rect 106349 65147 110759 65175
rect 110787 65147 110821 65175
rect 110849 65147 115259 65175
rect 115287 65147 115321 65175
rect 115349 65147 127625 65175
rect 127653 65147 127687 65175
rect 127715 65147 127749 65175
rect 127777 65147 127811 65175
rect 127839 65147 136625 65175
rect 136653 65147 136687 65175
rect 136715 65147 136749 65175
rect 136777 65147 136811 65175
rect 136839 65147 145625 65175
rect 145653 65147 145687 65175
rect 145715 65147 145749 65175
rect 145777 65147 145811 65175
rect 145839 65147 154625 65175
rect 154653 65147 154687 65175
rect 154715 65147 154749 65175
rect 154777 65147 154811 65175
rect 154839 65147 163625 65175
rect 163653 65147 163687 65175
rect 163715 65147 163749 65175
rect 163777 65147 163811 65175
rect 163839 65147 172625 65175
rect 172653 65147 172687 65175
rect 172715 65147 172749 65175
rect 172777 65147 172811 65175
rect 172839 65147 181625 65175
rect 181653 65147 181687 65175
rect 181715 65147 181749 65175
rect 181777 65147 181811 65175
rect 181839 65147 190625 65175
rect 190653 65147 190687 65175
rect 190715 65147 190749 65175
rect 190777 65147 190811 65175
rect 190839 65147 199625 65175
rect 199653 65147 199687 65175
rect 199715 65147 199749 65175
rect 199777 65147 199811 65175
rect 199839 65147 208625 65175
rect 208653 65147 208687 65175
rect 208715 65147 208749 65175
rect 208777 65147 208811 65175
rect 208839 65147 217625 65175
rect 217653 65147 217687 65175
rect 217715 65147 217749 65175
rect 217777 65147 217811 65175
rect 217839 65147 226625 65175
rect 226653 65147 226687 65175
rect 226715 65147 226749 65175
rect 226777 65147 226811 65175
rect 226839 65147 235625 65175
rect 235653 65147 235687 65175
rect 235715 65147 235749 65175
rect 235777 65147 235811 65175
rect 235839 65147 244625 65175
rect 244653 65147 244687 65175
rect 244715 65147 244749 65175
rect 244777 65147 244811 65175
rect 244839 65147 253625 65175
rect 253653 65147 253687 65175
rect 253715 65147 253749 65175
rect 253777 65147 253811 65175
rect 253839 65147 262625 65175
rect 262653 65147 262687 65175
rect 262715 65147 262749 65175
rect 262777 65147 262811 65175
rect 262839 65147 271625 65175
rect 271653 65147 271687 65175
rect 271715 65147 271749 65175
rect 271777 65147 271811 65175
rect 271839 65147 280625 65175
rect 280653 65147 280687 65175
rect 280715 65147 280749 65175
rect 280777 65147 280811 65175
rect 280839 65147 289625 65175
rect 289653 65147 289687 65175
rect 289715 65147 289749 65175
rect 289777 65147 289811 65175
rect 289839 65147 298248 65175
rect 298276 65147 298310 65175
rect 298338 65147 298372 65175
rect 298400 65147 298434 65175
rect 298462 65147 298990 65175
rect -958 65113 298990 65147
rect -958 65085 -430 65113
rect -402 65085 -368 65113
rect -340 65085 -306 65113
rect -278 65085 -244 65113
rect -216 65085 1625 65113
rect 1653 65085 1687 65113
rect 1715 65085 1749 65113
rect 1777 65085 1811 65113
rect 1839 65085 10625 65113
rect 10653 65085 10687 65113
rect 10715 65085 10749 65113
rect 10777 65085 10811 65113
rect 10839 65085 19625 65113
rect 19653 65085 19687 65113
rect 19715 65085 19749 65113
rect 19777 65085 19811 65113
rect 19839 65085 28625 65113
rect 28653 65085 28687 65113
rect 28715 65085 28749 65113
rect 28777 65085 28811 65113
rect 28839 65085 37625 65113
rect 37653 65085 37687 65113
rect 37715 65085 37749 65113
rect 37777 65085 37811 65113
rect 37839 65085 46625 65113
rect 46653 65085 46687 65113
rect 46715 65085 46749 65113
rect 46777 65085 46811 65113
rect 46839 65085 52259 65113
rect 52287 65085 52321 65113
rect 52349 65085 55625 65113
rect 55653 65085 55687 65113
rect 55715 65085 55749 65113
rect 55777 65085 55811 65113
rect 55839 65085 56759 65113
rect 56787 65085 56821 65113
rect 56849 65085 61259 65113
rect 61287 65085 61321 65113
rect 61349 65085 64625 65113
rect 64653 65085 64687 65113
rect 64715 65085 64749 65113
rect 64777 65085 64811 65113
rect 64839 65085 65759 65113
rect 65787 65085 65821 65113
rect 65849 65085 70259 65113
rect 70287 65085 70321 65113
rect 70349 65085 73625 65113
rect 73653 65085 73687 65113
rect 73715 65085 73749 65113
rect 73777 65085 73811 65113
rect 73839 65085 74759 65113
rect 74787 65085 74821 65113
rect 74849 65085 79259 65113
rect 79287 65085 79321 65113
rect 79349 65085 82625 65113
rect 82653 65085 82687 65113
rect 82715 65085 82749 65113
rect 82777 65085 82811 65113
rect 82839 65085 83759 65113
rect 83787 65085 83821 65113
rect 83849 65085 88259 65113
rect 88287 65085 88321 65113
rect 88349 65085 91625 65113
rect 91653 65085 91687 65113
rect 91715 65085 91749 65113
rect 91777 65085 91811 65113
rect 91839 65085 92759 65113
rect 92787 65085 92821 65113
rect 92849 65085 97259 65113
rect 97287 65085 97321 65113
rect 97349 65085 101759 65113
rect 101787 65085 101821 65113
rect 101849 65085 106259 65113
rect 106287 65085 106321 65113
rect 106349 65085 110759 65113
rect 110787 65085 110821 65113
rect 110849 65085 115259 65113
rect 115287 65085 115321 65113
rect 115349 65085 127625 65113
rect 127653 65085 127687 65113
rect 127715 65085 127749 65113
rect 127777 65085 127811 65113
rect 127839 65085 136625 65113
rect 136653 65085 136687 65113
rect 136715 65085 136749 65113
rect 136777 65085 136811 65113
rect 136839 65085 145625 65113
rect 145653 65085 145687 65113
rect 145715 65085 145749 65113
rect 145777 65085 145811 65113
rect 145839 65085 154625 65113
rect 154653 65085 154687 65113
rect 154715 65085 154749 65113
rect 154777 65085 154811 65113
rect 154839 65085 163625 65113
rect 163653 65085 163687 65113
rect 163715 65085 163749 65113
rect 163777 65085 163811 65113
rect 163839 65085 172625 65113
rect 172653 65085 172687 65113
rect 172715 65085 172749 65113
rect 172777 65085 172811 65113
rect 172839 65085 181625 65113
rect 181653 65085 181687 65113
rect 181715 65085 181749 65113
rect 181777 65085 181811 65113
rect 181839 65085 190625 65113
rect 190653 65085 190687 65113
rect 190715 65085 190749 65113
rect 190777 65085 190811 65113
rect 190839 65085 199625 65113
rect 199653 65085 199687 65113
rect 199715 65085 199749 65113
rect 199777 65085 199811 65113
rect 199839 65085 208625 65113
rect 208653 65085 208687 65113
rect 208715 65085 208749 65113
rect 208777 65085 208811 65113
rect 208839 65085 217625 65113
rect 217653 65085 217687 65113
rect 217715 65085 217749 65113
rect 217777 65085 217811 65113
rect 217839 65085 226625 65113
rect 226653 65085 226687 65113
rect 226715 65085 226749 65113
rect 226777 65085 226811 65113
rect 226839 65085 235625 65113
rect 235653 65085 235687 65113
rect 235715 65085 235749 65113
rect 235777 65085 235811 65113
rect 235839 65085 244625 65113
rect 244653 65085 244687 65113
rect 244715 65085 244749 65113
rect 244777 65085 244811 65113
rect 244839 65085 253625 65113
rect 253653 65085 253687 65113
rect 253715 65085 253749 65113
rect 253777 65085 253811 65113
rect 253839 65085 262625 65113
rect 262653 65085 262687 65113
rect 262715 65085 262749 65113
rect 262777 65085 262811 65113
rect 262839 65085 271625 65113
rect 271653 65085 271687 65113
rect 271715 65085 271749 65113
rect 271777 65085 271811 65113
rect 271839 65085 280625 65113
rect 280653 65085 280687 65113
rect 280715 65085 280749 65113
rect 280777 65085 280811 65113
rect 280839 65085 289625 65113
rect 289653 65085 289687 65113
rect 289715 65085 289749 65113
rect 289777 65085 289811 65113
rect 289839 65085 298248 65113
rect 298276 65085 298310 65113
rect 298338 65085 298372 65113
rect 298400 65085 298434 65113
rect 298462 65085 298990 65113
rect -958 65051 298990 65085
rect -958 65023 -430 65051
rect -402 65023 -368 65051
rect -340 65023 -306 65051
rect -278 65023 -244 65051
rect -216 65023 1625 65051
rect 1653 65023 1687 65051
rect 1715 65023 1749 65051
rect 1777 65023 1811 65051
rect 1839 65023 10625 65051
rect 10653 65023 10687 65051
rect 10715 65023 10749 65051
rect 10777 65023 10811 65051
rect 10839 65023 19625 65051
rect 19653 65023 19687 65051
rect 19715 65023 19749 65051
rect 19777 65023 19811 65051
rect 19839 65023 28625 65051
rect 28653 65023 28687 65051
rect 28715 65023 28749 65051
rect 28777 65023 28811 65051
rect 28839 65023 37625 65051
rect 37653 65023 37687 65051
rect 37715 65023 37749 65051
rect 37777 65023 37811 65051
rect 37839 65023 46625 65051
rect 46653 65023 46687 65051
rect 46715 65023 46749 65051
rect 46777 65023 46811 65051
rect 46839 65023 52259 65051
rect 52287 65023 52321 65051
rect 52349 65023 55625 65051
rect 55653 65023 55687 65051
rect 55715 65023 55749 65051
rect 55777 65023 55811 65051
rect 55839 65023 56759 65051
rect 56787 65023 56821 65051
rect 56849 65023 61259 65051
rect 61287 65023 61321 65051
rect 61349 65023 64625 65051
rect 64653 65023 64687 65051
rect 64715 65023 64749 65051
rect 64777 65023 64811 65051
rect 64839 65023 65759 65051
rect 65787 65023 65821 65051
rect 65849 65023 70259 65051
rect 70287 65023 70321 65051
rect 70349 65023 73625 65051
rect 73653 65023 73687 65051
rect 73715 65023 73749 65051
rect 73777 65023 73811 65051
rect 73839 65023 74759 65051
rect 74787 65023 74821 65051
rect 74849 65023 79259 65051
rect 79287 65023 79321 65051
rect 79349 65023 82625 65051
rect 82653 65023 82687 65051
rect 82715 65023 82749 65051
rect 82777 65023 82811 65051
rect 82839 65023 83759 65051
rect 83787 65023 83821 65051
rect 83849 65023 88259 65051
rect 88287 65023 88321 65051
rect 88349 65023 91625 65051
rect 91653 65023 91687 65051
rect 91715 65023 91749 65051
rect 91777 65023 91811 65051
rect 91839 65023 92759 65051
rect 92787 65023 92821 65051
rect 92849 65023 97259 65051
rect 97287 65023 97321 65051
rect 97349 65023 101759 65051
rect 101787 65023 101821 65051
rect 101849 65023 106259 65051
rect 106287 65023 106321 65051
rect 106349 65023 110759 65051
rect 110787 65023 110821 65051
rect 110849 65023 115259 65051
rect 115287 65023 115321 65051
rect 115349 65023 127625 65051
rect 127653 65023 127687 65051
rect 127715 65023 127749 65051
rect 127777 65023 127811 65051
rect 127839 65023 136625 65051
rect 136653 65023 136687 65051
rect 136715 65023 136749 65051
rect 136777 65023 136811 65051
rect 136839 65023 145625 65051
rect 145653 65023 145687 65051
rect 145715 65023 145749 65051
rect 145777 65023 145811 65051
rect 145839 65023 154625 65051
rect 154653 65023 154687 65051
rect 154715 65023 154749 65051
rect 154777 65023 154811 65051
rect 154839 65023 163625 65051
rect 163653 65023 163687 65051
rect 163715 65023 163749 65051
rect 163777 65023 163811 65051
rect 163839 65023 172625 65051
rect 172653 65023 172687 65051
rect 172715 65023 172749 65051
rect 172777 65023 172811 65051
rect 172839 65023 181625 65051
rect 181653 65023 181687 65051
rect 181715 65023 181749 65051
rect 181777 65023 181811 65051
rect 181839 65023 190625 65051
rect 190653 65023 190687 65051
rect 190715 65023 190749 65051
rect 190777 65023 190811 65051
rect 190839 65023 199625 65051
rect 199653 65023 199687 65051
rect 199715 65023 199749 65051
rect 199777 65023 199811 65051
rect 199839 65023 208625 65051
rect 208653 65023 208687 65051
rect 208715 65023 208749 65051
rect 208777 65023 208811 65051
rect 208839 65023 217625 65051
rect 217653 65023 217687 65051
rect 217715 65023 217749 65051
rect 217777 65023 217811 65051
rect 217839 65023 226625 65051
rect 226653 65023 226687 65051
rect 226715 65023 226749 65051
rect 226777 65023 226811 65051
rect 226839 65023 235625 65051
rect 235653 65023 235687 65051
rect 235715 65023 235749 65051
rect 235777 65023 235811 65051
rect 235839 65023 244625 65051
rect 244653 65023 244687 65051
rect 244715 65023 244749 65051
rect 244777 65023 244811 65051
rect 244839 65023 253625 65051
rect 253653 65023 253687 65051
rect 253715 65023 253749 65051
rect 253777 65023 253811 65051
rect 253839 65023 262625 65051
rect 262653 65023 262687 65051
rect 262715 65023 262749 65051
rect 262777 65023 262811 65051
rect 262839 65023 271625 65051
rect 271653 65023 271687 65051
rect 271715 65023 271749 65051
rect 271777 65023 271811 65051
rect 271839 65023 280625 65051
rect 280653 65023 280687 65051
rect 280715 65023 280749 65051
rect 280777 65023 280811 65051
rect 280839 65023 289625 65051
rect 289653 65023 289687 65051
rect 289715 65023 289749 65051
rect 289777 65023 289811 65051
rect 289839 65023 298248 65051
rect 298276 65023 298310 65051
rect 298338 65023 298372 65051
rect 298400 65023 298434 65051
rect 298462 65023 298990 65051
rect -958 64989 298990 65023
rect -958 64961 -430 64989
rect -402 64961 -368 64989
rect -340 64961 -306 64989
rect -278 64961 -244 64989
rect -216 64961 1625 64989
rect 1653 64961 1687 64989
rect 1715 64961 1749 64989
rect 1777 64961 1811 64989
rect 1839 64961 10625 64989
rect 10653 64961 10687 64989
rect 10715 64961 10749 64989
rect 10777 64961 10811 64989
rect 10839 64961 19625 64989
rect 19653 64961 19687 64989
rect 19715 64961 19749 64989
rect 19777 64961 19811 64989
rect 19839 64961 28625 64989
rect 28653 64961 28687 64989
rect 28715 64961 28749 64989
rect 28777 64961 28811 64989
rect 28839 64961 37625 64989
rect 37653 64961 37687 64989
rect 37715 64961 37749 64989
rect 37777 64961 37811 64989
rect 37839 64961 46625 64989
rect 46653 64961 46687 64989
rect 46715 64961 46749 64989
rect 46777 64961 46811 64989
rect 46839 64961 52259 64989
rect 52287 64961 52321 64989
rect 52349 64961 55625 64989
rect 55653 64961 55687 64989
rect 55715 64961 55749 64989
rect 55777 64961 55811 64989
rect 55839 64961 56759 64989
rect 56787 64961 56821 64989
rect 56849 64961 61259 64989
rect 61287 64961 61321 64989
rect 61349 64961 64625 64989
rect 64653 64961 64687 64989
rect 64715 64961 64749 64989
rect 64777 64961 64811 64989
rect 64839 64961 65759 64989
rect 65787 64961 65821 64989
rect 65849 64961 70259 64989
rect 70287 64961 70321 64989
rect 70349 64961 73625 64989
rect 73653 64961 73687 64989
rect 73715 64961 73749 64989
rect 73777 64961 73811 64989
rect 73839 64961 74759 64989
rect 74787 64961 74821 64989
rect 74849 64961 79259 64989
rect 79287 64961 79321 64989
rect 79349 64961 82625 64989
rect 82653 64961 82687 64989
rect 82715 64961 82749 64989
rect 82777 64961 82811 64989
rect 82839 64961 83759 64989
rect 83787 64961 83821 64989
rect 83849 64961 88259 64989
rect 88287 64961 88321 64989
rect 88349 64961 91625 64989
rect 91653 64961 91687 64989
rect 91715 64961 91749 64989
rect 91777 64961 91811 64989
rect 91839 64961 92759 64989
rect 92787 64961 92821 64989
rect 92849 64961 97259 64989
rect 97287 64961 97321 64989
rect 97349 64961 101759 64989
rect 101787 64961 101821 64989
rect 101849 64961 106259 64989
rect 106287 64961 106321 64989
rect 106349 64961 110759 64989
rect 110787 64961 110821 64989
rect 110849 64961 115259 64989
rect 115287 64961 115321 64989
rect 115349 64961 127625 64989
rect 127653 64961 127687 64989
rect 127715 64961 127749 64989
rect 127777 64961 127811 64989
rect 127839 64961 136625 64989
rect 136653 64961 136687 64989
rect 136715 64961 136749 64989
rect 136777 64961 136811 64989
rect 136839 64961 145625 64989
rect 145653 64961 145687 64989
rect 145715 64961 145749 64989
rect 145777 64961 145811 64989
rect 145839 64961 154625 64989
rect 154653 64961 154687 64989
rect 154715 64961 154749 64989
rect 154777 64961 154811 64989
rect 154839 64961 163625 64989
rect 163653 64961 163687 64989
rect 163715 64961 163749 64989
rect 163777 64961 163811 64989
rect 163839 64961 172625 64989
rect 172653 64961 172687 64989
rect 172715 64961 172749 64989
rect 172777 64961 172811 64989
rect 172839 64961 181625 64989
rect 181653 64961 181687 64989
rect 181715 64961 181749 64989
rect 181777 64961 181811 64989
rect 181839 64961 190625 64989
rect 190653 64961 190687 64989
rect 190715 64961 190749 64989
rect 190777 64961 190811 64989
rect 190839 64961 199625 64989
rect 199653 64961 199687 64989
rect 199715 64961 199749 64989
rect 199777 64961 199811 64989
rect 199839 64961 208625 64989
rect 208653 64961 208687 64989
rect 208715 64961 208749 64989
rect 208777 64961 208811 64989
rect 208839 64961 217625 64989
rect 217653 64961 217687 64989
rect 217715 64961 217749 64989
rect 217777 64961 217811 64989
rect 217839 64961 226625 64989
rect 226653 64961 226687 64989
rect 226715 64961 226749 64989
rect 226777 64961 226811 64989
rect 226839 64961 235625 64989
rect 235653 64961 235687 64989
rect 235715 64961 235749 64989
rect 235777 64961 235811 64989
rect 235839 64961 244625 64989
rect 244653 64961 244687 64989
rect 244715 64961 244749 64989
rect 244777 64961 244811 64989
rect 244839 64961 253625 64989
rect 253653 64961 253687 64989
rect 253715 64961 253749 64989
rect 253777 64961 253811 64989
rect 253839 64961 262625 64989
rect 262653 64961 262687 64989
rect 262715 64961 262749 64989
rect 262777 64961 262811 64989
rect 262839 64961 271625 64989
rect 271653 64961 271687 64989
rect 271715 64961 271749 64989
rect 271777 64961 271811 64989
rect 271839 64961 280625 64989
rect 280653 64961 280687 64989
rect 280715 64961 280749 64989
rect 280777 64961 280811 64989
rect 280839 64961 289625 64989
rect 289653 64961 289687 64989
rect 289715 64961 289749 64989
rect 289777 64961 289811 64989
rect 289839 64961 298248 64989
rect 298276 64961 298310 64989
rect 298338 64961 298372 64989
rect 298400 64961 298434 64989
rect 298462 64961 298990 64989
rect -958 64913 298990 64961
rect -958 59175 298990 59223
rect -958 59147 -910 59175
rect -882 59147 -848 59175
rect -820 59147 -786 59175
rect -758 59147 -724 59175
rect -696 59147 3485 59175
rect 3513 59147 3547 59175
rect 3575 59147 3609 59175
rect 3637 59147 3671 59175
rect 3699 59147 12485 59175
rect 12513 59147 12547 59175
rect 12575 59147 12609 59175
rect 12637 59147 12671 59175
rect 12699 59147 21485 59175
rect 21513 59147 21547 59175
rect 21575 59147 21609 59175
rect 21637 59147 21671 59175
rect 21699 59147 30485 59175
rect 30513 59147 30547 59175
rect 30575 59147 30609 59175
rect 30637 59147 30671 59175
rect 30699 59147 39485 59175
rect 39513 59147 39547 59175
rect 39575 59147 39609 59175
rect 39637 59147 39671 59175
rect 39699 59147 48485 59175
rect 48513 59147 48547 59175
rect 48575 59147 48609 59175
rect 48637 59147 48671 59175
rect 48699 59147 54509 59175
rect 54537 59147 54571 59175
rect 54599 59147 57485 59175
rect 57513 59147 57547 59175
rect 57575 59147 57609 59175
rect 57637 59147 57671 59175
rect 57699 59147 59009 59175
rect 59037 59147 59071 59175
rect 59099 59147 63509 59175
rect 63537 59147 63571 59175
rect 63599 59147 66485 59175
rect 66513 59147 66547 59175
rect 66575 59147 66609 59175
rect 66637 59147 66671 59175
rect 66699 59147 68009 59175
rect 68037 59147 68071 59175
rect 68099 59147 72509 59175
rect 72537 59147 72571 59175
rect 72599 59147 75485 59175
rect 75513 59147 75547 59175
rect 75575 59147 75609 59175
rect 75637 59147 75671 59175
rect 75699 59147 77009 59175
rect 77037 59147 77071 59175
rect 77099 59147 81509 59175
rect 81537 59147 81571 59175
rect 81599 59147 84485 59175
rect 84513 59147 84547 59175
rect 84575 59147 84609 59175
rect 84637 59147 84671 59175
rect 84699 59147 86009 59175
rect 86037 59147 86071 59175
rect 86099 59147 90509 59175
rect 90537 59147 90571 59175
rect 90599 59147 95009 59175
rect 95037 59147 95071 59175
rect 95099 59147 99509 59175
rect 99537 59147 99571 59175
rect 99599 59147 104009 59175
rect 104037 59147 104071 59175
rect 104099 59147 108509 59175
rect 108537 59147 108571 59175
rect 108599 59147 113009 59175
rect 113037 59147 113071 59175
rect 113099 59147 117509 59175
rect 117537 59147 117571 59175
rect 117599 59147 120485 59175
rect 120513 59147 120547 59175
rect 120575 59147 120609 59175
rect 120637 59147 120671 59175
rect 120699 59147 129485 59175
rect 129513 59147 129547 59175
rect 129575 59147 129609 59175
rect 129637 59147 129671 59175
rect 129699 59147 138485 59175
rect 138513 59147 138547 59175
rect 138575 59147 138609 59175
rect 138637 59147 138671 59175
rect 138699 59147 147485 59175
rect 147513 59147 147547 59175
rect 147575 59147 147609 59175
rect 147637 59147 147671 59175
rect 147699 59147 156485 59175
rect 156513 59147 156547 59175
rect 156575 59147 156609 59175
rect 156637 59147 156671 59175
rect 156699 59147 165485 59175
rect 165513 59147 165547 59175
rect 165575 59147 165609 59175
rect 165637 59147 165671 59175
rect 165699 59147 174485 59175
rect 174513 59147 174547 59175
rect 174575 59147 174609 59175
rect 174637 59147 174671 59175
rect 174699 59147 183485 59175
rect 183513 59147 183547 59175
rect 183575 59147 183609 59175
rect 183637 59147 183671 59175
rect 183699 59147 192485 59175
rect 192513 59147 192547 59175
rect 192575 59147 192609 59175
rect 192637 59147 192671 59175
rect 192699 59147 201485 59175
rect 201513 59147 201547 59175
rect 201575 59147 201609 59175
rect 201637 59147 201671 59175
rect 201699 59147 210485 59175
rect 210513 59147 210547 59175
rect 210575 59147 210609 59175
rect 210637 59147 210671 59175
rect 210699 59147 219485 59175
rect 219513 59147 219547 59175
rect 219575 59147 219609 59175
rect 219637 59147 219671 59175
rect 219699 59147 228485 59175
rect 228513 59147 228547 59175
rect 228575 59147 228609 59175
rect 228637 59147 228671 59175
rect 228699 59147 237485 59175
rect 237513 59147 237547 59175
rect 237575 59147 237609 59175
rect 237637 59147 237671 59175
rect 237699 59147 246485 59175
rect 246513 59147 246547 59175
rect 246575 59147 246609 59175
rect 246637 59147 246671 59175
rect 246699 59147 255485 59175
rect 255513 59147 255547 59175
rect 255575 59147 255609 59175
rect 255637 59147 255671 59175
rect 255699 59147 264485 59175
rect 264513 59147 264547 59175
rect 264575 59147 264609 59175
rect 264637 59147 264671 59175
rect 264699 59147 273485 59175
rect 273513 59147 273547 59175
rect 273575 59147 273609 59175
rect 273637 59147 273671 59175
rect 273699 59147 282485 59175
rect 282513 59147 282547 59175
rect 282575 59147 282609 59175
rect 282637 59147 282671 59175
rect 282699 59147 291485 59175
rect 291513 59147 291547 59175
rect 291575 59147 291609 59175
rect 291637 59147 291671 59175
rect 291699 59147 298728 59175
rect 298756 59147 298790 59175
rect 298818 59147 298852 59175
rect 298880 59147 298914 59175
rect 298942 59147 298990 59175
rect -958 59113 298990 59147
rect -958 59085 -910 59113
rect -882 59085 -848 59113
rect -820 59085 -786 59113
rect -758 59085 -724 59113
rect -696 59085 3485 59113
rect 3513 59085 3547 59113
rect 3575 59085 3609 59113
rect 3637 59085 3671 59113
rect 3699 59085 12485 59113
rect 12513 59085 12547 59113
rect 12575 59085 12609 59113
rect 12637 59085 12671 59113
rect 12699 59085 21485 59113
rect 21513 59085 21547 59113
rect 21575 59085 21609 59113
rect 21637 59085 21671 59113
rect 21699 59085 30485 59113
rect 30513 59085 30547 59113
rect 30575 59085 30609 59113
rect 30637 59085 30671 59113
rect 30699 59085 39485 59113
rect 39513 59085 39547 59113
rect 39575 59085 39609 59113
rect 39637 59085 39671 59113
rect 39699 59085 48485 59113
rect 48513 59085 48547 59113
rect 48575 59085 48609 59113
rect 48637 59085 48671 59113
rect 48699 59085 54509 59113
rect 54537 59085 54571 59113
rect 54599 59085 57485 59113
rect 57513 59085 57547 59113
rect 57575 59085 57609 59113
rect 57637 59085 57671 59113
rect 57699 59085 59009 59113
rect 59037 59085 59071 59113
rect 59099 59085 63509 59113
rect 63537 59085 63571 59113
rect 63599 59085 66485 59113
rect 66513 59085 66547 59113
rect 66575 59085 66609 59113
rect 66637 59085 66671 59113
rect 66699 59085 68009 59113
rect 68037 59085 68071 59113
rect 68099 59085 72509 59113
rect 72537 59085 72571 59113
rect 72599 59085 75485 59113
rect 75513 59085 75547 59113
rect 75575 59085 75609 59113
rect 75637 59085 75671 59113
rect 75699 59085 77009 59113
rect 77037 59085 77071 59113
rect 77099 59085 81509 59113
rect 81537 59085 81571 59113
rect 81599 59085 84485 59113
rect 84513 59085 84547 59113
rect 84575 59085 84609 59113
rect 84637 59085 84671 59113
rect 84699 59085 86009 59113
rect 86037 59085 86071 59113
rect 86099 59085 90509 59113
rect 90537 59085 90571 59113
rect 90599 59085 95009 59113
rect 95037 59085 95071 59113
rect 95099 59085 99509 59113
rect 99537 59085 99571 59113
rect 99599 59085 104009 59113
rect 104037 59085 104071 59113
rect 104099 59085 108509 59113
rect 108537 59085 108571 59113
rect 108599 59085 113009 59113
rect 113037 59085 113071 59113
rect 113099 59085 117509 59113
rect 117537 59085 117571 59113
rect 117599 59085 120485 59113
rect 120513 59085 120547 59113
rect 120575 59085 120609 59113
rect 120637 59085 120671 59113
rect 120699 59085 129485 59113
rect 129513 59085 129547 59113
rect 129575 59085 129609 59113
rect 129637 59085 129671 59113
rect 129699 59085 138485 59113
rect 138513 59085 138547 59113
rect 138575 59085 138609 59113
rect 138637 59085 138671 59113
rect 138699 59085 147485 59113
rect 147513 59085 147547 59113
rect 147575 59085 147609 59113
rect 147637 59085 147671 59113
rect 147699 59085 156485 59113
rect 156513 59085 156547 59113
rect 156575 59085 156609 59113
rect 156637 59085 156671 59113
rect 156699 59085 165485 59113
rect 165513 59085 165547 59113
rect 165575 59085 165609 59113
rect 165637 59085 165671 59113
rect 165699 59085 174485 59113
rect 174513 59085 174547 59113
rect 174575 59085 174609 59113
rect 174637 59085 174671 59113
rect 174699 59085 183485 59113
rect 183513 59085 183547 59113
rect 183575 59085 183609 59113
rect 183637 59085 183671 59113
rect 183699 59085 192485 59113
rect 192513 59085 192547 59113
rect 192575 59085 192609 59113
rect 192637 59085 192671 59113
rect 192699 59085 201485 59113
rect 201513 59085 201547 59113
rect 201575 59085 201609 59113
rect 201637 59085 201671 59113
rect 201699 59085 210485 59113
rect 210513 59085 210547 59113
rect 210575 59085 210609 59113
rect 210637 59085 210671 59113
rect 210699 59085 219485 59113
rect 219513 59085 219547 59113
rect 219575 59085 219609 59113
rect 219637 59085 219671 59113
rect 219699 59085 228485 59113
rect 228513 59085 228547 59113
rect 228575 59085 228609 59113
rect 228637 59085 228671 59113
rect 228699 59085 237485 59113
rect 237513 59085 237547 59113
rect 237575 59085 237609 59113
rect 237637 59085 237671 59113
rect 237699 59085 246485 59113
rect 246513 59085 246547 59113
rect 246575 59085 246609 59113
rect 246637 59085 246671 59113
rect 246699 59085 255485 59113
rect 255513 59085 255547 59113
rect 255575 59085 255609 59113
rect 255637 59085 255671 59113
rect 255699 59085 264485 59113
rect 264513 59085 264547 59113
rect 264575 59085 264609 59113
rect 264637 59085 264671 59113
rect 264699 59085 273485 59113
rect 273513 59085 273547 59113
rect 273575 59085 273609 59113
rect 273637 59085 273671 59113
rect 273699 59085 282485 59113
rect 282513 59085 282547 59113
rect 282575 59085 282609 59113
rect 282637 59085 282671 59113
rect 282699 59085 291485 59113
rect 291513 59085 291547 59113
rect 291575 59085 291609 59113
rect 291637 59085 291671 59113
rect 291699 59085 298728 59113
rect 298756 59085 298790 59113
rect 298818 59085 298852 59113
rect 298880 59085 298914 59113
rect 298942 59085 298990 59113
rect -958 59051 298990 59085
rect -958 59023 -910 59051
rect -882 59023 -848 59051
rect -820 59023 -786 59051
rect -758 59023 -724 59051
rect -696 59023 3485 59051
rect 3513 59023 3547 59051
rect 3575 59023 3609 59051
rect 3637 59023 3671 59051
rect 3699 59023 12485 59051
rect 12513 59023 12547 59051
rect 12575 59023 12609 59051
rect 12637 59023 12671 59051
rect 12699 59023 21485 59051
rect 21513 59023 21547 59051
rect 21575 59023 21609 59051
rect 21637 59023 21671 59051
rect 21699 59023 30485 59051
rect 30513 59023 30547 59051
rect 30575 59023 30609 59051
rect 30637 59023 30671 59051
rect 30699 59023 39485 59051
rect 39513 59023 39547 59051
rect 39575 59023 39609 59051
rect 39637 59023 39671 59051
rect 39699 59023 48485 59051
rect 48513 59023 48547 59051
rect 48575 59023 48609 59051
rect 48637 59023 48671 59051
rect 48699 59023 54509 59051
rect 54537 59023 54571 59051
rect 54599 59023 57485 59051
rect 57513 59023 57547 59051
rect 57575 59023 57609 59051
rect 57637 59023 57671 59051
rect 57699 59023 59009 59051
rect 59037 59023 59071 59051
rect 59099 59023 63509 59051
rect 63537 59023 63571 59051
rect 63599 59023 66485 59051
rect 66513 59023 66547 59051
rect 66575 59023 66609 59051
rect 66637 59023 66671 59051
rect 66699 59023 68009 59051
rect 68037 59023 68071 59051
rect 68099 59023 72509 59051
rect 72537 59023 72571 59051
rect 72599 59023 75485 59051
rect 75513 59023 75547 59051
rect 75575 59023 75609 59051
rect 75637 59023 75671 59051
rect 75699 59023 77009 59051
rect 77037 59023 77071 59051
rect 77099 59023 81509 59051
rect 81537 59023 81571 59051
rect 81599 59023 84485 59051
rect 84513 59023 84547 59051
rect 84575 59023 84609 59051
rect 84637 59023 84671 59051
rect 84699 59023 86009 59051
rect 86037 59023 86071 59051
rect 86099 59023 90509 59051
rect 90537 59023 90571 59051
rect 90599 59023 95009 59051
rect 95037 59023 95071 59051
rect 95099 59023 99509 59051
rect 99537 59023 99571 59051
rect 99599 59023 104009 59051
rect 104037 59023 104071 59051
rect 104099 59023 108509 59051
rect 108537 59023 108571 59051
rect 108599 59023 113009 59051
rect 113037 59023 113071 59051
rect 113099 59023 117509 59051
rect 117537 59023 117571 59051
rect 117599 59023 120485 59051
rect 120513 59023 120547 59051
rect 120575 59023 120609 59051
rect 120637 59023 120671 59051
rect 120699 59023 129485 59051
rect 129513 59023 129547 59051
rect 129575 59023 129609 59051
rect 129637 59023 129671 59051
rect 129699 59023 138485 59051
rect 138513 59023 138547 59051
rect 138575 59023 138609 59051
rect 138637 59023 138671 59051
rect 138699 59023 147485 59051
rect 147513 59023 147547 59051
rect 147575 59023 147609 59051
rect 147637 59023 147671 59051
rect 147699 59023 156485 59051
rect 156513 59023 156547 59051
rect 156575 59023 156609 59051
rect 156637 59023 156671 59051
rect 156699 59023 165485 59051
rect 165513 59023 165547 59051
rect 165575 59023 165609 59051
rect 165637 59023 165671 59051
rect 165699 59023 174485 59051
rect 174513 59023 174547 59051
rect 174575 59023 174609 59051
rect 174637 59023 174671 59051
rect 174699 59023 183485 59051
rect 183513 59023 183547 59051
rect 183575 59023 183609 59051
rect 183637 59023 183671 59051
rect 183699 59023 192485 59051
rect 192513 59023 192547 59051
rect 192575 59023 192609 59051
rect 192637 59023 192671 59051
rect 192699 59023 201485 59051
rect 201513 59023 201547 59051
rect 201575 59023 201609 59051
rect 201637 59023 201671 59051
rect 201699 59023 210485 59051
rect 210513 59023 210547 59051
rect 210575 59023 210609 59051
rect 210637 59023 210671 59051
rect 210699 59023 219485 59051
rect 219513 59023 219547 59051
rect 219575 59023 219609 59051
rect 219637 59023 219671 59051
rect 219699 59023 228485 59051
rect 228513 59023 228547 59051
rect 228575 59023 228609 59051
rect 228637 59023 228671 59051
rect 228699 59023 237485 59051
rect 237513 59023 237547 59051
rect 237575 59023 237609 59051
rect 237637 59023 237671 59051
rect 237699 59023 246485 59051
rect 246513 59023 246547 59051
rect 246575 59023 246609 59051
rect 246637 59023 246671 59051
rect 246699 59023 255485 59051
rect 255513 59023 255547 59051
rect 255575 59023 255609 59051
rect 255637 59023 255671 59051
rect 255699 59023 264485 59051
rect 264513 59023 264547 59051
rect 264575 59023 264609 59051
rect 264637 59023 264671 59051
rect 264699 59023 273485 59051
rect 273513 59023 273547 59051
rect 273575 59023 273609 59051
rect 273637 59023 273671 59051
rect 273699 59023 282485 59051
rect 282513 59023 282547 59051
rect 282575 59023 282609 59051
rect 282637 59023 282671 59051
rect 282699 59023 291485 59051
rect 291513 59023 291547 59051
rect 291575 59023 291609 59051
rect 291637 59023 291671 59051
rect 291699 59023 298728 59051
rect 298756 59023 298790 59051
rect 298818 59023 298852 59051
rect 298880 59023 298914 59051
rect 298942 59023 298990 59051
rect -958 58989 298990 59023
rect -958 58961 -910 58989
rect -882 58961 -848 58989
rect -820 58961 -786 58989
rect -758 58961 -724 58989
rect -696 58961 3485 58989
rect 3513 58961 3547 58989
rect 3575 58961 3609 58989
rect 3637 58961 3671 58989
rect 3699 58961 12485 58989
rect 12513 58961 12547 58989
rect 12575 58961 12609 58989
rect 12637 58961 12671 58989
rect 12699 58961 21485 58989
rect 21513 58961 21547 58989
rect 21575 58961 21609 58989
rect 21637 58961 21671 58989
rect 21699 58961 30485 58989
rect 30513 58961 30547 58989
rect 30575 58961 30609 58989
rect 30637 58961 30671 58989
rect 30699 58961 39485 58989
rect 39513 58961 39547 58989
rect 39575 58961 39609 58989
rect 39637 58961 39671 58989
rect 39699 58961 48485 58989
rect 48513 58961 48547 58989
rect 48575 58961 48609 58989
rect 48637 58961 48671 58989
rect 48699 58961 54509 58989
rect 54537 58961 54571 58989
rect 54599 58961 57485 58989
rect 57513 58961 57547 58989
rect 57575 58961 57609 58989
rect 57637 58961 57671 58989
rect 57699 58961 59009 58989
rect 59037 58961 59071 58989
rect 59099 58961 63509 58989
rect 63537 58961 63571 58989
rect 63599 58961 66485 58989
rect 66513 58961 66547 58989
rect 66575 58961 66609 58989
rect 66637 58961 66671 58989
rect 66699 58961 68009 58989
rect 68037 58961 68071 58989
rect 68099 58961 72509 58989
rect 72537 58961 72571 58989
rect 72599 58961 75485 58989
rect 75513 58961 75547 58989
rect 75575 58961 75609 58989
rect 75637 58961 75671 58989
rect 75699 58961 77009 58989
rect 77037 58961 77071 58989
rect 77099 58961 81509 58989
rect 81537 58961 81571 58989
rect 81599 58961 84485 58989
rect 84513 58961 84547 58989
rect 84575 58961 84609 58989
rect 84637 58961 84671 58989
rect 84699 58961 86009 58989
rect 86037 58961 86071 58989
rect 86099 58961 90509 58989
rect 90537 58961 90571 58989
rect 90599 58961 95009 58989
rect 95037 58961 95071 58989
rect 95099 58961 99509 58989
rect 99537 58961 99571 58989
rect 99599 58961 104009 58989
rect 104037 58961 104071 58989
rect 104099 58961 108509 58989
rect 108537 58961 108571 58989
rect 108599 58961 113009 58989
rect 113037 58961 113071 58989
rect 113099 58961 117509 58989
rect 117537 58961 117571 58989
rect 117599 58961 120485 58989
rect 120513 58961 120547 58989
rect 120575 58961 120609 58989
rect 120637 58961 120671 58989
rect 120699 58961 129485 58989
rect 129513 58961 129547 58989
rect 129575 58961 129609 58989
rect 129637 58961 129671 58989
rect 129699 58961 138485 58989
rect 138513 58961 138547 58989
rect 138575 58961 138609 58989
rect 138637 58961 138671 58989
rect 138699 58961 147485 58989
rect 147513 58961 147547 58989
rect 147575 58961 147609 58989
rect 147637 58961 147671 58989
rect 147699 58961 156485 58989
rect 156513 58961 156547 58989
rect 156575 58961 156609 58989
rect 156637 58961 156671 58989
rect 156699 58961 165485 58989
rect 165513 58961 165547 58989
rect 165575 58961 165609 58989
rect 165637 58961 165671 58989
rect 165699 58961 174485 58989
rect 174513 58961 174547 58989
rect 174575 58961 174609 58989
rect 174637 58961 174671 58989
rect 174699 58961 183485 58989
rect 183513 58961 183547 58989
rect 183575 58961 183609 58989
rect 183637 58961 183671 58989
rect 183699 58961 192485 58989
rect 192513 58961 192547 58989
rect 192575 58961 192609 58989
rect 192637 58961 192671 58989
rect 192699 58961 201485 58989
rect 201513 58961 201547 58989
rect 201575 58961 201609 58989
rect 201637 58961 201671 58989
rect 201699 58961 210485 58989
rect 210513 58961 210547 58989
rect 210575 58961 210609 58989
rect 210637 58961 210671 58989
rect 210699 58961 219485 58989
rect 219513 58961 219547 58989
rect 219575 58961 219609 58989
rect 219637 58961 219671 58989
rect 219699 58961 228485 58989
rect 228513 58961 228547 58989
rect 228575 58961 228609 58989
rect 228637 58961 228671 58989
rect 228699 58961 237485 58989
rect 237513 58961 237547 58989
rect 237575 58961 237609 58989
rect 237637 58961 237671 58989
rect 237699 58961 246485 58989
rect 246513 58961 246547 58989
rect 246575 58961 246609 58989
rect 246637 58961 246671 58989
rect 246699 58961 255485 58989
rect 255513 58961 255547 58989
rect 255575 58961 255609 58989
rect 255637 58961 255671 58989
rect 255699 58961 264485 58989
rect 264513 58961 264547 58989
rect 264575 58961 264609 58989
rect 264637 58961 264671 58989
rect 264699 58961 273485 58989
rect 273513 58961 273547 58989
rect 273575 58961 273609 58989
rect 273637 58961 273671 58989
rect 273699 58961 282485 58989
rect 282513 58961 282547 58989
rect 282575 58961 282609 58989
rect 282637 58961 282671 58989
rect 282699 58961 291485 58989
rect 291513 58961 291547 58989
rect 291575 58961 291609 58989
rect 291637 58961 291671 58989
rect 291699 58961 298728 58989
rect 298756 58961 298790 58989
rect 298818 58961 298852 58989
rect 298880 58961 298914 58989
rect 298942 58961 298990 58989
rect -958 58913 298990 58961
rect -958 56175 298990 56223
rect -958 56147 -430 56175
rect -402 56147 -368 56175
rect -340 56147 -306 56175
rect -278 56147 -244 56175
rect -216 56147 1625 56175
rect 1653 56147 1687 56175
rect 1715 56147 1749 56175
rect 1777 56147 1811 56175
rect 1839 56147 10625 56175
rect 10653 56147 10687 56175
rect 10715 56147 10749 56175
rect 10777 56147 10811 56175
rect 10839 56147 19625 56175
rect 19653 56147 19687 56175
rect 19715 56147 19749 56175
rect 19777 56147 19811 56175
rect 19839 56147 28625 56175
rect 28653 56147 28687 56175
rect 28715 56147 28749 56175
rect 28777 56147 28811 56175
rect 28839 56147 37625 56175
rect 37653 56147 37687 56175
rect 37715 56147 37749 56175
rect 37777 56147 37811 56175
rect 37839 56147 46625 56175
rect 46653 56147 46687 56175
rect 46715 56147 46749 56175
rect 46777 56147 46811 56175
rect 46839 56147 52259 56175
rect 52287 56147 52321 56175
rect 52349 56147 55625 56175
rect 55653 56147 55687 56175
rect 55715 56147 55749 56175
rect 55777 56147 55811 56175
rect 55839 56147 56759 56175
rect 56787 56147 56821 56175
rect 56849 56147 61259 56175
rect 61287 56147 61321 56175
rect 61349 56147 64625 56175
rect 64653 56147 64687 56175
rect 64715 56147 64749 56175
rect 64777 56147 64811 56175
rect 64839 56147 65759 56175
rect 65787 56147 65821 56175
rect 65849 56147 70259 56175
rect 70287 56147 70321 56175
rect 70349 56147 73625 56175
rect 73653 56147 73687 56175
rect 73715 56147 73749 56175
rect 73777 56147 73811 56175
rect 73839 56147 74759 56175
rect 74787 56147 74821 56175
rect 74849 56147 79259 56175
rect 79287 56147 79321 56175
rect 79349 56147 82625 56175
rect 82653 56147 82687 56175
rect 82715 56147 82749 56175
rect 82777 56147 82811 56175
rect 82839 56147 83759 56175
rect 83787 56147 83821 56175
rect 83849 56147 88259 56175
rect 88287 56147 88321 56175
rect 88349 56147 91625 56175
rect 91653 56147 91687 56175
rect 91715 56147 91749 56175
rect 91777 56147 91811 56175
rect 91839 56147 92759 56175
rect 92787 56147 92821 56175
rect 92849 56147 97259 56175
rect 97287 56147 97321 56175
rect 97349 56147 101759 56175
rect 101787 56147 101821 56175
rect 101849 56147 106259 56175
rect 106287 56147 106321 56175
rect 106349 56147 110759 56175
rect 110787 56147 110821 56175
rect 110849 56147 115259 56175
rect 115287 56147 115321 56175
rect 115349 56147 127625 56175
rect 127653 56147 127687 56175
rect 127715 56147 127749 56175
rect 127777 56147 127811 56175
rect 127839 56147 136625 56175
rect 136653 56147 136687 56175
rect 136715 56147 136749 56175
rect 136777 56147 136811 56175
rect 136839 56147 145625 56175
rect 145653 56147 145687 56175
rect 145715 56147 145749 56175
rect 145777 56147 145811 56175
rect 145839 56147 154625 56175
rect 154653 56147 154687 56175
rect 154715 56147 154749 56175
rect 154777 56147 154811 56175
rect 154839 56147 163625 56175
rect 163653 56147 163687 56175
rect 163715 56147 163749 56175
rect 163777 56147 163811 56175
rect 163839 56147 172625 56175
rect 172653 56147 172687 56175
rect 172715 56147 172749 56175
rect 172777 56147 172811 56175
rect 172839 56147 181625 56175
rect 181653 56147 181687 56175
rect 181715 56147 181749 56175
rect 181777 56147 181811 56175
rect 181839 56147 190625 56175
rect 190653 56147 190687 56175
rect 190715 56147 190749 56175
rect 190777 56147 190811 56175
rect 190839 56147 199625 56175
rect 199653 56147 199687 56175
rect 199715 56147 199749 56175
rect 199777 56147 199811 56175
rect 199839 56147 208625 56175
rect 208653 56147 208687 56175
rect 208715 56147 208749 56175
rect 208777 56147 208811 56175
rect 208839 56147 217625 56175
rect 217653 56147 217687 56175
rect 217715 56147 217749 56175
rect 217777 56147 217811 56175
rect 217839 56147 226625 56175
rect 226653 56147 226687 56175
rect 226715 56147 226749 56175
rect 226777 56147 226811 56175
rect 226839 56147 235625 56175
rect 235653 56147 235687 56175
rect 235715 56147 235749 56175
rect 235777 56147 235811 56175
rect 235839 56147 244625 56175
rect 244653 56147 244687 56175
rect 244715 56147 244749 56175
rect 244777 56147 244811 56175
rect 244839 56147 253625 56175
rect 253653 56147 253687 56175
rect 253715 56147 253749 56175
rect 253777 56147 253811 56175
rect 253839 56147 262625 56175
rect 262653 56147 262687 56175
rect 262715 56147 262749 56175
rect 262777 56147 262811 56175
rect 262839 56147 271625 56175
rect 271653 56147 271687 56175
rect 271715 56147 271749 56175
rect 271777 56147 271811 56175
rect 271839 56147 280625 56175
rect 280653 56147 280687 56175
rect 280715 56147 280749 56175
rect 280777 56147 280811 56175
rect 280839 56147 289625 56175
rect 289653 56147 289687 56175
rect 289715 56147 289749 56175
rect 289777 56147 289811 56175
rect 289839 56147 298248 56175
rect 298276 56147 298310 56175
rect 298338 56147 298372 56175
rect 298400 56147 298434 56175
rect 298462 56147 298990 56175
rect -958 56113 298990 56147
rect -958 56085 -430 56113
rect -402 56085 -368 56113
rect -340 56085 -306 56113
rect -278 56085 -244 56113
rect -216 56085 1625 56113
rect 1653 56085 1687 56113
rect 1715 56085 1749 56113
rect 1777 56085 1811 56113
rect 1839 56085 10625 56113
rect 10653 56085 10687 56113
rect 10715 56085 10749 56113
rect 10777 56085 10811 56113
rect 10839 56085 19625 56113
rect 19653 56085 19687 56113
rect 19715 56085 19749 56113
rect 19777 56085 19811 56113
rect 19839 56085 28625 56113
rect 28653 56085 28687 56113
rect 28715 56085 28749 56113
rect 28777 56085 28811 56113
rect 28839 56085 37625 56113
rect 37653 56085 37687 56113
rect 37715 56085 37749 56113
rect 37777 56085 37811 56113
rect 37839 56085 46625 56113
rect 46653 56085 46687 56113
rect 46715 56085 46749 56113
rect 46777 56085 46811 56113
rect 46839 56085 52259 56113
rect 52287 56085 52321 56113
rect 52349 56085 55625 56113
rect 55653 56085 55687 56113
rect 55715 56085 55749 56113
rect 55777 56085 55811 56113
rect 55839 56085 56759 56113
rect 56787 56085 56821 56113
rect 56849 56085 61259 56113
rect 61287 56085 61321 56113
rect 61349 56085 64625 56113
rect 64653 56085 64687 56113
rect 64715 56085 64749 56113
rect 64777 56085 64811 56113
rect 64839 56085 65759 56113
rect 65787 56085 65821 56113
rect 65849 56085 70259 56113
rect 70287 56085 70321 56113
rect 70349 56085 73625 56113
rect 73653 56085 73687 56113
rect 73715 56085 73749 56113
rect 73777 56085 73811 56113
rect 73839 56085 74759 56113
rect 74787 56085 74821 56113
rect 74849 56085 79259 56113
rect 79287 56085 79321 56113
rect 79349 56085 82625 56113
rect 82653 56085 82687 56113
rect 82715 56085 82749 56113
rect 82777 56085 82811 56113
rect 82839 56085 83759 56113
rect 83787 56085 83821 56113
rect 83849 56085 88259 56113
rect 88287 56085 88321 56113
rect 88349 56085 91625 56113
rect 91653 56085 91687 56113
rect 91715 56085 91749 56113
rect 91777 56085 91811 56113
rect 91839 56085 92759 56113
rect 92787 56085 92821 56113
rect 92849 56085 97259 56113
rect 97287 56085 97321 56113
rect 97349 56085 101759 56113
rect 101787 56085 101821 56113
rect 101849 56085 106259 56113
rect 106287 56085 106321 56113
rect 106349 56085 110759 56113
rect 110787 56085 110821 56113
rect 110849 56085 115259 56113
rect 115287 56085 115321 56113
rect 115349 56085 127625 56113
rect 127653 56085 127687 56113
rect 127715 56085 127749 56113
rect 127777 56085 127811 56113
rect 127839 56085 136625 56113
rect 136653 56085 136687 56113
rect 136715 56085 136749 56113
rect 136777 56085 136811 56113
rect 136839 56085 145625 56113
rect 145653 56085 145687 56113
rect 145715 56085 145749 56113
rect 145777 56085 145811 56113
rect 145839 56085 154625 56113
rect 154653 56085 154687 56113
rect 154715 56085 154749 56113
rect 154777 56085 154811 56113
rect 154839 56085 163625 56113
rect 163653 56085 163687 56113
rect 163715 56085 163749 56113
rect 163777 56085 163811 56113
rect 163839 56085 172625 56113
rect 172653 56085 172687 56113
rect 172715 56085 172749 56113
rect 172777 56085 172811 56113
rect 172839 56085 181625 56113
rect 181653 56085 181687 56113
rect 181715 56085 181749 56113
rect 181777 56085 181811 56113
rect 181839 56085 190625 56113
rect 190653 56085 190687 56113
rect 190715 56085 190749 56113
rect 190777 56085 190811 56113
rect 190839 56085 199625 56113
rect 199653 56085 199687 56113
rect 199715 56085 199749 56113
rect 199777 56085 199811 56113
rect 199839 56085 208625 56113
rect 208653 56085 208687 56113
rect 208715 56085 208749 56113
rect 208777 56085 208811 56113
rect 208839 56085 217625 56113
rect 217653 56085 217687 56113
rect 217715 56085 217749 56113
rect 217777 56085 217811 56113
rect 217839 56085 226625 56113
rect 226653 56085 226687 56113
rect 226715 56085 226749 56113
rect 226777 56085 226811 56113
rect 226839 56085 235625 56113
rect 235653 56085 235687 56113
rect 235715 56085 235749 56113
rect 235777 56085 235811 56113
rect 235839 56085 244625 56113
rect 244653 56085 244687 56113
rect 244715 56085 244749 56113
rect 244777 56085 244811 56113
rect 244839 56085 253625 56113
rect 253653 56085 253687 56113
rect 253715 56085 253749 56113
rect 253777 56085 253811 56113
rect 253839 56085 262625 56113
rect 262653 56085 262687 56113
rect 262715 56085 262749 56113
rect 262777 56085 262811 56113
rect 262839 56085 271625 56113
rect 271653 56085 271687 56113
rect 271715 56085 271749 56113
rect 271777 56085 271811 56113
rect 271839 56085 280625 56113
rect 280653 56085 280687 56113
rect 280715 56085 280749 56113
rect 280777 56085 280811 56113
rect 280839 56085 289625 56113
rect 289653 56085 289687 56113
rect 289715 56085 289749 56113
rect 289777 56085 289811 56113
rect 289839 56085 298248 56113
rect 298276 56085 298310 56113
rect 298338 56085 298372 56113
rect 298400 56085 298434 56113
rect 298462 56085 298990 56113
rect -958 56051 298990 56085
rect -958 56023 -430 56051
rect -402 56023 -368 56051
rect -340 56023 -306 56051
rect -278 56023 -244 56051
rect -216 56023 1625 56051
rect 1653 56023 1687 56051
rect 1715 56023 1749 56051
rect 1777 56023 1811 56051
rect 1839 56023 10625 56051
rect 10653 56023 10687 56051
rect 10715 56023 10749 56051
rect 10777 56023 10811 56051
rect 10839 56023 19625 56051
rect 19653 56023 19687 56051
rect 19715 56023 19749 56051
rect 19777 56023 19811 56051
rect 19839 56023 28625 56051
rect 28653 56023 28687 56051
rect 28715 56023 28749 56051
rect 28777 56023 28811 56051
rect 28839 56023 37625 56051
rect 37653 56023 37687 56051
rect 37715 56023 37749 56051
rect 37777 56023 37811 56051
rect 37839 56023 46625 56051
rect 46653 56023 46687 56051
rect 46715 56023 46749 56051
rect 46777 56023 46811 56051
rect 46839 56023 52259 56051
rect 52287 56023 52321 56051
rect 52349 56023 55625 56051
rect 55653 56023 55687 56051
rect 55715 56023 55749 56051
rect 55777 56023 55811 56051
rect 55839 56023 56759 56051
rect 56787 56023 56821 56051
rect 56849 56023 61259 56051
rect 61287 56023 61321 56051
rect 61349 56023 64625 56051
rect 64653 56023 64687 56051
rect 64715 56023 64749 56051
rect 64777 56023 64811 56051
rect 64839 56023 65759 56051
rect 65787 56023 65821 56051
rect 65849 56023 70259 56051
rect 70287 56023 70321 56051
rect 70349 56023 73625 56051
rect 73653 56023 73687 56051
rect 73715 56023 73749 56051
rect 73777 56023 73811 56051
rect 73839 56023 74759 56051
rect 74787 56023 74821 56051
rect 74849 56023 79259 56051
rect 79287 56023 79321 56051
rect 79349 56023 82625 56051
rect 82653 56023 82687 56051
rect 82715 56023 82749 56051
rect 82777 56023 82811 56051
rect 82839 56023 83759 56051
rect 83787 56023 83821 56051
rect 83849 56023 88259 56051
rect 88287 56023 88321 56051
rect 88349 56023 91625 56051
rect 91653 56023 91687 56051
rect 91715 56023 91749 56051
rect 91777 56023 91811 56051
rect 91839 56023 92759 56051
rect 92787 56023 92821 56051
rect 92849 56023 97259 56051
rect 97287 56023 97321 56051
rect 97349 56023 101759 56051
rect 101787 56023 101821 56051
rect 101849 56023 106259 56051
rect 106287 56023 106321 56051
rect 106349 56023 110759 56051
rect 110787 56023 110821 56051
rect 110849 56023 115259 56051
rect 115287 56023 115321 56051
rect 115349 56023 127625 56051
rect 127653 56023 127687 56051
rect 127715 56023 127749 56051
rect 127777 56023 127811 56051
rect 127839 56023 136625 56051
rect 136653 56023 136687 56051
rect 136715 56023 136749 56051
rect 136777 56023 136811 56051
rect 136839 56023 145625 56051
rect 145653 56023 145687 56051
rect 145715 56023 145749 56051
rect 145777 56023 145811 56051
rect 145839 56023 154625 56051
rect 154653 56023 154687 56051
rect 154715 56023 154749 56051
rect 154777 56023 154811 56051
rect 154839 56023 163625 56051
rect 163653 56023 163687 56051
rect 163715 56023 163749 56051
rect 163777 56023 163811 56051
rect 163839 56023 172625 56051
rect 172653 56023 172687 56051
rect 172715 56023 172749 56051
rect 172777 56023 172811 56051
rect 172839 56023 181625 56051
rect 181653 56023 181687 56051
rect 181715 56023 181749 56051
rect 181777 56023 181811 56051
rect 181839 56023 190625 56051
rect 190653 56023 190687 56051
rect 190715 56023 190749 56051
rect 190777 56023 190811 56051
rect 190839 56023 199625 56051
rect 199653 56023 199687 56051
rect 199715 56023 199749 56051
rect 199777 56023 199811 56051
rect 199839 56023 208625 56051
rect 208653 56023 208687 56051
rect 208715 56023 208749 56051
rect 208777 56023 208811 56051
rect 208839 56023 217625 56051
rect 217653 56023 217687 56051
rect 217715 56023 217749 56051
rect 217777 56023 217811 56051
rect 217839 56023 226625 56051
rect 226653 56023 226687 56051
rect 226715 56023 226749 56051
rect 226777 56023 226811 56051
rect 226839 56023 235625 56051
rect 235653 56023 235687 56051
rect 235715 56023 235749 56051
rect 235777 56023 235811 56051
rect 235839 56023 244625 56051
rect 244653 56023 244687 56051
rect 244715 56023 244749 56051
rect 244777 56023 244811 56051
rect 244839 56023 253625 56051
rect 253653 56023 253687 56051
rect 253715 56023 253749 56051
rect 253777 56023 253811 56051
rect 253839 56023 262625 56051
rect 262653 56023 262687 56051
rect 262715 56023 262749 56051
rect 262777 56023 262811 56051
rect 262839 56023 271625 56051
rect 271653 56023 271687 56051
rect 271715 56023 271749 56051
rect 271777 56023 271811 56051
rect 271839 56023 280625 56051
rect 280653 56023 280687 56051
rect 280715 56023 280749 56051
rect 280777 56023 280811 56051
rect 280839 56023 289625 56051
rect 289653 56023 289687 56051
rect 289715 56023 289749 56051
rect 289777 56023 289811 56051
rect 289839 56023 298248 56051
rect 298276 56023 298310 56051
rect 298338 56023 298372 56051
rect 298400 56023 298434 56051
rect 298462 56023 298990 56051
rect -958 55989 298990 56023
rect -958 55961 -430 55989
rect -402 55961 -368 55989
rect -340 55961 -306 55989
rect -278 55961 -244 55989
rect -216 55961 1625 55989
rect 1653 55961 1687 55989
rect 1715 55961 1749 55989
rect 1777 55961 1811 55989
rect 1839 55961 10625 55989
rect 10653 55961 10687 55989
rect 10715 55961 10749 55989
rect 10777 55961 10811 55989
rect 10839 55961 19625 55989
rect 19653 55961 19687 55989
rect 19715 55961 19749 55989
rect 19777 55961 19811 55989
rect 19839 55961 28625 55989
rect 28653 55961 28687 55989
rect 28715 55961 28749 55989
rect 28777 55961 28811 55989
rect 28839 55961 37625 55989
rect 37653 55961 37687 55989
rect 37715 55961 37749 55989
rect 37777 55961 37811 55989
rect 37839 55961 46625 55989
rect 46653 55961 46687 55989
rect 46715 55961 46749 55989
rect 46777 55961 46811 55989
rect 46839 55961 52259 55989
rect 52287 55961 52321 55989
rect 52349 55961 55625 55989
rect 55653 55961 55687 55989
rect 55715 55961 55749 55989
rect 55777 55961 55811 55989
rect 55839 55961 56759 55989
rect 56787 55961 56821 55989
rect 56849 55961 61259 55989
rect 61287 55961 61321 55989
rect 61349 55961 64625 55989
rect 64653 55961 64687 55989
rect 64715 55961 64749 55989
rect 64777 55961 64811 55989
rect 64839 55961 65759 55989
rect 65787 55961 65821 55989
rect 65849 55961 70259 55989
rect 70287 55961 70321 55989
rect 70349 55961 73625 55989
rect 73653 55961 73687 55989
rect 73715 55961 73749 55989
rect 73777 55961 73811 55989
rect 73839 55961 74759 55989
rect 74787 55961 74821 55989
rect 74849 55961 79259 55989
rect 79287 55961 79321 55989
rect 79349 55961 82625 55989
rect 82653 55961 82687 55989
rect 82715 55961 82749 55989
rect 82777 55961 82811 55989
rect 82839 55961 83759 55989
rect 83787 55961 83821 55989
rect 83849 55961 88259 55989
rect 88287 55961 88321 55989
rect 88349 55961 91625 55989
rect 91653 55961 91687 55989
rect 91715 55961 91749 55989
rect 91777 55961 91811 55989
rect 91839 55961 92759 55989
rect 92787 55961 92821 55989
rect 92849 55961 97259 55989
rect 97287 55961 97321 55989
rect 97349 55961 101759 55989
rect 101787 55961 101821 55989
rect 101849 55961 106259 55989
rect 106287 55961 106321 55989
rect 106349 55961 110759 55989
rect 110787 55961 110821 55989
rect 110849 55961 115259 55989
rect 115287 55961 115321 55989
rect 115349 55961 127625 55989
rect 127653 55961 127687 55989
rect 127715 55961 127749 55989
rect 127777 55961 127811 55989
rect 127839 55961 136625 55989
rect 136653 55961 136687 55989
rect 136715 55961 136749 55989
rect 136777 55961 136811 55989
rect 136839 55961 145625 55989
rect 145653 55961 145687 55989
rect 145715 55961 145749 55989
rect 145777 55961 145811 55989
rect 145839 55961 154625 55989
rect 154653 55961 154687 55989
rect 154715 55961 154749 55989
rect 154777 55961 154811 55989
rect 154839 55961 163625 55989
rect 163653 55961 163687 55989
rect 163715 55961 163749 55989
rect 163777 55961 163811 55989
rect 163839 55961 172625 55989
rect 172653 55961 172687 55989
rect 172715 55961 172749 55989
rect 172777 55961 172811 55989
rect 172839 55961 181625 55989
rect 181653 55961 181687 55989
rect 181715 55961 181749 55989
rect 181777 55961 181811 55989
rect 181839 55961 190625 55989
rect 190653 55961 190687 55989
rect 190715 55961 190749 55989
rect 190777 55961 190811 55989
rect 190839 55961 199625 55989
rect 199653 55961 199687 55989
rect 199715 55961 199749 55989
rect 199777 55961 199811 55989
rect 199839 55961 208625 55989
rect 208653 55961 208687 55989
rect 208715 55961 208749 55989
rect 208777 55961 208811 55989
rect 208839 55961 217625 55989
rect 217653 55961 217687 55989
rect 217715 55961 217749 55989
rect 217777 55961 217811 55989
rect 217839 55961 226625 55989
rect 226653 55961 226687 55989
rect 226715 55961 226749 55989
rect 226777 55961 226811 55989
rect 226839 55961 235625 55989
rect 235653 55961 235687 55989
rect 235715 55961 235749 55989
rect 235777 55961 235811 55989
rect 235839 55961 244625 55989
rect 244653 55961 244687 55989
rect 244715 55961 244749 55989
rect 244777 55961 244811 55989
rect 244839 55961 253625 55989
rect 253653 55961 253687 55989
rect 253715 55961 253749 55989
rect 253777 55961 253811 55989
rect 253839 55961 262625 55989
rect 262653 55961 262687 55989
rect 262715 55961 262749 55989
rect 262777 55961 262811 55989
rect 262839 55961 271625 55989
rect 271653 55961 271687 55989
rect 271715 55961 271749 55989
rect 271777 55961 271811 55989
rect 271839 55961 280625 55989
rect 280653 55961 280687 55989
rect 280715 55961 280749 55989
rect 280777 55961 280811 55989
rect 280839 55961 289625 55989
rect 289653 55961 289687 55989
rect 289715 55961 289749 55989
rect 289777 55961 289811 55989
rect 289839 55961 298248 55989
rect 298276 55961 298310 55989
rect 298338 55961 298372 55989
rect 298400 55961 298434 55989
rect 298462 55961 298990 55989
rect -958 55913 298990 55961
rect -958 50175 298990 50223
rect -958 50147 -910 50175
rect -882 50147 -848 50175
rect -820 50147 -786 50175
rect -758 50147 -724 50175
rect -696 50147 3485 50175
rect 3513 50147 3547 50175
rect 3575 50147 3609 50175
rect 3637 50147 3671 50175
rect 3699 50147 12485 50175
rect 12513 50147 12547 50175
rect 12575 50147 12609 50175
rect 12637 50147 12671 50175
rect 12699 50147 21485 50175
rect 21513 50147 21547 50175
rect 21575 50147 21609 50175
rect 21637 50147 21671 50175
rect 21699 50147 30485 50175
rect 30513 50147 30547 50175
rect 30575 50147 30609 50175
rect 30637 50147 30671 50175
rect 30699 50147 39485 50175
rect 39513 50147 39547 50175
rect 39575 50147 39609 50175
rect 39637 50147 39671 50175
rect 39699 50147 48485 50175
rect 48513 50147 48547 50175
rect 48575 50147 48609 50175
rect 48637 50147 48671 50175
rect 48699 50147 57485 50175
rect 57513 50147 57547 50175
rect 57575 50147 57609 50175
rect 57637 50147 57671 50175
rect 57699 50147 66485 50175
rect 66513 50147 66547 50175
rect 66575 50147 66609 50175
rect 66637 50147 66671 50175
rect 66699 50147 75485 50175
rect 75513 50147 75547 50175
rect 75575 50147 75609 50175
rect 75637 50147 75671 50175
rect 75699 50147 84485 50175
rect 84513 50147 84547 50175
rect 84575 50147 84609 50175
rect 84637 50147 84671 50175
rect 84699 50147 120485 50175
rect 120513 50147 120547 50175
rect 120575 50147 120609 50175
rect 120637 50147 120671 50175
rect 120699 50147 129485 50175
rect 129513 50147 129547 50175
rect 129575 50147 129609 50175
rect 129637 50147 129671 50175
rect 129699 50147 138485 50175
rect 138513 50147 138547 50175
rect 138575 50147 138609 50175
rect 138637 50147 138671 50175
rect 138699 50147 147485 50175
rect 147513 50147 147547 50175
rect 147575 50147 147609 50175
rect 147637 50147 147671 50175
rect 147699 50147 156485 50175
rect 156513 50147 156547 50175
rect 156575 50147 156609 50175
rect 156637 50147 156671 50175
rect 156699 50147 165485 50175
rect 165513 50147 165547 50175
rect 165575 50147 165609 50175
rect 165637 50147 165671 50175
rect 165699 50147 174485 50175
rect 174513 50147 174547 50175
rect 174575 50147 174609 50175
rect 174637 50147 174671 50175
rect 174699 50147 183485 50175
rect 183513 50147 183547 50175
rect 183575 50147 183609 50175
rect 183637 50147 183671 50175
rect 183699 50147 192485 50175
rect 192513 50147 192547 50175
rect 192575 50147 192609 50175
rect 192637 50147 192671 50175
rect 192699 50147 201485 50175
rect 201513 50147 201547 50175
rect 201575 50147 201609 50175
rect 201637 50147 201671 50175
rect 201699 50147 210485 50175
rect 210513 50147 210547 50175
rect 210575 50147 210609 50175
rect 210637 50147 210671 50175
rect 210699 50147 219485 50175
rect 219513 50147 219547 50175
rect 219575 50147 219609 50175
rect 219637 50147 219671 50175
rect 219699 50147 228485 50175
rect 228513 50147 228547 50175
rect 228575 50147 228609 50175
rect 228637 50147 228671 50175
rect 228699 50147 237485 50175
rect 237513 50147 237547 50175
rect 237575 50147 237609 50175
rect 237637 50147 237671 50175
rect 237699 50147 246485 50175
rect 246513 50147 246547 50175
rect 246575 50147 246609 50175
rect 246637 50147 246671 50175
rect 246699 50147 255485 50175
rect 255513 50147 255547 50175
rect 255575 50147 255609 50175
rect 255637 50147 255671 50175
rect 255699 50147 264485 50175
rect 264513 50147 264547 50175
rect 264575 50147 264609 50175
rect 264637 50147 264671 50175
rect 264699 50147 273485 50175
rect 273513 50147 273547 50175
rect 273575 50147 273609 50175
rect 273637 50147 273671 50175
rect 273699 50147 282485 50175
rect 282513 50147 282547 50175
rect 282575 50147 282609 50175
rect 282637 50147 282671 50175
rect 282699 50147 291485 50175
rect 291513 50147 291547 50175
rect 291575 50147 291609 50175
rect 291637 50147 291671 50175
rect 291699 50147 298728 50175
rect 298756 50147 298790 50175
rect 298818 50147 298852 50175
rect 298880 50147 298914 50175
rect 298942 50147 298990 50175
rect -958 50113 298990 50147
rect -958 50085 -910 50113
rect -882 50085 -848 50113
rect -820 50085 -786 50113
rect -758 50085 -724 50113
rect -696 50085 3485 50113
rect 3513 50085 3547 50113
rect 3575 50085 3609 50113
rect 3637 50085 3671 50113
rect 3699 50085 12485 50113
rect 12513 50085 12547 50113
rect 12575 50085 12609 50113
rect 12637 50085 12671 50113
rect 12699 50085 21485 50113
rect 21513 50085 21547 50113
rect 21575 50085 21609 50113
rect 21637 50085 21671 50113
rect 21699 50085 30485 50113
rect 30513 50085 30547 50113
rect 30575 50085 30609 50113
rect 30637 50085 30671 50113
rect 30699 50085 39485 50113
rect 39513 50085 39547 50113
rect 39575 50085 39609 50113
rect 39637 50085 39671 50113
rect 39699 50085 48485 50113
rect 48513 50085 48547 50113
rect 48575 50085 48609 50113
rect 48637 50085 48671 50113
rect 48699 50085 57485 50113
rect 57513 50085 57547 50113
rect 57575 50085 57609 50113
rect 57637 50085 57671 50113
rect 57699 50085 66485 50113
rect 66513 50085 66547 50113
rect 66575 50085 66609 50113
rect 66637 50085 66671 50113
rect 66699 50085 75485 50113
rect 75513 50085 75547 50113
rect 75575 50085 75609 50113
rect 75637 50085 75671 50113
rect 75699 50085 84485 50113
rect 84513 50085 84547 50113
rect 84575 50085 84609 50113
rect 84637 50085 84671 50113
rect 84699 50085 120485 50113
rect 120513 50085 120547 50113
rect 120575 50085 120609 50113
rect 120637 50085 120671 50113
rect 120699 50085 129485 50113
rect 129513 50085 129547 50113
rect 129575 50085 129609 50113
rect 129637 50085 129671 50113
rect 129699 50085 138485 50113
rect 138513 50085 138547 50113
rect 138575 50085 138609 50113
rect 138637 50085 138671 50113
rect 138699 50085 147485 50113
rect 147513 50085 147547 50113
rect 147575 50085 147609 50113
rect 147637 50085 147671 50113
rect 147699 50085 156485 50113
rect 156513 50085 156547 50113
rect 156575 50085 156609 50113
rect 156637 50085 156671 50113
rect 156699 50085 165485 50113
rect 165513 50085 165547 50113
rect 165575 50085 165609 50113
rect 165637 50085 165671 50113
rect 165699 50085 174485 50113
rect 174513 50085 174547 50113
rect 174575 50085 174609 50113
rect 174637 50085 174671 50113
rect 174699 50085 183485 50113
rect 183513 50085 183547 50113
rect 183575 50085 183609 50113
rect 183637 50085 183671 50113
rect 183699 50085 192485 50113
rect 192513 50085 192547 50113
rect 192575 50085 192609 50113
rect 192637 50085 192671 50113
rect 192699 50085 201485 50113
rect 201513 50085 201547 50113
rect 201575 50085 201609 50113
rect 201637 50085 201671 50113
rect 201699 50085 210485 50113
rect 210513 50085 210547 50113
rect 210575 50085 210609 50113
rect 210637 50085 210671 50113
rect 210699 50085 219485 50113
rect 219513 50085 219547 50113
rect 219575 50085 219609 50113
rect 219637 50085 219671 50113
rect 219699 50085 228485 50113
rect 228513 50085 228547 50113
rect 228575 50085 228609 50113
rect 228637 50085 228671 50113
rect 228699 50085 237485 50113
rect 237513 50085 237547 50113
rect 237575 50085 237609 50113
rect 237637 50085 237671 50113
rect 237699 50085 246485 50113
rect 246513 50085 246547 50113
rect 246575 50085 246609 50113
rect 246637 50085 246671 50113
rect 246699 50085 255485 50113
rect 255513 50085 255547 50113
rect 255575 50085 255609 50113
rect 255637 50085 255671 50113
rect 255699 50085 264485 50113
rect 264513 50085 264547 50113
rect 264575 50085 264609 50113
rect 264637 50085 264671 50113
rect 264699 50085 273485 50113
rect 273513 50085 273547 50113
rect 273575 50085 273609 50113
rect 273637 50085 273671 50113
rect 273699 50085 282485 50113
rect 282513 50085 282547 50113
rect 282575 50085 282609 50113
rect 282637 50085 282671 50113
rect 282699 50085 291485 50113
rect 291513 50085 291547 50113
rect 291575 50085 291609 50113
rect 291637 50085 291671 50113
rect 291699 50085 298728 50113
rect 298756 50085 298790 50113
rect 298818 50085 298852 50113
rect 298880 50085 298914 50113
rect 298942 50085 298990 50113
rect -958 50051 298990 50085
rect -958 50023 -910 50051
rect -882 50023 -848 50051
rect -820 50023 -786 50051
rect -758 50023 -724 50051
rect -696 50023 3485 50051
rect 3513 50023 3547 50051
rect 3575 50023 3609 50051
rect 3637 50023 3671 50051
rect 3699 50023 12485 50051
rect 12513 50023 12547 50051
rect 12575 50023 12609 50051
rect 12637 50023 12671 50051
rect 12699 50023 21485 50051
rect 21513 50023 21547 50051
rect 21575 50023 21609 50051
rect 21637 50023 21671 50051
rect 21699 50023 30485 50051
rect 30513 50023 30547 50051
rect 30575 50023 30609 50051
rect 30637 50023 30671 50051
rect 30699 50023 39485 50051
rect 39513 50023 39547 50051
rect 39575 50023 39609 50051
rect 39637 50023 39671 50051
rect 39699 50023 48485 50051
rect 48513 50023 48547 50051
rect 48575 50023 48609 50051
rect 48637 50023 48671 50051
rect 48699 50023 57485 50051
rect 57513 50023 57547 50051
rect 57575 50023 57609 50051
rect 57637 50023 57671 50051
rect 57699 50023 66485 50051
rect 66513 50023 66547 50051
rect 66575 50023 66609 50051
rect 66637 50023 66671 50051
rect 66699 50023 75485 50051
rect 75513 50023 75547 50051
rect 75575 50023 75609 50051
rect 75637 50023 75671 50051
rect 75699 50023 84485 50051
rect 84513 50023 84547 50051
rect 84575 50023 84609 50051
rect 84637 50023 84671 50051
rect 84699 50023 120485 50051
rect 120513 50023 120547 50051
rect 120575 50023 120609 50051
rect 120637 50023 120671 50051
rect 120699 50023 129485 50051
rect 129513 50023 129547 50051
rect 129575 50023 129609 50051
rect 129637 50023 129671 50051
rect 129699 50023 138485 50051
rect 138513 50023 138547 50051
rect 138575 50023 138609 50051
rect 138637 50023 138671 50051
rect 138699 50023 147485 50051
rect 147513 50023 147547 50051
rect 147575 50023 147609 50051
rect 147637 50023 147671 50051
rect 147699 50023 156485 50051
rect 156513 50023 156547 50051
rect 156575 50023 156609 50051
rect 156637 50023 156671 50051
rect 156699 50023 165485 50051
rect 165513 50023 165547 50051
rect 165575 50023 165609 50051
rect 165637 50023 165671 50051
rect 165699 50023 174485 50051
rect 174513 50023 174547 50051
rect 174575 50023 174609 50051
rect 174637 50023 174671 50051
rect 174699 50023 183485 50051
rect 183513 50023 183547 50051
rect 183575 50023 183609 50051
rect 183637 50023 183671 50051
rect 183699 50023 192485 50051
rect 192513 50023 192547 50051
rect 192575 50023 192609 50051
rect 192637 50023 192671 50051
rect 192699 50023 201485 50051
rect 201513 50023 201547 50051
rect 201575 50023 201609 50051
rect 201637 50023 201671 50051
rect 201699 50023 210485 50051
rect 210513 50023 210547 50051
rect 210575 50023 210609 50051
rect 210637 50023 210671 50051
rect 210699 50023 219485 50051
rect 219513 50023 219547 50051
rect 219575 50023 219609 50051
rect 219637 50023 219671 50051
rect 219699 50023 228485 50051
rect 228513 50023 228547 50051
rect 228575 50023 228609 50051
rect 228637 50023 228671 50051
rect 228699 50023 237485 50051
rect 237513 50023 237547 50051
rect 237575 50023 237609 50051
rect 237637 50023 237671 50051
rect 237699 50023 246485 50051
rect 246513 50023 246547 50051
rect 246575 50023 246609 50051
rect 246637 50023 246671 50051
rect 246699 50023 255485 50051
rect 255513 50023 255547 50051
rect 255575 50023 255609 50051
rect 255637 50023 255671 50051
rect 255699 50023 264485 50051
rect 264513 50023 264547 50051
rect 264575 50023 264609 50051
rect 264637 50023 264671 50051
rect 264699 50023 273485 50051
rect 273513 50023 273547 50051
rect 273575 50023 273609 50051
rect 273637 50023 273671 50051
rect 273699 50023 282485 50051
rect 282513 50023 282547 50051
rect 282575 50023 282609 50051
rect 282637 50023 282671 50051
rect 282699 50023 291485 50051
rect 291513 50023 291547 50051
rect 291575 50023 291609 50051
rect 291637 50023 291671 50051
rect 291699 50023 298728 50051
rect 298756 50023 298790 50051
rect 298818 50023 298852 50051
rect 298880 50023 298914 50051
rect 298942 50023 298990 50051
rect -958 49989 298990 50023
rect -958 49961 -910 49989
rect -882 49961 -848 49989
rect -820 49961 -786 49989
rect -758 49961 -724 49989
rect -696 49961 3485 49989
rect 3513 49961 3547 49989
rect 3575 49961 3609 49989
rect 3637 49961 3671 49989
rect 3699 49961 12485 49989
rect 12513 49961 12547 49989
rect 12575 49961 12609 49989
rect 12637 49961 12671 49989
rect 12699 49961 21485 49989
rect 21513 49961 21547 49989
rect 21575 49961 21609 49989
rect 21637 49961 21671 49989
rect 21699 49961 30485 49989
rect 30513 49961 30547 49989
rect 30575 49961 30609 49989
rect 30637 49961 30671 49989
rect 30699 49961 39485 49989
rect 39513 49961 39547 49989
rect 39575 49961 39609 49989
rect 39637 49961 39671 49989
rect 39699 49961 48485 49989
rect 48513 49961 48547 49989
rect 48575 49961 48609 49989
rect 48637 49961 48671 49989
rect 48699 49961 57485 49989
rect 57513 49961 57547 49989
rect 57575 49961 57609 49989
rect 57637 49961 57671 49989
rect 57699 49961 66485 49989
rect 66513 49961 66547 49989
rect 66575 49961 66609 49989
rect 66637 49961 66671 49989
rect 66699 49961 75485 49989
rect 75513 49961 75547 49989
rect 75575 49961 75609 49989
rect 75637 49961 75671 49989
rect 75699 49961 84485 49989
rect 84513 49961 84547 49989
rect 84575 49961 84609 49989
rect 84637 49961 84671 49989
rect 84699 49961 120485 49989
rect 120513 49961 120547 49989
rect 120575 49961 120609 49989
rect 120637 49961 120671 49989
rect 120699 49961 129485 49989
rect 129513 49961 129547 49989
rect 129575 49961 129609 49989
rect 129637 49961 129671 49989
rect 129699 49961 138485 49989
rect 138513 49961 138547 49989
rect 138575 49961 138609 49989
rect 138637 49961 138671 49989
rect 138699 49961 147485 49989
rect 147513 49961 147547 49989
rect 147575 49961 147609 49989
rect 147637 49961 147671 49989
rect 147699 49961 156485 49989
rect 156513 49961 156547 49989
rect 156575 49961 156609 49989
rect 156637 49961 156671 49989
rect 156699 49961 165485 49989
rect 165513 49961 165547 49989
rect 165575 49961 165609 49989
rect 165637 49961 165671 49989
rect 165699 49961 174485 49989
rect 174513 49961 174547 49989
rect 174575 49961 174609 49989
rect 174637 49961 174671 49989
rect 174699 49961 183485 49989
rect 183513 49961 183547 49989
rect 183575 49961 183609 49989
rect 183637 49961 183671 49989
rect 183699 49961 192485 49989
rect 192513 49961 192547 49989
rect 192575 49961 192609 49989
rect 192637 49961 192671 49989
rect 192699 49961 201485 49989
rect 201513 49961 201547 49989
rect 201575 49961 201609 49989
rect 201637 49961 201671 49989
rect 201699 49961 210485 49989
rect 210513 49961 210547 49989
rect 210575 49961 210609 49989
rect 210637 49961 210671 49989
rect 210699 49961 219485 49989
rect 219513 49961 219547 49989
rect 219575 49961 219609 49989
rect 219637 49961 219671 49989
rect 219699 49961 228485 49989
rect 228513 49961 228547 49989
rect 228575 49961 228609 49989
rect 228637 49961 228671 49989
rect 228699 49961 237485 49989
rect 237513 49961 237547 49989
rect 237575 49961 237609 49989
rect 237637 49961 237671 49989
rect 237699 49961 246485 49989
rect 246513 49961 246547 49989
rect 246575 49961 246609 49989
rect 246637 49961 246671 49989
rect 246699 49961 255485 49989
rect 255513 49961 255547 49989
rect 255575 49961 255609 49989
rect 255637 49961 255671 49989
rect 255699 49961 264485 49989
rect 264513 49961 264547 49989
rect 264575 49961 264609 49989
rect 264637 49961 264671 49989
rect 264699 49961 273485 49989
rect 273513 49961 273547 49989
rect 273575 49961 273609 49989
rect 273637 49961 273671 49989
rect 273699 49961 282485 49989
rect 282513 49961 282547 49989
rect 282575 49961 282609 49989
rect 282637 49961 282671 49989
rect 282699 49961 291485 49989
rect 291513 49961 291547 49989
rect 291575 49961 291609 49989
rect 291637 49961 291671 49989
rect 291699 49961 298728 49989
rect 298756 49961 298790 49989
rect 298818 49961 298852 49989
rect 298880 49961 298914 49989
rect 298942 49961 298990 49989
rect -958 49913 298990 49961
rect -958 47175 298990 47223
rect -958 47147 -430 47175
rect -402 47147 -368 47175
rect -340 47147 -306 47175
rect -278 47147 -244 47175
rect -216 47147 1625 47175
rect 1653 47147 1687 47175
rect 1715 47147 1749 47175
rect 1777 47147 1811 47175
rect 1839 47147 10625 47175
rect 10653 47147 10687 47175
rect 10715 47147 10749 47175
rect 10777 47147 10811 47175
rect 10839 47147 19625 47175
rect 19653 47147 19687 47175
rect 19715 47147 19749 47175
rect 19777 47147 19811 47175
rect 19839 47147 28625 47175
rect 28653 47147 28687 47175
rect 28715 47147 28749 47175
rect 28777 47147 28811 47175
rect 28839 47147 37625 47175
rect 37653 47147 37687 47175
rect 37715 47147 37749 47175
rect 37777 47147 37811 47175
rect 37839 47147 46625 47175
rect 46653 47147 46687 47175
rect 46715 47147 46749 47175
rect 46777 47147 46811 47175
rect 46839 47147 55625 47175
rect 55653 47147 55687 47175
rect 55715 47147 55749 47175
rect 55777 47147 55811 47175
rect 55839 47147 64625 47175
rect 64653 47147 64687 47175
rect 64715 47147 64749 47175
rect 64777 47147 64811 47175
rect 64839 47147 73625 47175
rect 73653 47147 73687 47175
rect 73715 47147 73749 47175
rect 73777 47147 73811 47175
rect 73839 47147 82625 47175
rect 82653 47147 82687 47175
rect 82715 47147 82749 47175
rect 82777 47147 82811 47175
rect 82839 47147 91625 47175
rect 91653 47147 91687 47175
rect 91715 47147 91749 47175
rect 91777 47147 91811 47175
rect 91839 47147 100625 47175
rect 100653 47147 100687 47175
rect 100715 47147 100749 47175
rect 100777 47147 100811 47175
rect 100839 47147 109625 47175
rect 109653 47147 109687 47175
rect 109715 47147 109749 47175
rect 109777 47147 109811 47175
rect 109839 47147 118625 47175
rect 118653 47147 118687 47175
rect 118715 47147 118749 47175
rect 118777 47147 118811 47175
rect 118839 47147 127625 47175
rect 127653 47147 127687 47175
rect 127715 47147 127749 47175
rect 127777 47147 127811 47175
rect 127839 47147 136625 47175
rect 136653 47147 136687 47175
rect 136715 47147 136749 47175
rect 136777 47147 136811 47175
rect 136839 47147 145625 47175
rect 145653 47147 145687 47175
rect 145715 47147 145749 47175
rect 145777 47147 145811 47175
rect 145839 47147 154625 47175
rect 154653 47147 154687 47175
rect 154715 47147 154749 47175
rect 154777 47147 154811 47175
rect 154839 47147 163625 47175
rect 163653 47147 163687 47175
rect 163715 47147 163749 47175
rect 163777 47147 163811 47175
rect 163839 47147 172625 47175
rect 172653 47147 172687 47175
rect 172715 47147 172749 47175
rect 172777 47147 172811 47175
rect 172839 47147 181625 47175
rect 181653 47147 181687 47175
rect 181715 47147 181749 47175
rect 181777 47147 181811 47175
rect 181839 47147 190625 47175
rect 190653 47147 190687 47175
rect 190715 47147 190749 47175
rect 190777 47147 190811 47175
rect 190839 47147 199625 47175
rect 199653 47147 199687 47175
rect 199715 47147 199749 47175
rect 199777 47147 199811 47175
rect 199839 47147 208625 47175
rect 208653 47147 208687 47175
rect 208715 47147 208749 47175
rect 208777 47147 208811 47175
rect 208839 47147 217625 47175
rect 217653 47147 217687 47175
rect 217715 47147 217749 47175
rect 217777 47147 217811 47175
rect 217839 47147 226625 47175
rect 226653 47147 226687 47175
rect 226715 47147 226749 47175
rect 226777 47147 226811 47175
rect 226839 47147 235625 47175
rect 235653 47147 235687 47175
rect 235715 47147 235749 47175
rect 235777 47147 235811 47175
rect 235839 47147 244625 47175
rect 244653 47147 244687 47175
rect 244715 47147 244749 47175
rect 244777 47147 244811 47175
rect 244839 47147 253625 47175
rect 253653 47147 253687 47175
rect 253715 47147 253749 47175
rect 253777 47147 253811 47175
rect 253839 47147 262625 47175
rect 262653 47147 262687 47175
rect 262715 47147 262749 47175
rect 262777 47147 262811 47175
rect 262839 47147 271625 47175
rect 271653 47147 271687 47175
rect 271715 47147 271749 47175
rect 271777 47147 271811 47175
rect 271839 47147 280625 47175
rect 280653 47147 280687 47175
rect 280715 47147 280749 47175
rect 280777 47147 280811 47175
rect 280839 47147 289625 47175
rect 289653 47147 289687 47175
rect 289715 47147 289749 47175
rect 289777 47147 289811 47175
rect 289839 47147 298248 47175
rect 298276 47147 298310 47175
rect 298338 47147 298372 47175
rect 298400 47147 298434 47175
rect 298462 47147 298990 47175
rect -958 47113 298990 47147
rect -958 47085 -430 47113
rect -402 47085 -368 47113
rect -340 47085 -306 47113
rect -278 47085 -244 47113
rect -216 47085 1625 47113
rect 1653 47085 1687 47113
rect 1715 47085 1749 47113
rect 1777 47085 1811 47113
rect 1839 47085 10625 47113
rect 10653 47085 10687 47113
rect 10715 47085 10749 47113
rect 10777 47085 10811 47113
rect 10839 47085 19625 47113
rect 19653 47085 19687 47113
rect 19715 47085 19749 47113
rect 19777 47085 19811 47113
rect 19839 47085 28625 47113
rect 28653 47085 28687 47113
rect 28715 47085 28749 47113
rect 28777 47085 28811 47113
rect 28839 47085 37625 47113
rect 37653 47085 37687 47113
rect 37715 47085 37749 47113
rect 37777 47085 37811 47113
rect 37839 47085 46625 47113
rect 46653 47085 46687 47113
rect 46715 47085 46749 47113
rect 46777 47085 46811 47113
rect 46839 47085 55625 47113
rect 55653 47085 55687 47113
rect 55715 47085 55749 47113
rect 55777 47085 55811 47113
rect 55839 47085 64625 47113
rect 64653 47085 64687 47113
rect 64715 47085 64749 47113
rect 64777 47085 64811 47113
rect 64839 47085 73625 47113
rect 73653 47085 73687 47113
rect 73715 47085 73749 47113
rect 73777 47085 73811 47113
rect 73839 47085 82625 47113
rect 82653 47085 82687 47113
rect 82715 47085 82749 47113
rect 82777 47085 82811 47113
rect 82839 47085 91625 47113
rect 91653 47085 91687 47113
rect 91715 47085 91749 47113
rect 91777 47085 91811 47113
rect 91839 47085 100625 47113
rect 100653 47085 100687 47113
rect 100715 47085 100749 47113
rect 100777 47085 100811 47113
rect 100839 47085 109625 47113
rect 109653 47085 109687 47113
rect 109715 47085 109749 47113
rect 109777 47085 109811 47113
rect 109839 47085 118625 47113
rect 118653 47085 118687 47113
rect 118715 47085 118749 47113
rect 118777 47085 118811 47113
rect 118839 47085 127625 47113
rect 127653 47085 127687 47113
rect 127715 47085 127749 47113
rect 127777 47085 127811 47113
rect 127839 47085 136625 47113
rect 136653 47085 136687 47113
rect 136715 47085 136749 47113
rect 136777 47085 136811 47113
rect 136839 47085 145625 47113
rect 145653 47085 145687 47113
rect 145715 47085 145749 47113
rect 145777 47085 145811 47113
rect 145839 47085 154625 47113
rect 154653 47085 154687 47113
rect 154715 47085 154749 47113
rect 154777 47085 154811 47113
rect 154839 47085 163625 47113
rect 163653 47085 163687 47113
rect 163715 47085 163749 47113
rect 163777 47085 163811 47113
rect 163839 47085 172625 47113
rect 172653 47085 172687 47113
rect 172715 47085 172749 47113
rect 172777 47085 172811 47113
rect 172839 47085 181625 47113
rect 181653 47085 181687 47113
rect 181715 47085 181749 47113
rect 181777 47085 181811 47113
rect 181839 47085 190625 47113
rect 190653 47085 190687 47113
rect 190715 47085 190749 47113
rect 190777 47085 190811 47113
rect 190839 47085 199625 47113
rect 199653 47085 199687 47113
rect 199715 47085 199749 47113
rect 199777 47085 199811 47113
rect 199839 47085 208625 47113
rect 208653 47085 208687 47113
rect 208715 47085 208749 47113
rect 208777 47085 208811 47113
rect 208839 47085 217625 47113
rect 217653 47085 217687 47113
rect 217715 47085 217749 47113
rect 217777 47085 217811 47113
rect 217839 47085 226625 47113
rect 226653 47085 226687 47113
rect 226715 47085 226749 47113
rect 226777 47085 226811 47113
rect 226839 47085 235625 47113
rect 235653 47085 235687 47113
rect 235715 47085 235749 47113
rect 235777 47085 235811 47113
rect 235839 47085 244625 47113
rect 244653 47085 244687 47113
rect 244715 47085 244749 47113
rect 244777 47085 244811 47113
rect 244839 47085 253625 47113
rect 253653 47085 253687 47113
rect 253715 47085 253749 47113
rect 253777 47085 253811 47113
rect 253839 47085 262625 47113
rect 262653 47085 262687 47113
rect 262715 47085 262749 47113
rect 262777 47085 262811 47113
rect 262839 47085 271625 47113
rect 271653 47085 271687 47113
rect 271715 47085 271749 47113
rect 271777 47085 271811 47113
rect 271839 47085 280625 47113
rect 280653 47085 280687 47113
rect 280715 47085 280749 47113
rect 280777 47085 280811 47113
rect 280839 47085 289625 47113
rect 289653 47085 289687 47113
rect 289715 47085 289749 47113
rect 289777 47085 289811 47113
rect 289839 47085 298248 47113
rect 298276 47085 298310 47113
rect 298338 47085 298372 47113
rect 298400 47085 298434 47113
rect 298462 47085 298990 47113
rect -958 47051 298990 47085
rect -958 47023 -430 47051
rect -402 47023 -368 47051
rect -340 47023 -306 47051
rect -278 47023 -244 47051
rect -216 47023 1625 47051
rect 1653 47023 1687 47051
rect 1715 47023 1749 47051
rect 1777 47023 1811 47051
rect 1839 47023 10625 47051
rect 10653 47023 10687 47051
rect 10715 47023 10749 47051
rect 10777 47023 10811 47051
rect 10839 47023 19625 47051
rect 19653 47023 19687 47051
rect 19715 47023 19749 47051
rect 19777 47023 19811 47051
rect 19839 47023 28625 47051
rect 28653 47023 28687 47051
rect 28715 47023 28749 47051
rect 28777 47023 28811 47051
rect 28839 47023 37625 47051
rect 37653 47023 37687 47051
rect 37715 47023 37749 47051
rect 37777 47023 37811 47051
rect 37839 47023 46625 47051
rect 46653 47023 46687 47051
rect 46715 47023 46749 47051
rect 46777 47023 46811 47051
rect 46839 47023 55625 47051
rect 55653 47023 55687 47051
rect 55715 47023 55749 47051
rect 55777 47023 55811 47051
rect 55839 47023 64625 47051
rect 64653 47023 64687 47051
rect 64715 47023 64749 47051
rect 64777 47023 64811 47051
rect 64839 47023 73625 47051
rect 73653 47023 73687 47051
rect 73715 47023 73749 47051
rect 73777 47023 73811 47051
rect 73839 47023 82625 47051
rect 82653 47023 82687 47051
rect 82715 47023 82749 47051
rect 82777 47023 82811 47051
rect 82839 47023 91625 47051
rect 91653 47023 91687 47051
rect 91715 47023 91749 47051
rect 91777 47023 91811 47051
rect 91839 47023 100625 47051
rect 100653 47023 100687 47051
rect 100715 47023 100749 47051
rect 100777 47023 100811 47051
rect 100839 47023 109625 47051
rect 109653 47023 109687 47051
rect 109715 47023 109749 47051
rect 109777 47023 109811 47051
rect 109839 47023 118625 47051
rect 118653 47023 118687 47051
rect 118715 47023 118749 47051
rect 118777 47023 118811 47051
rect 118839 47023 127625 47051
rect 127653 47023 127687 47051
rect 127715 47023 127749 47051
rect 127777 47023 127811 47051
rect 127839 47023 136625 47051
rect 136653 47023 136687 47051
rect 136715 47023 136749 47051
rect 136777 47023 136811 47051
rect 136839 47023 145625 47051
rect 145653 47023 145687 47051
rect 145715 47023 145749 47051
rect 145777 47023 145811 47051
rect 145839 47023 154625 47051
rect 154653 47023 154687 47051
rect 154715 47023 154749 47051
rect 154777 47023 154811 47051
rect 154839 47023 163625 47051
rect 163653 47023 163687 47051
rect 163715 47023 163749 47051
rect 163777 47023 163811 47051
rect 163839 47023 172625 47051
rect 172653 47023 172687 47051
rect 172715 47023 172749 47051
rect 172777 47023 172811 47051
rect 172839 47023 181625 47051
rect 181653 47023 181687 47051
rect 181715 47023 181749 47051
rect 181777 47023 181811 47051
rect 181839 47023 190625 47051
rect 190653 47023 190687 47051
rect 190715 47023 190749 47051
rect 190777 47023 190811 47051
rect 190839 47023 199625 47051
rect 199653 47023 199687 47051
rect 199715 47023 199749 47051
rect 199777 47023 199811 47051
rect 199839 47023 208625 47051
rect 208653 47023 208687 47051
rect 208715 47023 208749 47051
rect 208777 47023 208811 47051
rect 208839 47023 217625 47051
rect 217653 47023 217687 47051
rect 217715 47023 217749 47051
rect 217777 47023 217811 47051
rect 217839 47023 226625 47051
rect 226653 47023 226687 47051
rect 226715 47023 226749 47051
rect 226777 47023 226811 47051
rect 226839 47023 235625 47051
rect 235653 47023 235687 47051
rect 235715 47023 235749 47051
rect 235777 47023 235811 47051
rect 235839 47023 244625 47051
rect 244653 47023 244687 47051
rect 244715 47023 244749 47051
rect 244777 47023 244811 47051
rect 244839 47023 253625 47051
rect 253653 47023 253687 47051
rect 253715 47023 253749 47051
rect 253777 47023 253811 47051
rect 253839 47023 262625 47051
rect 262653 47023 262687 47051
rect 262715 47023 262749 47051
rect 262777 47023 262811 47051
rect 262839 47023 271625 47051
rect 271653 47023 271687 47051
rect 271715 47023 271749 47051
rect 271777 47023 271811 47051
rect 271839 47023 280625 47051
rect 280653 47023 280687 47051
rect 280715 47023 280749 47051
rect 280777 47023 280811 47051
rect 280839 47023 289625 47051
rect 289653 47023 289687 47051
rect 289715 47023 289749 47051
rect 289777 47023 289811 47051
rect 289839 47023 298248 47051
rect 298276 47023 298310 47051
rect 298338 47023 298372 47051
rect 298400 47023 298434 47051
rect 298462 47023 298990 47051
rect -958 46989 298990 47023
rect -958 46961 -430 46989
rect -402 46961 -368 46989
rect -340 46961 -306 46989
rect -278 46961 -244 46989
rect -216 46961 1625 46989
rect 1653 46961 1687 46989
rect 1715 46961 1749 46989
rect 1777 46961 1811 46989
rect 1839 46961 10625 46989
rect 10653 46961 10687 46989
rect 10715 46961 10749 46989
rect 10777 46961 10811 46989
rect 10839 46961 19625 46989
rect 19653 46961 19687 46989
rect 19715 46961 19749 46989
rect 19777 46961 19811 46989
rect 19839 46961 28625 46989
rect 28653 46961 28687 46989
rect 28715 46961 28749 46989
rect 28777 46961 28811 46989
rect 28839 46961 37625 46989
rect 37653 46961 37687 46989
rect 37715 46961 37749 46989
rect 37777 46961 37811 46989
rect 37839 46961 46625 46989
rect 46653 46961 46687 46989
rect 46715 46961 46749 46989
rect 46777 46961 46811 46989
rect 46839 46961 55625 46989
rect 55653 46961 55687 46989
rect 55715 46961 55749 46989
rect 55777 46961 55811 46989
rect 55839 46961 64625 46989
rect 64653 46961 64687 46989
rect 64715 46961 64749 46989
rect 64777 46961 64811 46989
rect 64839 46961 73625 46989
rect 73653 46961 73687 46989
rect 73715 46961 73749 46989
rect 73777 46961 73811 46989
rect 73839 46961 82625 46989
rect 82653 46961 82687 46989
rect 82715 46961 82749 46989
rect 82777 46961 82811 46989
rect 82839 46961 91625 46989
rect 91653 46961 91687 46989
rect 91715 46961 91749 46989
rect 91777 46961 91811 46989
rect 91839 46961 100625 46989
rect 100653 46961 100687 46989
rect 100715 46961 100749 46989
rect 100777 46961 100811 46989
rect 100839 46961 109625 46989
rect 109653 46961 109687 46989
rect 109715 46961 109749 46989
rect 109777 46961 109811 46989
rect 109839 46961 118625 46989
rect 118653 46961 118687 46989
rect 118715 46961 118749 46989
rect 118777 46961 118811 46989
rect 118839 46961 127625 46989
rect 127653 46961 127687 46989
rect 127715 46961 127749 46989
rect 127777 46961 127811 46989
rect 127839 46961 136625 46989
rect 136653 46961 136687 46989
rect 136715 46961 136749 46989
rect 136777 46961 136811 46989
rect 136839 46961 145625 46989
rect 145653 46961 145687 46989
rect 145715 46961 145749 46989
rect 145777 46961 145811 46989
rect 145839 46961 154625 46989
rect 154653 46961 154687 46989
rect 154715 46961 154749 46989
rect 154777 46961 154811 46989
rect 154839 46961 163625 46989
rect 163653 46961 163687 46989
rect 163715 46961 163749 46989
rect 163777 46961 163811 46989
rect 163839 46961 172625 46989
rect 172653 46961 172687 46989
rect 172715 46961 172749 46989
rect 172777 46961 172811 46989
rect 172839 46961 181625 46989
rect 181653 46961 181687 46989
rect 181715 46961 181749 46989
rect 181777 46961 181811 46989
rect 181839 46961 190625 46989
rect 190653 46961 190687 46989
rect 190715 46961 190749 46989
rect 190777 46961 190811 46989
rect 190839 46961 199625 46989
rect 199653 46961 199687 46989
rect 199715 46961 199749 46989
rect 199777 46961 199811 46989
rect 199839 46961 208625 46989
rect 208653 46961 208687 46989
rect 208715 46961 208749 46989
rect 208777 46961 208811 46989
rect 208839 46961 217625 46989
rect 217653 46961 217687 46989
rect 217715 46961 217749 46989
rect 217777 46961 217811 46989
rect 217839 46961 226625 46989
rect 226653 46961 226687 46989
rect 226715 46961 226749 46989
rect 226777 46961 226811 46989
rect 226839 46961 235625 46989
rect 235653 46961 235687 46989
rect 235715 46961 235749 46989
rect 235777 46961 235811 46989
rect 235839 46961 244625 46989
rect 244653 46961 244687 46989
rect 244715 46961 244749 46989
rect 244777 46961 244811 46989
rect 244839 46961 253625 46989
rect 253653 46961 253687 46989
rect 253715 46961 253749 46989
rect 253777 46961 253811 46989
rect 253839 46961 262625 46989
rect 262653 46961 262687 46989
rect 262715 46961 262749 46989
rect 262777 46961 262811 46989
rect 262839 46961 271625 46989
rect 271653 46961 271687 46989
rect 271715 46961 271749 46989
rect 271777 46961 271811 46989
rect 271839 46961 280625 46989
rect 280653 46961 280687 46989
rect 280715 46961 280749 46989
rect 280777 46961 280811 46989
rect 280839 46961 289625 46989
rect 289653 46961 289687 46989
rect 289715 46961 289749 46989
rect 289777 46961 289811 46989
rect 289839 46961 298248 46989
rect 298276 46961 298310 46989
rect 298338 46961 298372 46989
rect 298400 46961 298434 46989
rect 298462 46961 298990 46989
rect -958 46913 298990 46961
rect -958 41175 298990 41223
rect -958 41147 -910 41175
rect -882 41147 -848 41175
rect -820 41147 -786 41175
rect -758 41147 -724 41175
rect -696 41147 3485 41175
rect 3513 41147 3547 41175
rect 3575 41147 3609 41175
rect 3637 41147 3671 41175
rect 3699 41147 12485 41175
rect 12513 41147 12547 41175
rect 12575 41147 12609 41175
rect 12637 41147 12671 41175
rect 12699 41147 21485 41175
rect 21513 41147 21547 41175
rect 21575 41147 21609 41175
rect 21637 41147 21671 41175
rect 21699 41147 30485 41175
rect 30513 41147 30547 41175
rect 30575 41147 30609 41175
rect 30637 41147 30671 41175
rect 30699 41147 39485 41175
rect 39513 41147 39547 41175
rect 39575 41147 39609 41175
rect 39637 41147 39671 41175
rect 39699 41147 48485 41175
rect 48513 41147 48547 41175
rect 48575 41147 48609 41175
rect 48637 41147 48671 41175
rect 48699 41147 57485 41175
rect 57513 41147 57547 41175
rect 57575 41147 57609 41175
rect 57637 41147 57671 41175
rect 57699 41147 66485 41175
rect 66513 41147 66547 41175
rect 66575 41147 66609 41175
rect 66637 41147 66671 41175
rect 66699 41147 75485 41175
rect 75513 41147 75547 41175
rect 75575 41147 75609 41175
rect 75637 41147 75671 41175
rect 75699 41147 84485 41175
rect 84513 41147 84547 41175
rect 84575 41147 84609 41175
rect 84637 41147 84671 41175
rect 84699 41147 93485 41175
rect 93513 41147 93547 41175
rect 93575 41147 93609 41175
rect 93637 41147 93671 41175
rect 93699 41147 102485 41175
rect 102513 41147 102547 41175
rect 102575 41147 102609 41175
rect 102637 41147 102671 41175
rect 102699 41147 111485 41175
rect 111513 41147 111547 41175
rect 111575 41147 111609 41175
rect 111637 41147 111671 41175
rect 111699 41147 120485 41175
rect 120513 41147 120547 41175
rect 120575 41147 120609 41175
rect 120637 41147 120671 41175
rect 120699 41147 129485 41175
rect 129513 41147 129547 41175
rect 129575 41147 129609 41175
rect 129637 41147 129671 41175
rect 129699 41147 138485 41175
rect 138513 41147 138547 41175
rect 138575 41147 138609 41175
rect 138637 41147 138671 41175
rect 138699 41147 147485 41175
rect 147513 41147 147547 41175
rect 147575 41147 147609 41175
rect 147637 41147 147671 41175
rect 147699 41147 156485 41175
rect 156513 41147 156547 41175
rect 156575 41147 156609 41175
rect 156637 41147 156671 41175
rect 156699 41147 165485 41175
rect 165513 41147 165547 41175
rect 165575 41147 165609 41175
rect 165637 41147 165671 41175
rect 165699 41147 174485 41175
rect 174513 41147 174547 41175
rect 174575 41147 174609 41175
rect 174637 41147 174671 41175
rect 174699 41147 183485 41175
rect 183513 41147 183547 41175
rect 183575 41147 183609 41175
rect 183637 41147 183671 41175
rect 183699 41147 192485 41175
rect 192513 41147 192547 41175
rect 192575 41147 192609 41175
rect 192637 41147 192671 41175
rect 192699 41147 201485 41175
rect 201513 41147 201547 41175
rect 201575 41147 201609 41175
rect 201637 41147 201671 41175
rect 201699 41147 210485 41175
rect 210513 41147 210547 41175
rect 210575 41147 210609 41175
rect 210637 41147 210671 41175
rect 210699 41147 219485 41175
rect 219513 41147 219547 41175
rect 219575 41147 219609 41175
rect 219637 41147 219671 41175
rect 219699 41147 228485 41175
rect 228513 41147 228547 41175
rect 228575 41147 228609 41175
rect 228637 41147 228671 41175
rect 228699 41147 237485 41175
rect 237513 41147 237547 41175
rect 237575 41147 237609 41175
rect 237637 41147 237671 41175
rect 237699 41147 246485 41175
rect 246513 41147 246547 41175
rect 246575 41147 246609 41175
rect 246637 41147 246671 41175
rect 246699 41147 255485 41175
rect 255513 41147 255547 41175
rect 255575 41147 255609 41175
rect 255637 41147 255671 41175
rect 255699 41147 264485 41175
rect 264513 41147 264547 41175
rect 264575 41147 264609 41175
rect 264637 41147 264671 41175
rect 264699 41147 273485 41175
rect 273513 41147 273547 41175
rect 273575 41147 273609 41175
rect 273637 41147 273671 41175
rect 273699 41147 282485 41175
rect 282513 41147 282547 41175
rect 282575 41147 282609 41175
rect 282637 41147 282671 41175
rect 282699 41147 291485 41175
rect 291513 41147 291547 41175
rect 291575 41147 291609 41175
rect 291637 41147 291671 41175
rect 291699 41147 298728 41175
rect 298756 41147 298790 41175
rect 298818 41147 298852 41175
rect 298880 41147 298914 41175
rect 298942 41147 298990 41175
rect -958 41113 298990 41147
rect -958 41085 -910 41113
rect -882 41085 -848 41113
rect -820 41085 -786 41113
rect -758 41085 -724 41113
rect -696 41085 3485 41113
rect 3513 41085 3547 41113
rect 3575 41085 3609 41113
rect 3637 41085 3671 41113
rect 3699 41085 12485 41113
rect 12513 41085 12547 41113
rect 12575 41085 12609 41113
rect 12637 41085 12671 41113
rect 12699 41085 21485 41113
rect 21513 41085 21547 41113
rect 21575 41085 21609 41113
rect 21637 41085 21671 41113
rect 21699 41085 30485 41113
rect 30513 41085 30547 41113
rect 30575 41085 30609 41113
rect 30637 41085 30671 41113
rect 30699 41085 39485 41113
rect 39513 41085 39547 41113
rect 39575 41085 39609 41113
rect 39637 41085 39671 41113
rect 39699 41085 48485 41113
rect 48513 41085 48547 41113
rect 48575 41085 48609 41113
rect 48637 41085 48671 41113
rect 48699 41085 57485 41113
rect 57513 41085 57547 41113
rect 57575 41085 57609 41113
rect 57637 41085 57671 41113
rect 57699 41085 66485 41113
rect 66513 41085 66547 41113
rect 66575 41085 66609 41113
rect 66637 41085 66671 41113
rect 66699 41085 75485 41113
rect 75513 41085 75547 41113
rect 75575 41085 75609 41113
rect 75637 41085 75671 41113
rect 75699 41085 84485 41113
rect 84513 41085 84547 41113
rect 84575 41085 84609 41113
rect 84637 41085 84671 41113
rect 84699 41085 93485 41113
rect 93513 41085 93547 41113
rect 93575 41085 93609 41113
rect 93637 41085 93671 41113
rect 93699 41085 102485 41113
rect 102513 41085 102547 41113
rect 102575 41085 102609 41113
rect 102637 41085 102671 41113
rect 102699 41085 111485 41113
rect 111513 41085 111547 41113
rect 111575 41085 111609 41113
rect 111637 41085 111671 41113
rect 111699 41085 120485 41113
rect 120513 41085 120547 41113
rect 120575 41085 120609 41113
rect 120637 41085 120671 41113
rect 120699 41085 129485 41113
rect 129513 41085 129547 41113
rect 129575 41085 129609 41113
rect 129637 41085 129671 41113
rect 129699 41085 138485 41113
rect 138513 41085 138547 41113
rect 138575 41085 138609 41113
rect 138637 41085 138671 41113
rect 138699 41085 147485 41113
rect 147513 41085 147547 41113
rect 147575 41085 147609 41113
rect 147637 41085 147671 41113
rect 147699 41085 156485 41113
rect 156513 41085 156547 41113
rect 156575 41085 156609 41113
rect 156637 41085 156671 41113
rect 156699 41085 165485 41113
rect 165513 41085 165547 41113
rect 165575 41085 165609 41113
rect 165637 41085 165671 41113
rect 165699 41085 174485 41113
rect 174513 41085 174547 41113
rect 174575 41085 174609 41113
rect 174637 41085 174671 41113
rect 174699 41085 183485 41113
rect 183513 41085 183547 41113
rect 183575 41085 183609 41113
rect 183637 41085 183671 41113
rect 183699 41085 192485 41113
rect 192513 41085 192547 41113
rect 192575 41085 192609 41113
rect 192637 41085 192671 41113
rect 192699 41085 201485 41113
rect 201513 41085 201547 41113
rect 201575 41085 201609 41113
rect 201637 41085 201671 41113
rect 201699 41085 210485 41113
rect 210513 41085 210547 41113
rect 210575 41085 210609 41113
rect 210637 41085 210671 41113
rect 210699 41085 219485 41113
rect 219513 41085 219547 41113
rect 219575 41085 219609 41113
rect 219637 41085 219671 41113
rect 219699 41085 228485 41113
rect 228513 41085 228547 41113
rect 228575 41085 228609 41113
rect 228637 41085 228671 41113
rect 228699 41085 237485 41113
rect 237513 41085 237547 41113
rect 237575 41085 237609 41113
rect 237637 41085 237671 41113
rect 237699 41085 246485 41113
rect 246513 41085 246547 41113
rect 246575 41085 246609 41113
rect 246637 41085 246671 41113
rect 246699 41085 255485 41113
rect 255513 41085 255547 41113
rect 255575 41085 255609 41113
rect 255637 41085 255671 41113
rect 255699 41085 264485 41113
rect 264513 41085 264547 41113
rect 264575 41085 264609 41113
rect 264637 41085 264671 41113
rect 264699 41085 273485 41113
rect 273513 41085 273547 41113
rect 273575 41085 273609 41113
rect 273637 41085 273671 41113
rect 273699 41085 282485 41113
rect 282513 41085 282547 41113
rect 282575 41085 282609 41113
rect 282637 41085 282671 41113
rect 282699 41085 291485 41113
rect 291513 41085 291547 41113
rect 291575 41085 291609 41113
rect 291637 41085 291671 41113
rect 291699 41085 298728 41113
rect 298756 41085 298790 41113
rect 298818 41085 298852 41113
rect 298880 41085 298914 41113
rect 298942 41085 298990 41113
rect -958 41051 298990 41085
rect -958 41023 -910 41051
rect -882 41023 -848 41051
rect -820 41023 -786 41051
rect -758 41023 -724 41051
rect -696 41023 3485 41051
rect 3513 41023 3547 41051
rect 3575 41023 3609 41051
rect 3637 41023 3671 41051
rect 3699 41023 12485 41051
rect 12513 41023 12547 41051
rect 12575 41023 12609 41051
rect 12637 41023 12671 41051
rect 12699 41023 21485 41051
rect 21513 41023 21547 41051
rect 21575 41023 21609 41051
rect 21637 41023 21671 41051
rect 21699 41023 30485 41051
rect 30513 41023 30547 41051
rect 30575 41023 30609 41051
rect 30637 41023 30671 41051
rect 30699 41023 39485 41051
rect 39513 41023 39547 41051
rect 39575 41023 39609 41051
rect 39637 41023 39671 41051
rect 39699 41023 48485 41051
rect 48513 41023 48547 41051
rect 48575 41023 48609 41051
rect 48637 41023 48671 41051
rect 48699 41023 57485 41051
rect 57513 41023 57547 41051
rect 57575 41023 57609 41051
rect 57637 41023 57671 41051
rect 57699 41023 66485 41051
rect 66513 41023 66547 41051
rect 66575 41023 66609 41051
rect 66637 41023 66671 41051
rect 66699 41023 75485 41051
rect 75513 41023 75547 41051
rect 75575 41023 75609 41051
rect 75637 41023 75671 41051
rect 75699 41023 84485 41051
rect 84513 41023 84547 41051
rect 84575 41023 84609 41051
rect 84637 41023 84671 41051
rect 84699 41023 93485 41051
rect 93513 41023 93547 41051
rect 93575 41023 93609 41051
rect 93637 41023 93671 41051
rect 93699 41023 102485 41051
rect 102513 41023 102547 41051
rect 102575 41023 102609 41051
rect 102637 41023 102671 41051
rect 102699 41023 111485 41051
rect 111513 41023 111547 41051
rect 111575 41023 111609 41051
rect 111637 41023 111671 41051
rect 111699 41023 120485 41051
rect 120513 41023 120547 41051
rect 120575 41023 120609 41051
rect 120637 41023 120671 41051
rect 120699 41023 129485 41051
rect 129513 41023 129547 41051
rect 129575 41023 129609 41051
rect 129637 41023 129671 41051
rect 129699 41023 138485 41051
rect 138513 41023 138547 41051
rect 138575 41023 138609 41051
rect 138637 41023 138671 41051
rect 138699 41023 147485 41051
rect 147513 41023 147547 41051
rect 147575 41023 147609 41051
rect 147637 41023 147671 41051
rect 147699 41023 156485 41051
rect 156513 41023 156547 41051
rect 156575 41023 156609 41051
rect 156637 41023 156671 41051
rect 156699 41023 165485 41051
rect 165513 41023 165547 41051
rect 165575 41023 165609 41051
rect 165637 41023 165671 41051
rect 165699 41023 174485 41051
rect 174513 41023 174547 41051
rect 174575 41023 174609 41051
rect 174637 41023 174671 41051
rect 174699 41023 183485 41051
rect 183513 41023 183547 41051
rect 183575 41023 183609 41051
rect 183637 41023 183671 41051
rect 183699 41023 192485 41051
rect 192513 41023 192547 41051
rect 192575 41023 192609 41051
rect 192637 41023 192671 41051
rect 192699 41023 201485 41051
rect 201513 41023 201547 41051
rect 201575 41023 201609 41051
rect 201637 41023 201671 41051
rect 201699 41023 210485 41051
rect 210513 41023 210547 41051
rect 210575 41023 210609 41051
rect 210637 41023 210671 41051
rect 210699 41023 219485 41051
rect 219513 41023 219547 41051
rect 219575 41023 219609 41051
rect 219637 41023 219671 41051
rect 219699 41023 228485 41051
rect 228513 41023 228547 41051
rect 228575 41023 228609 41051
rect 228637 41023 228671 41051
rect 228699 41023 237485 41051
rect 237513 41023 237547 41051
rect 237575 41023 237609 41051
rect 237637 41023 237671 41051
rect 237699 41023 246485 41051
rect 246513 41023 246547 41051
rect 246575 41023 246609 41051
rect 246637 41023 246671 41051
rect 246699 41023 255485 41051
rect 255513 41023 255547 41051
rect 255575 41023 255609 41051
rect 255637 41023 255671 41051
rect 255699 41023 264485 41051
rect 264513 41023 264547 41051
rect 264575 41023 264609 41051
rect 264637 41023 264671 41051
rect 264699 41023 273485 41051
rect 273513 41023 273547 41051
rect 273575 41023 273609 41051
rect 273637 41023 273671 41051
rect 273699 41023 282485 41051
rect 282513 41023 282547 41051
rect 282575 41023 282609 41051
rect 282637 41023 282671 41051
rect 282699 41023 291485 41051
rect 291513 41023 291547 41051
rect 291575 41023 291609 41051
rect 291637 41023 291671 41051
rect 291699 41023 298728 41051
rect 298756 41023 298790 41051
rect 298818 41023 298852 41051
rect 298880 41023 298914 41051
rect 298942 41023 298990 41051
rect -958 40989 298990 41023
rect -958 40961 -910 40989
rect -882 40961 -848 40989
rect -820 40961 -786 40989
rect -758 40961 -724 40989
rect -696 40961 3485 40989
rect 3513 40961 3547 40989
rect 3575 40961 3609 40989
rect 3637 40961 3671 40989
rect 3699 40961 12485 40989
rect 12513 40961 12547 40989
rect 12575 40961 12609 40989
rect 12637 40961 12671 40989
rect 12699 40961 21485 40989
rect 21513 40961 21547 40989
rect 21575 40961 21609 40989
rect 21637 40961 21671 40989
rect 21699 40961 30485 40989
rect 30513 40961 30547 40989
rect 30575 40961 30609 40989
rect 30637 40961 30671 40989
rect 30699 40961 39485 40989
rect 39513 40961 39547 40989
rect 39575 40961 39609 40989
rect 39637 40961 39671 40989
rect 39699 40961 48485 40989
rect 48513 40961 48547 40989
rect 48575 40961 48609 40989
rect 48637 40961 48671 40989
rect 48699 40961 57485 40989
rect 57513 40961 57547 40989
rect 57575 40961 57609 40989
rect 57637 40961 57671 40989
rect 57699 40961 66485 40989
rect 66513 40961 66547 40989
rect 66575 40961 66609 40989
rect 66637 40961 66671 40989
rect 66699 40961 75485 40989
rect 75513 40961 75547 40989
rect 75575 40961 75609 40989
rect 75637 40961 75671 40989
rect 75699 40961 84485 40989
rect 84513 40961 84547 40989
rect 84575 40961 84609 40989
rect 84637 40961 84671 40989
rect 84699 40961 93485 40989
rect 93513 40961 93547 40989
rect 93575 40961 93609 40989
rect 93637 40961 93671 40989
rect 93699 40961 102485 40989
rect 102513 40961 102547 40989
rect 102575 40961 102609 40989
rect 102637 40961 102671 40989
rect 102699 40961 111485 40989
rect 111513 40961 111547 40989
rect 111575 40961 111609 40989
rect 111637 40961 111671 40989
rect 111699 40961 120485 40989
rect 120513 40961 120547 40989
rect 120575 40961 120609 40989
rect 120637 40961 120671 40989
rect 120699 40961 129485 40989
rect 129513 40961 129547 40989
rect 129575 40961 129609 40989
rect 129637 40961 129671 40989
rect 129699 40961 138485 40989
rect 138513 40961 138547 40989
rect 138575 40961 138609 40989
rect 138637 40961 138671 40989
rect 138699 40961 147485 40989
rect 147513 40961 147547 40989
rect 147575 40961 147609 40989
rect 147637 40961 147671 40989
rect 147699 40961 156485 40989
rect 156513 40961 156547 40989
rect 156575 40961 156609 40989
rect 156637 40961 156671 40989
rect 156699 40961 165485 40989
rect 165513 40961 165547 40989
rect 165575 40961 165609 40989
rect 165637 40961 165671 40989
rect 165699 40961 174485 40989
rect 174513 40961 174547 40989
rect 174575 40961 174609 40989
rect 174637 40961 174671 40989
rect 174699 40961 183485 40989
rect 183513 40961 183547 40989
rect 183575 40961 183609 40989
rect 183637 40961 183671 40989
rect 183699 40961 192485 40989
rect 192513 40961 192547 40989
rect 192575 40961 192609 40989
rect 192637 40961 192671 40989
rect 192699 40961 201485 40989
rect 201513 40961 201547 40989
rect 201575 40961 201609 40989
rect 201637 40961 201671 40989
rect 201699 40961 210485 40989
rect 210513 40961 210547 40989
rect 210575 40961 210609 40989
rect 210637 40961 210671 40989
rect 210699 40961 219485 40989
rect 219513 40961 219547 40989
rect 219575 40961 219609 40989
rect 219637 40961 219671 40989
rect 219699 40961 228485 40989
rect 228513 40961 228547 40989
rect 228575 40961 228609 40989
rect 228637 40961 228671 40989
rect 228699 40961 237485 40989
rect 237513 40961 237547 40989
rect 237575 40961 237609 40989
rect 237637 40961 237671 40989
rect 237699 40961 246485 40989
rect 246513 40961 246547 40989
rect 246575 40961 246609 40989
rect 246637 40961 246671 40989
rect 246699 40961 255485 40989
rect 255513 40961 255547 40989
rect 255575 40961 255609 40989
rect 255637 40961 255671 40989
rect 255699 40961 264485 40989
rect 264513 40961 264547 40989
rect 264575 40961 264609 40989
rect 264637 40961 264671 40989
rect 264699 40961 273485 40989
rect 273513 40961 273547 40989
rect 273575 40961 273609 40989
rect 273637 40961 273671 40989
rect 273699 40961 282485 40989
rect 282513 40961 282547 40989
rect 282575 40961 282609 40989
rect 282637 40961 282671 40989
rect 282699 40961 291485 40989
rect 291513 40961 291547 40989
rect 291575 40961 291609 40989
rect 291637 40961 291671 40989
rect 291699 40961 298728 40989
rect 298756 40961 298790 40989
rect 298818 40961 298852 40989
rect 298880 40961 298914 40989
rect 298942 40961 298990 40989
rect -958 40913 298990 40961
rect -958 38175 298990 38223
rect -958 38147 -430 38175
rect -402 38147 -368 38175
rect -340 38147 -306 38175
rect -278 38147 -244 38175
rect -216 38147 1625 38175
rect 1653 38147 1687 38175
rect 1715 38147 1749 38175
rect 1777 38147 1811 38175
rect 1839 38147 10625 38175
rect 10653 38147 10687 38175
rect 10715 38147 10749 38175
rect 10777 38147 10811 38175
rect 10839 38147 19625 38175
rect 19653 38147 19687 38175
rect 19715 38147 19749 38175
rect 19777 38147 19811 38175
rect 19839 38147 28625 38175
rect 28653 38147 28687 38175
rect 28715 38147 28749 38175
rect 28777 38147 28811 38175
rect 28839 38147 37625 38175
rect 37653 38147 37687 38175
rect 37715 38147 37749 38175
rect 37777 38147 37811 38175
rect 37839 38147 46625 38175
rect 46653 38147 46687 38175
rect 46715 38147 46749 38175
rect 46777 38147 46811 38175
rect 46839 38147 55625 38175
rect 55653 38147 55687 38175
rect 55715 38147 55749 38175
rect 55777 38147 55811 38175
rect 55839 38147 64625 38175
rect 64653 38147 64687 38175
rect 64715 38147 64749 38175
rect 64777 38147 64811 38175
rect 64839 38147 73625 38175
rect 73653 38147 73687 38175
rect 73715 38147 73749 38175
rect 73777 38147 73811 38175
rect 73839 38147 82625 38175
rect 82653 38147 82687 38175
rect 82715 38147 82749 38175
rect 82777 38147 82811 38175
rect 82839 38147 91625 38175
rect 91653 38147 91687 38175
rect 91715 38147 91749 38175
rect 91777 38147 91811 38175
rect 91839 38147 100625 38175
rect 100653 38147 100687 38175
rect 100715 38147 100749 38175
rect 100777 38147 100811 38175
rect 100839 38147 109625 38175
rect 109653 38147 109687 38175
rect 109715 38147 109749 38175
rect 109777 38147 109811 38175
rect 109839 38147 118625 38175
rect 118653 38147 118687 38175
rect 118715 38147 118749 38175
rect 118777 38147 118811 38175
rect 118839 38147 127625 38175
rect 127653 38147 127687 38175
rect 127715 38147 127749 38175
rect 127777 38147 127811 38175
rect 127839 38147 136625 38175
rect 136653 38147 136687 38175
rect 136715 38147 136749 38175
rect 136777 38147 136811 38175
rect 136839 38147 145625 38175
rect 145653 38147 145687 38175
rect 145715 38147 145749 38175
rect 145777 38147 145811 38175
rect 145839 38147 154625 38175
rect 154653 38147 154687 38175
rect 154715 38147 154749 38175
rect 154777 38147 154811 38175
rect 154839 38147 163625 38175
rect 163653 38147 163687 38175
rect 163715 38147 163749 38175
rect 163777 38147 163811 38175
rect 163839 38147 172625 38175
rect 172653 38147 172687 38175
rect 172715 38147 172749 38175
rect 172777 38147 172811 38175
rect 172839 38147 181625 38175
rect 181653 38147 181687 38175
rect 181715 38147 181749 38175
rect 181777 38147 181811 38175
rect 181839 38147 190625 38175
rect 190653 38147 190687 38175
rect 190715 38147 190749 38175
rect 190777 38147 190811 38175
rect 190839 38147 199625 38175
rect 199653 38147 199687 38175
rect 199715 38147 199749 38175
rect 199777 38147 199811 38175
rect 199839 38147 208625 38175
rect 208653 38147 208687 38175
rect 208715 38147 208749 38175
rect 208777 38147 208811 38175
rect 208839 38147 217625 38175
rect 217653 38147 217687 38175
rect 217715 38147 217749 38175
rect 217777 38147 217811 38175
rect 217839 38147 226625 38175
rect 226653 38147 226687 38175
rect 226715 38147 226749 38175
rect 226777 38147 226811 38175
rect 226839 38147 235625 38175
rect 235653 38147 235687 38175
rect 235715 38147 235749 38175
rect 235777 38147 235811 38175
rect 235839 38147 244625 38175
rect 244653 38147 244687 38175
rect 244715 38147 244749 38175
rect 244777 38147 244811 38175
rect 244839 38147 253625 38175
rect 253653 38147 253687 38175
rect 253715 38147 253749 38175
rect 253777 38147 253811 38175
rect 253839 38147 262625 38175
rect 262653 38147 262687 38175
rect 262715 38147 262749 38175
rect 262777 38147 262811 38175
rect 262839 38147 271625 38175
rect 271653 38147 271687 38175
rect 271715 38147 271749 38175
rect 271777 38147 271811 38175
rect 271839 38147 280625 38175
rect 280653 38147 280687 38175
rect 280715 38147 280749 38175
rect 280777 38147 280811 38175
rect 280839 38147 289625 38175
rect 289653 38147 289687 38175
rect 289715 38147 289749 38175
rect 289777 38147 289811 38175
rect 289839 38147 298248 38175
rect 298276 38147 298310 38175
rect 298338 38147 298372 38175
rect 298400 38147 298434 38175
rect 298462 38147 298990 38175
rect -958 38113 298990 38147
rect -958 38085 -430 38113
rect -402 38085 -368 38113
rect -340 38085 -306 38113
rect -278 38085 -244 38113
rect -216 38085 1625 38113
rect 1653 38085 1687 38113
rect 1715 38085 1749 38113
rect 1777 38085 1811 38113
rect 1839 38085 10625 38113
rect 10653 38085 10687 38113
rect 10715 38085 10749 38113
rect 10777 38085 10811 38113
rect 10839 38085 19625 38113
rect 19653 38085 19687 38113
rect 19715 38085 19749 38113
rect 19777 38085 19811 38113
rect 19839 38085 28625 38113
rect 28653 38085 28687 38113
rect 28715 38085 28749 38113
rect 28777 38085 28811 38113
rect 28839 38085 37625 38113
rect 37653 38085 37687 38113
rect 37715 38085 37749 38113
rect 37777 38085 37811 38113
rect 37839 38085 46625 38113
rect 46653 38085 46687 38113
rect 46715 38085 46749 38113
rect 46777 38085 46811 38113
rect 46839 38085 55625 38113
rect 55653 38085 55687 38113
rect 55715 38085 55749 38113
rect 55777 38085 55811 38113
rect 55839 38085 64625 38113
rect 64653 38085 64687 38113
rect 64715 38085 64749 38113
rect 64777 38085 64811 38113
rect 64839 38085 73625 38113
rect 73653 38085 73687 38113
rect 73715 38085 73749 38113
rect 73777 38085 73811 38113
rect 73839 38085 82625 38113
rect 82653 38085 82687 38113
rect 82715 38085 82749 38113
rect 82777 38085 82811 38113
rect 82839 38085 91625 38113
rect 91653 38085 91687 38113
rect 91715 38085 91749 38113
rect 91777 38085 91811 38113
rect 91839 38085 100625 38113
rect 100653 38085 100687 38113
rect 100715 38085 100749 38113
rect 100777 38085 100811 38113
rect 100839 38085 109625 38113
rect 109653 38085 109687 38113
rect 109715 38085 109749 38113
rect 109777 38085 109811 38113
rect 109839 38085 118625 38113
rect 118653 38085 118687 38113
rect 118715 38085 118749 38113
rect 118777 38085 118811 38113
rect 118839 38085 127625 38113
rect 127653 38085 127687 38113
rect 127715 38085 127749 38113
rect 127777 38085 127811 38113
rect 127839 38085 136625 38113
rect 136653 38085 136687 38113
rect 136715 38085 136749 38113
rect 136777 38085 136811 38113
rect 136839 38085 145625 38113
rect 145653 38085 145687 38113
rect 145715 38085 145749 38113
rect 145777 38085 145811 38113
rect 145839 38085 154625 38113
rect 154653 38085 154687 38113
rect 154715 38085 154749 38113
rect 154777 38085 154811 38113
rect 154839 38085 163625 38113
rect 163653 38085 163687 38113
rect 163715 38085 163749 38113
rect 163777 38085 163811 38113
rect 163839 38085 172625 38113
rect 172653 38085 172687 38113
rect 172715 38085 172749 38113
rect 172777 38085 172811 38113
rect 172839 38085 181625 38113
rect 181653 38085 181687 38113
rect 181715 38085 181749 38113
rect 181777 38085 181811 38113
rect 181839 38085 190625 38113
rect 190653 38085 190687 38113
rect 190715 38085 190749 38113
rect 190777 38085 190811 38113
rect 190839 38085 199625 38113
rect 199653 38085 199687 38113
rect 199715 38085 199749 38113
rect 199777 38085 199811 38113
rect 199839 38085 208625 38113
rect 208653 38085 208687 38113
rect 208715 38085 208749 38113
rect 208777 38085 208811 38113
rect 208839 38085 217625 38113
rect 217653 38085 217687 38113
rect 217715 38085 217749 38113
rect 217777 38085 217811 38113
rect 217839 38085 226625 38113
rect 226653 38085 226687 38113
rect 226715 38085 226749 38113
rect 226777 38085 226811 38113
rect 226839 38085 235625 38113
rect 235653 38085 235687 38113
rect 235715 38085 235749 38113
rect 235777 38085 235811 38113
rect 235839 38085 244625 38113
rect 244653 38085 244687 38113
rect 244715 38085 244749 38113
rect 244777 38085 244811 38113
rect 244839 38085 253625 38113
rect 253653 38085 253687 38113
rect 253715 38085 253749 38113
rect 253777 38085 253811 38113
rect 253839 38085 262625 38113
rect 262653 38085 262687 38113
rect 262715 38085 262749 38113
rect 262777 38085 262811 38113
rect 262839 38085 271625 38113
rect 271653 38085 271687 38113
rect 271715 38085 271749 38113
rect 271777 38085 271811 38113
rect 271839 38085 280625 38113
rect 280653 38085 280687 38113
rect 280715 38085 280749 38113
rect 280777 38085 280811 38113
rect 280839 38085 289625 38113
rect 289653 38085 289687 38113
rect 289715 38085 289749 38113
rect 289777 38085 289811 38113
rect 289839 38085 298248 38113
rect 298276 38085 298310 38113
rect 298338 38085 298372 38113
rect 298400 38085 298434 38113
rect 298462 38085 298990 38113
rect -958 38051 298990 38085
rect -958 38023 -430 38051
rect -402 38023 -368 38051
rect -340 38023 -306 38051
rect -278 38023 -244 38051
rect -216 38023 1625 38051
rect 1653 38023 1687 38051
rect 1715 38023 1749 38051
rect 1777 38023 1811 38051
rect 1839 38023 10625 38051
rect 10653 38023 10687 38051
rect 10715 38023 10749 38051
rect 10777 38023 10811 38051
rect 10839 38023 19625 38051
rect 19653 38023 19687 38051
rect 19715 38023 19749 38051
rect 19777 38023 19811 38051
rect 19839 38023 28625 38051
rect 28653 38023 28687 38051
rect 28715 38023 28749 38051
rect 28777 38023 28811 38051
rect 28839 38023 37625 38051
rect 37653 38023 37687 38051
rect 37715 38023 37749 38051
rect 37777 38023 37811 38051
rect 37839 38023 46625 38051
rect 46653 38023 46687 38051
rect 46715 38023 46749 38051
rect 46777 38023 46811 38051
rect 46839 38023 55625 38051
rect 55653 38023 55687 38051
rect 55715 38023 55749 38051
rect 55777 38023 55811 38051
rect 55839 38023 64625 38051
rect 64653 38023 64687 38051
rect 64715 38023 64749 38051
rect 64777 38023 64811 38051
rect 64839 38023 73625 38051
rect 73653 38023 73687 38051
rect 73715 38023 73749 38051
rect 73777 38023 73811 38051
rect 73839 38023 82625 38051
rect 82653 38023 82687 38051
rect 82715 38023 82749 38051
rect 82777 38023 82811 38051
rect 82839 38023 91625 38051
rect 91653 38023 91687 38051
rect 91715 38023 91749 38051
rect 91777 38023 91811 38051
rect 91839 38023 100625 38051
rect 100653 38023 100687 38051
rect 100715 38023 100749 38051
rect 100777 38023 100811 38051
rect 100839 38023 109625 38051
rect 109653 38023 109687 38051
rect 109715 38023 109749 38051
rect 109777 38023 109811 38051
rect 109839 38023 118625 38051
rect 118653 38023 118687 38051
rect 118715 38023 118749 38051
rect 118777 38023 118811 38051
rect 118839 38023 127625 38051
rect 127653 38023 127687 38051
rect 127715 38023 127749 38051
rect 127777 38023 127811 38051
rect 127839 38023 136625 38051
rect 136653 38023 136687 38051
rect 136715 38023 136749 38051
rect 136777 38023 136811 38051
rect 136839 38023 145625 38051
rect 145653 38023 145687 38051
rect 145715 38023 145749 38051
rect 145777 38023 145811 38051
rect 145839 38023 154625 38051
rect 154653 38023 154687 38051
rect 154715 38023 154749 38051
rect 154777 38023 154811 38051
rect 154839 38023 163625 38051
rect 163653 38023 163687 38051
rect 163715 38023 163749 38051
rect 163777 38023 163811 38051
rect 163839 38023 172625 38051
rect 172653 38023 172687 38051
rect 172715 38023 172749 38051
rect 172777 38023 172811 38051
rect 172839 38023 181625 38051
rect 181653 38023 181687 38051
rect 181715 38023 181749 38051
rect 181777 38023 181811 38051
rect 181839 38023 190625 38051
rect 190653 38023 190687 38051
rect 190715 38023 190749 38051
rect 190777 38023 190811 38051
rect 190839 38023 199625 38051
rect 199653 38023 199687 38051
rect 199715 38023 199749 38051
rect 199777 38023 199811 38051
rect 199839 38023 208625 38051
rect 208653 38023 208687 38051
rect 208715 38023 208749 38051
rect 208777 38023 208811 38051
rect 208839 38023 217625 38051
rect 217653 38023 217687 38051
rect 217715 38023 217749 38051
rect 217777 38023 217811 38051
rect 217839 38023 226625 38051
rect 226653 38023 226687 38051
rect 226715 38023 226749 38051
rect 226777 38023 226811 38051
rect 226839 38023 235625 38051
rect 235653 38023 235687 38051
rect 235715 38023 235749 38051
rect 235777 38023 235811 38051
rect 235839 38023 244625 38051
rect 244653 38023 244687 38051
rect 244715 38023 244749 38051
rect 244777 38023 244811 38051
rect 244839 38023 253625 38051
rect 253653 38023 253687 38051
rect 253715 38023 253749 38051
rect 253777 38023 253811 38051
rect 253839 38023 262625 38051
rect 262653 38023 262687 38051
rect 262715 38023 262749 38051
rect 262777 38023 262811 38051
rect 262839 38023 271625 38051
rect 271653 38023 271687 38051
rect 271715 38023 271749 38051
rect 271777 38023 271811 38051
rect 271839 38023 280625 38051
rect 280653 38023 280687 38051
rect 280715 38023 280749 38051
rect 280777 38023 280811 38051
rect 280839 38023 289625 38051
rect 289653 38023 289687 38051
rect 289715 38023 289749 38051
rect 289777 38023 289811 38051
rect 289839 38023 298248 38051
rect 298276 38023 298310 38051
rect 298338 38023 298372 38051
rect 298400 38023 298434 38051
rect 298462 38023 298990 38051
rect -958 37989 298990 38023
rect -958 37961 -430 37989
rect -402 37961 -368 37989
rect -340 37961 -306 37989
rect -278 37961 -244 37989
rect -216 37961 1625 37989
rect 1653 37961 1687 37989
rect 1715 37961 1749 37989
rect 1777 37961 1811 37989
rect 1839 37961 10625 37989
rect 10653 37961 10687 37989
rect 10715 37961 10749 37989
rect 10777 37961 10811 37989
rect 10839 37961 19625 37989
rect 19653 37961 19687 37989
rect 19715 37961 19749 37989
rect 19777 37961 19811 37989
rect 19839 37961 28625 37989
rect 28653 37961 28687 37989
rect 28715 37961 28749 37989
rect 28777 37961 28811 37989
rect 28839 37961 37625 37989
rect 37653 37961 37687 37989
rect 37715 37961 37749 37989
rect 37777 37961 37811 37989
rect 37839 37961 46625 37989
rect 46653 37961 46687 37989
rect 46715 37961 46749 37989
rect 46777 37961 46811 37989
rect 46839 37961 55625 37989
rect 55653 37961 55687 37989
rect 55715 37961 55749 37989
rect 55777 37961 55811 37989
rect 55839 37961 64625 37989
rect 64653 37961 64687 37989
rect 64715 37961 64749 37989
rect 64777 37961 64811 37989
rect 64839 37961 73625 37989
rect 73653 37961 73687 37989
rect 73715 37961 73749 37989
rect 73777 37961 73811 37989
rect 73839 37961 82625 37989
rect 82653 37961 82687 37989
rect 82715 37961 82749 37989
rect 82777 37961 82811 37989
rect 82839 37961 91625 37989
rect 91653 37961 91687 37989
rect 91715 37961 91749 37989
rect 91777 37961 91811 37989
rect 91839 37961 100625 37989
rect 100653 37961 100687 37989
rect 100715 37961 100749 37989
rect 100777 37961 100811 37989
rect 100839 37961 109625 37989
rect 109653 37961 109687 37989
rect 109715 37961 109749 37989
rect 109777 37961 109811 37989
rect 109839 37961 118625 37989
rect 118653 37961 118687 37989
rect 118715 37961 118749 37989
rect 118777 37961 118811 37989
rect 118839 37961 127625 37989
rect 127653 37961 127687 37989
rect 127715 37961 127749 37989
rect 127777 37961 127811 37989
rect 127839 37961 136625 37989
rect 136653 37961 136687 37989
rect 136715 37961 136749 37989
rect 136777 37961 136811 37989
rect 136839 37961 145625 37989
rect 145653 37961 145687 37989
rect 145715 37961 145749 37989
rect 145777 37961 145811 37989
rect 145839 37961 154625 37989
rect 154653 37961 154687 37989
rect 154715 37961 154749 37989
rect 154777 37961 154811 37989
rect 154839 37961 163625 37989
rect 163653 37961 163687 37989
rect 163715 37961 163749 37989
rect 163777 37961 163811 37989
rect 163839 37961 172625 37989
rect 172653 37961 172687 37989
rect 172715 37961 172749 37989
rect 172777 37961 172811 37989
rect 172839 37961 181625 37989
rect 181653 37961 181687 37989
rect 181715 37961 181749 37989
rect 181777 37961 181811 37989
rect 181839 37961 190625 37989
rect 190653 37961 190687 37989
rect 190715 37961 190749 37989
rect 190777 37961 190811 37989
rect 190839 37961 199625 37989
rect 199653 37961 199687 37989
rect 199715 37961 199749 37989
rect 199777 37961 199811 37989
rect 199839 37961 208625 37989
rect 208653 37961 208687 37989
rect 208715 37961 208749 37989
rect 208777 37961 208811 37989
rect 208839 37961 217625 37989
rect 217653 37961 217687 37989
rect 217715 37961 217749 37989
rect 217777 37961 217811 37989
rect 217839 37961 226625 37989
rect 226653 37961 226687 37989
rect 226715 37961 226749 37989
rect 226777 37961 226811 37989
rect 226839 37961 235625 37989
rect 235653 37961 235687 37989
rect 235715 37961 235749 37989
rect 235777 37961 235811 37989
rect 235839 37961 244625 37989
rect 244653 37961 244687 37989
rect 244715 37961 244749 37989
rect 244777 37961 244811 37989
rect 244839 37961 253625 37989
rect 253653 37961 253687 37989
rect 253715 37961 253749 37989
rect 253777 37961 253811 37989
rect 253839 37961 262625 37989
rect 262653 37961 262687 37989
rect 262715 37961 262749 37989
rect 262777 37961 262811 37989
rect 262839 37961 271625 37989
rect 271653 37961 271687 37989
rect 271715 37961 271749 37989
rect 271777 37961 271811 37989
rect 271839 37961 280625 37989
rect 280653 37961 280687 37989
rect 280715 37961 280749 37989
rect 280777 37961 280811 37989
rect 280839 37961 289625 37989
rect 289653 37961 289687 37989
rect 289715 37961 289749 37989
rect 289777 37961 289811 37989
rect 289839 37961 298248 37989
rect 298276 37961 298310 37989
rect 298338 37961 298372 37989
rect 298400 37961 298434 37989
rect 298462 37961 298990 37989
rect -958 37913 298990 37961
rect -958 32175 298990 32223
rect -958 32147 -910 32175
rect -882 32147 -848 32175
rect -820 32147 -786 32175
rect -758 32147 -724 32175
rect -696 32147 3485 32175
rect 3513 32147 3547 32175
rect 3575 32147 3609 32175
rect 3637 32147 3671 32175
rect 3699 32147 12485 32175
rect 12513 32147 12547 32175
rect 12575 32147 12609 32175
rect 12637 32147 12671 32175
rect 12699 32147 21485 32175
rect 21513 32147 21547 32175
rect 21575 32147 21609 32175
rect 21637 32147 21671 32175
rect 21699 32147 30485 32175
rect 30513 32147 30547 32175
rect 30575 32147 30609 32175
rect 30637 32147 30671 32175
rect 30699 32147 39485 32175
rect 39513 32147 39547 32175
rect 39575 32147 39609 32175
rect 39637 32147 39671 32175
rect 39699 32147 48485 32175
rect 48513 32147 48547 32175
rect 48575 32147 48609 32175
rect 48637 32147 48671 32175
rect 48699 32147 57485 32175
rect 57513 32147 57547 32175
rect 57575 32147 57609 32175
rect 57637 32147 57671 32175
rect 57699 32147 66485 32175
rect 66513 32147 66547 32175
rect 66575 32147 66609 32175
rect 66637 32147 66671 32175
rect 66699 32147 75485 32175
rect 75513 32147 75547 32175
rect 75575 32147 75609 32175
rect 75637 32147 75671 32175
rect 75699 32147 84485 32175
rect 84513 32147 84547 32175
rect 84575 32147 84609 32175
rect 84637 32147 84671 32175
rect 84699 32147 93485 32175
rect 93513 32147 93547 32175
rect 93575 32147 93609 32175
rect 93637 32147 93671 32175
rect 93699 32147 102485 32175
rect 102513 32147 102547 32175
rect 102575 32147 102609 32175
rect 102637 32147 102671 32175
rect 102699 32147 111485 32175
rect 111513 32147 111547 32175
rect 111575 32147 111609 32175
rect 111637 32147 111671 32175
rect 111699 32147 120485 32175
rect 120513 32147 120547 32175
rect 120575 32147 120609 32175
rect 120637 32147 120671 32175
rect 120699 32147 129485 32175
rect 129513 32147 129547 32175
rect 129575 32147 129609 32175
rect 129637 32147 129671 32175
rect 129699 32147 138485 32175
rect 138513 32147 138547 32175
rect 138575 32147 138609 32175
rect 138637 32147 138671 32175
rect 138699 32147 147485 32175
rect 147513 32147 147547 32175
rect 147575 32147 147609 32175
rect 147637 32147 147671 32175
rect 147699 32147 156485 32175
rect 156513 32147 156547 32175
rect 156575 32147 156609 32175
rect 156637 32147 156671 32175
rect 156699 32147 165485 32175
rect 165513 32147 165547 32175
rect 165575 32147 165609 32175
rect 165637 32147 165671 32175
rect 165699 32147 174485 32175
rect 174513 32147 174547 32175
rect 174575 32147 174609 32175
rect 174637 32147 174671 32175
rect 174699 32147 183485 32175
rect 183513 32147 183547 32175
rect 183575 32147 183609 32175
rect 183637 32147 183671 32175
rect 183699 32147 192485 32175
rect 192513 32147 192547 32175
rect 192575 32147 192609 32175
rect 192637 32147 192671 32175
rect 192699 32147 201485 32175
rect 201513 32147 201547 32175
rect 201575 32147 201609 32175
rect 201637 32147 201671 32175
rect 201699 32147 210485 32175
rect 210513 32147 210547 32175
rect 210575 32147 210609 32175
rect 210637 32147 210671 32175
rect 210699 32147 219485 32175
rect 219513 32147 219547 32175
rect 219575 32147 219609 32175
rect 219637 32147 219671 32175
rect 219699 32147 228485 32175
rect 228513 32147 228547 32175
rect 228575 32147 228609 32175
rect 228637 32147 228671 32175
rect 228699 32147 237485 32175
rect 237513 32147 237547 32175
rect 237575 32147 237609 32175
rect 237637 32147 237671 32175
rect 237699 32147 246485 32175
rect 246513 32147 246547 32175
rect 246575 32147 246609 32175
rect 246637 32147 246671 32175
rect 246699 32147 255485 32175
rect 255513 32147 255547 32175
rect 255575 32147 255609 32175
rect 255637 32147 255671 32175
rect 255699 32147 264485 32175
rect 264513 32147 264547 32175
rect 264575 32147 264609 32175
rect 264637 32147 264671 32175
rect 264699 32147 273485 32175
rect 273513 32147 273547 32175
rect 273575 32147 273609 32175
rect 273637 32147 273671 32175
rect 273699 32147 282485 32175
rect 282513 32147 282547 32175
rect 282575 32147 282609 32175
rect 282637 32147 282671 32175
rect 282699 32147 291485 32175
rect 291513 32147 291547 32175
rect 291575 32147 291609 32175
rect 291637 32147 291671 32175
rect 291699 32147 298728 32175
rect 298756 32147 298790 32175
rect 298818 32147 298852 32175
rect 298880 32147 298914 32175
rect 298942 32147 298990 32175
rect -958 32113 298990 32147
rect -958 32085 -910 32113
rect -882 32085 -848 32113
rect -820 32085 -786 32113
rect -758 32085 -724 32113
rect -696 32085 3485 32113
rect 3513 32085 3547 32113
rect 3575 32085 3609 32113
rect 3637 32085 3671 32113
rect 3699 32085 12485 32113
rect 12513 32085 12547 32113
rect 12575 32085 12609 32113
rect 12637 32085 12671 32113
rect 12699 32085 21485 32113
rect 21513 32085 21547 32113
rect 21575 32085 21609 32113
rect 21637 32085 21671 32113
rect 21699 32085 30485 32113
rect 30513 32085 30547 32113
rect 30575 32085 30609 32113
rect 30637 32085 30671 32113
rect 30699 32085 39485 32113
rect 39513 32085 39547 32113
rect 39575 32085 39609 32113
rect 39637 32085 39671 32113
rect 39699 32085 48485 32113
rect 48513 32085 48547 32113
rect 48575 32085 48609 32113
rect 48637 32085 48671 32113
rect 48699 32085 57485 32113
rect 57513 32085 57547 32113
rect 57575 32085 57609 32113
rect 57637 32085 57671 32113
rect 57699 32085 66485 32113
rect 66513 32085 66547 32113
rect 66575 32085 66609 32113
rect 66637 32085 66671 32113
rect 66699 32085 75485 32113
rect 75513 32085 75547 32113
rect 75575 32085 75609 32113
rect 75637 32085 75671 32113
rect 75699 32085 84485 32113
rect 84513 32085 84547 32113
rect 84575 32085 84609 32113
rect 84637 32085 84671 32113
rect 84699 32085 93485 32113
rect 93513 32085 93547 32113
rect 93575 32085 93609 32113
rect 93637 32085 93671 32113
rect 93699 32085 102485 32113
rect 102513 32085 102547 32113
rect 102575 32085 102609 32113
rect 102637 32085 102671 32113
rect 102699 32085 111485 32113
rect 111513 32085 111547 32113
rect 111575 32085 111609 32113
rect 111637 32085 111671 32113
rect 111699 32085 120485 32113
rect 120513 32085 120547 32113
rect 120575 32085 120609 32113
rect 120637 32085 120671 32113
rect 120699 32085 129485 32113
rect 129513 32085 129547 32113
rect 129575 32085 129609 32113
rect 129637 32085 129671 32113
rect 129699 32085 138485 32113
rect 138513 32085 138547 32113
rect 138575 32085 138609 32113
rect 138637 32085 138671 32113
rect 138699 32085 147485 32113
rect 147513 32085 147547 32113
rect 147575 32085 147609 32113
rect 147637 32085 147671 32113
rect 147699 32085 156485 32113
rect 156513 32085 156547 32113
rect 156575 32085 156609 32113
rect 156637 32085 156671 32113
rect 156699 32085 165485 32113
rect 165513 32085 165547 32113
rect 165575 32085 165609 32113
rect 165637 32085 165671 32113
rect 165699 32085 174485 32113
rect 174513 32085 174547 32113
rect 174575 32085 174609 32113
rect 174637 32085 174671 32113
rect 174699 32085 183485 32113
rect 183513 32085 183547 32113
rect 183575 32085 183609 32113
rect 183637 32085 183671 32113
rect 183699 32085 192485 32113
rect 192513 32085 192547 32113
rect 192575 32085 192609 32113
rect 192637 32085 192671 32113
rect 192699 32085 201485 32113
rect 201513 32085 201547 32113
rect 201575 32085 201609 32113
rect 201637 32085 201671 32113
rect 201699 32085 210485 32113
rect 210513 32085 210547 32113
rect 210575 32085 210609 32113
rect 210637 32085 210671 32113
rect 210699 32085 219485 32113
rect 219513 32085 219547 32113
rect 219575 32085 219609 32113
rect 219637 32085 219671 32113
rect 219699 32085 228485 32113
rect 228513 32085 228547 32113
rect 228575 32085 228609 32113
rect 228637 32085 228671 32113
rect 228699 32085 237485 32113
rect 237513 32085 237547 32113
rect 237575 32085 237609 32113
rect 237637 32085 237671 32113
rect 237699 32085 246485 32113
rect 246513 32085 246547 32113
rect 246575 32085 246609 32113
rect 246637 32085 246671 32113
rect 246699 32085 255485 32113
rect 255513 32085 255547 32113
rect 255575 32085 255609 32113
rect 255637 32085 255671 32113
rect 255699 32085 264485 32113
rect 264513 32085 264547 32113
rect 264575 32085 264609 32113
rect 264637 32085 264671 32113
rect 264699 32085 273485 32113
rect 273513 32085 273547 32113
rect 273575 32085 273609 32113
rect 273637 32085 273671 32113
rect 273699 32085 282485 32113
rect 282513 32085 282547 32113
rect 282575 32085 282609 32113
rect 282637 32085 282671 32113
rect 282699 32085 291485 32113
rect 291513 32085 291547 32113
rect 291575 32085 291609 32113
rect 291637 32085 291671 32113
rect 291699 32085 298728 32113
rect 298756 32085 298790 32113
rect 298818 32085 298852 32113
rect 298880 32085 298914 32113
rect 298942 32085 298990 32113
rect -958 32051 298990 32085
rect -958 32023 -910 32051
rect -882 32023 -848 32051
rect -820 32023 -786 32051
rect -758 32023 -724 32051
rect -696 32023 3485 32051
rect 3513 32023 3547 32051
rect 3575 32023 3609 32051
rect 3637 32023 3671 32051
rect 3699 32023 12485 32051
rect 12513 32023 12547 32051
rect 12575 32023 12609 32051
rect 12637 32023 12671 32051
rect 12699 32023 21485 32051
rect 21513 32023 21547 32051
rect 21575 32023 21609 32051
rect 21637 32023 21671 32051
rect 21699 32023 30485 32051
rect 30513 32023 30547 32051
rect 30575 32023 30609 32051
rect 30637 32023 30671 32051
rect 30699 32023 39485 32051
rect 39513 32023 39547 32051
rect 39575 32023 39609 32051
rect 39637 32023 39671 32051
rect 39699 32023 48485 32051
rect 48513 32023 48547 32051
rect 48575 32023 48609 32051
rect 48637 32023 48671 32051
rect 48699 32023 57485 32051
rect 57513 32023 57547 32051
rect 57575 32023 57609 32051
rect 57637 32023 57671 32051
rect 57699 32023 66485 32051
rect 66513 32023 66547 32051
rect 66575 32023 66609 32051
rect 66637 32023 66671 32051
rect 66699 32023 75485 32051
rect 75513 32023 75547 32051
rect 75575 32023 75609 32051
rect 75637 32023 75671 32051
rect 75699 32023 84485 32051
rect 84513 32023 84547 32051
rect 84575 32023 84609 32051
rect 84637 32023 84671 32051
rect 84699 32023 93485 32051
rect 93513 32023 93547 32051
rect 93575 32023 93609 32051
rect 93637 32023 93671 32051
rect 93699 32023 102485 32051
rect 102513 32023 102547 32051
rect 102575 32023 102609 32051
rect 102637 32023 102671 32051
rect 102699 32023 111485 32051
rect 111513 32023 111547 32051
rect 111575 32023 111609 32051
rect 111637 32023 111671 32051
rect 111699 32023 120485 32051
rect 120513 32023 120547 32051
rect 120575 32023 120609 32051
rect 120637 32023 120671 32051
rect 120699 32023 129485 32051
rect 129513 32023 129547 32051
rect 129575 32023 129609 32051
rect 129637 32023 129671 32051
rect 129699 32023 138485 32051
rect 138513 32023 138547 32051
rect 138575 32023 138609 32051
rect 138637 32023 138671 32051
rect 138699 32023 147485 32051
rect 147513 32023 147547 32051
rect 147575 32023 147609 32051
rect 147637 32023 147671 32051
rect 147699 32023 156485 32051
rect 156513 32023 156547 32051
rect 156575 32023 156609 32051
rect 156637 32023 156671 32051
rect 156699 32023 165485 32051
rect 165513 32023 165547 32051
rect 165575 32023 165609 32051
rect 165637 32023 165671 32051
rect 165699 32023 174485 32051
rect 174513 32023 174547 32051
rect 174575 32023 174609 32051
rect 174637 32023 174671 32051
rect 174699 32023 183485 32051
rect 183513 32023 183547 32051
rect 183575 32023 183609 32051
rect 183637 32023 183671 32051
rect 183699 32023 192485 32051
rect 192513 32023 192547 32051
rect 192575 32023 192609 32051
rect 192637 32023 192671 32051
rect 192699 32023 201485 32051
rect 201513 32023 201547 32051
rect 201575 32023 201609 32051
rect 201637 32023 201671 32051
rect 201699 32023 210485 32051
rect 210513 32023 210547 32051
rect 210575 32023 210609 32051
rect 210637 32023 210671 32051
rect 210699 32023 219485 32051
rect 219513 32023 219547 32051
rect 219575 32023 219609 32051
rect 219637 32023 219671 32051
rect 219699 32023 228485 32051
rect 228513 32023 228547 32051
rect 228575 32023 228609 32051
rect 228637 32023 228671 32051
rect 228699 32023 237485 32051
rect 237513 32023 237547 32051
rect 237575 32023 237609 32051
rect 237637 32023 237671 32051
rect 237699 32023 246485 32051
rect 246513 32023 246547 32051
rect 246575 32023 246609 32051
rect 246637 32023 246671 32051
rect 246699 32023 255485 32051
rect 255513 32023 255547 32051
rect 255575 32023 255609 32051
rect 255637 32023 255671 32051
rect 255699 32023 264485 32051
rect 264513 32023 264547 32051
rect 264575 32023 264609 32051
rect 264637 32023 264671 32051
rect 264699 32023 273485 32051
rect 273513 32023 273547 32051
rect 273575 32023 273609 32051
rect 273637 32023 273671 32051
rect 273699 32023 282485 32051
rect 282513 32023 282547 32051
rect 282575 32023 282609 32051
rect 282637 32023 282671 32051
rect 282699 32023 291485 32051
rect 291513 32023 291547 32051
rect 291575 32023 291609 32051
rect 291637 32023 291671 32051
rect 291699 32023 298728 32051
rect 298756 32023 298790 32051
rect 298818 32023 298852 32051
rect 298880 32023 298914 32051
rect 298942 32023 298990 32051
rect -958 31989 298990 32023
rect -958 31961 -910 31989
rect -882 31961 -848 31989
rect -820 31961 -786 31989
rect -758 31961 -724 31989
rect -696 31961 3485 31989
rect 3513 31961 3547 31989
rect 3575 31961 3609 31989
rect 3637 31961 3671 31989
rect 3699 31961 12485 31989
rect 12513 31961 12547 31989
rect 12575 31961 12609 31989
rect 12637 31961 12671 31989
rect 12699 31961 21485 31989
rect 21513 31961 21547 31989
rect 21575 31961 21609 31989
rect 21637 31961 21671 31989
rect 21699 31961 30485 31989
rect 30513 31961 30547 31989
rect 30575 31961 30609 31989
rect 30637 31961 30671 31989
rect 30699 31961 39485 31989
rect 39513 31961 39547 31989
rect 39575 31961 39609 31989
rect 39637 31961 39671 31989
rect 39699 31961 48485 31989
rect 48513 31961 48547 31989
rect 48575 31961 48609 31989
rect 48637 31961 48671 31989
rect 48699 31961 57485 31989
rect 57513 31961 57547 31989
rect 57575 31961 57609 31989
rect 57637 31961 57671 31989
rect 57699 31961 66485 31989
rect 66513 31961 66547 31989
rect 66575 31961 66609 31989
rect 66637 31961 66671 31989
rect 66699 31961 75485 31989
rect 75513 31961 75547 31989
rect 75575 31961 75609 31989
rect 75637 31961 75671 31989
rect 75699 31961 84485 31989
rect 84513 31961 84547 31989
rect 84575 31961 84609 31989
rect 84637 31961 84671 31989
rect 84699 31961 93485 31989
rect 93513 31961 93547 31989
rect 93575 31961 93609 31989
rect 93637 31961 93671 31989
rect 93699 31961 102485 31989
rect 102513 31961 102547 31989
rect 102575 31961 102609 31989
rect 102637 31961 102671 31989
rect 102699 31961 111485 31989
rect 111513 31961 111547 31989
rect 111575 31961 111609 31989
rect 111637 31961 111671 31989
rect 111699 31961 120485 31989
rect 120513 31961 120547 31989
rect 120575 31961 120609 31989
rect 120637 31961 120671 31989
rect 120699 31961 129485 31989
rect 129513 31961 129547 31989
rect 129575 31961 129609 31989
rect 129637 31961 129671 31989
rect 129699 31961 138485 31989
rect 138513 31961 138547 31989
rect 138575 31961 138609 31989
rect 138637 31961 138671 31989
rect 138699 31961 147485 31989
rect 147513 31961 147547 31989
rect 147575 31961 147609 31989
rect 147637 31961 147671 31989
rect 147699 31961 156485 31989
rect 156513 31961 156547 31989
rect 156575 31961 156609 31989
rect 156637 31961 156671 31989
rect 156699 31961 165485 31989
rect 165513 31961 165547 31989
rect 165575 31961 165609 31989
rect 165637 31961 165671 31989
rect 165699 31961 174485 31989
rect 174513 31961 174547 31989
rect 174575 31961 174609 31989
rect 174637 31961 174671 31989
rect 174699 31961 183485 31989
rect 183513 31961 183547 31989
rect 183575 31961 183609 31989
rect 183637 31961 183671 31989
rect 183699 31961 192485 31989
rect 192513 31961 192547 31989
rect 192575 31961 192609 31989
rect 192637 31961 192671 31989
rect 192699 31961 201485 31989
rect 201513 31961 201547 31989
rect 201575 31961 201609 31989
rect 201637 31961 201671 31989
rect 201699 31961 210485 31989
rect 210513 31961 210547 31989
rect 210575 31961 210609 31989
rect 210637 31961 210671 31989
rect 210699 31961 219485 31989
rect 219513 31961 219547 31989
rect 219575 31961 219609 31989
rect 219637 31961 219671 31989
rect 219699 31961 228485 31989
rect 228513 31961 228547 31989
rect 228575 31961 228609 31989
rect 228637 31961 228671 31989
rect 228699 31961 237485 31989
rect 237513 31961 237547 31989
rect 237575 31961 237609 31989
rect 237637 31961 237671 31989
rect 237699 31961 246485 31989
rect 246513 31961 246547 31989
rect 246575 31961 246609 31989
rect 246637 31961 246671 31989
rect 246699 31961 255485 31989
rect 255513 31961 255547 31989
rect 255575 31961 255609 31989
rect 255637 31961 255671 31989
rect 255699 31961 264485 31989
rect 264513 31961 264547 31989
rect 264575 31961 264609 31989
rect 264637 31961 264671 31989
rect 264699 31961 273485 31989
rect 273513 31961 273547 31989
rect 273575 31961 273609 31989
rect 273637 31961 273671 31989
rect 273699 31961 282485 31989
rect 282513 31961 282547 31989
rect 282575 31961 282609 31989
rect 282637 31961 282671 31989
rect 282699 31961 291485 31989
rect 291513 31961 291547 31989
rect 291575 31961 291609 31989
rect 291637 31961 291671 31989
rect 291699 31961 298728 31989
rect 298756 31961 298790 31989
rect 298818 31961 298852 31989
rect 298880 31961 298914 31989
rect 298942 31961 298990 31989
rect -958 31913 298990 31961
rect -958 29175 298990 29223
rect -958 29147 -430 29175
rect -402 29147 -368 29175
rect -340 29147 -306 29175
rect -278 29147 -244 29175
rect -216 29147 1625 29175
rect 1653 29147 1687 29175
rect 1715 29147 1749 29175
rect 1777 29147 1811 29175
rect 1839 29147 10625 29175
rect 10653 29147 10687 29175
rect 10715 29147 10749 29175
rect 10777 29147 10811 29175
rect 10839 29147 19625 29175
rect 19653 29147 19687 29175
rect 19715 29147 19749 29175
rect 19777 29147 19811 29175
rect 19839 29147 28625 29175
rect 28653 29147 28687 29175
rect 28715 29147 28749 29175
rect 28777 29147 28811 29175
rect 28839 29147 37625 29175
rect 37653 29147 37687 29175
rect 37715 29147 37749 29175
rect 37777 29147 37811 29175
rect 37839 29147 46625 29175
rect 46653 29147 46687 29175
rect 46715 29147 46749 29175
rect 46777 29147 46811 29175
rect 46839 29147 55625 29175
rect 55653 29147 55687 29175
rect 55715 29147 55749 29175
rect 55777 29147 55811 29175
rect 55839 29147 64625 29175
rect 64653 29147 64687 29175
rect 64715 29147 64749 29175
rect 64777 29147 64811 29175
rect 64839 29147 73625 29175
rect 73653 29147 73687 29175
rect 73715 29147 73749 29175
rect 73777 29147 73811 29175
rect 73839 29147 82625 29175
rect 82653 29147 82687 29175
rect 82715 29147 82749 29175
rect 82777 29147 82811 29175
rect 82839 29147 91625 29175
rect 91653 29147 91687 29175
rect 91715 29147 91749 29175
rect 91777 29147 91811 29175
rect 91839 29147 100625 29175
rect 100653 29147 100687 29175
rect 100715 29147 100749 29175
rect 100777 29147 100811 29175
rect 100839 29147 109625 29175
rect 109653 29147 109687 29175
rect 109715 29147 109749 29175
rect 109777 29147 109811 29175
rect 109839 29147 118625 29175
rect 118653 29147 118687 29175
rect 118715 29147 118749 29175
rect 118777 29147 118811 29175
rect 118839 29147 127625 29175
rect 127653 29147 127687 29175
rect 127715 29147 127749 29175
rect 127777 29147 127811 29175
rect 127839 29147 136625 29175
rect 136653 29147 136687 29175
rect 136715 29147 136749 29175
rect 136777 29147 136811 29175
rect 136839 29147 145625 29175
rect 145653 29147 145687 29175
rect 145715 29147 145749 29175
rect 145777 29147 145811 29175
rect 145839 29147 154625 29175
rect 154653 29147 154687 29175
rect 154715 29147 154749 29175
rect 154777 29147 154811 29175
rect 154839 29147 163625 29175
rect 163653 29147 163687 29175
rect 163715 29147 163749 29175
rect 163777 29147 163811 29175
rect 163839 29147 172625 29175
rect 172653 29147 172687 29175
rect 172715 29147 172749 29175
rect 172777 29147 172811 29175
rect 172839 29147 181625 29175
rect 181653 29147 181687 29175
rect 181715 29147 181749 29175
rect 181777 29147 181811 29175
rect 181839 29147 190625 29175
rect 190653 29147 190687 29175
rect 190715 29147 190749 29175
rect 190777 29147 190811 29175
rect 190839 29147 199625 29175
rect 199653 29147 199687 29175
rect 199715 29147 199749 29175
rect 199777 29147 199811 29175
rect 199839 29147 208625 29175
rect 208653 29147 208687 29175
rect 208715 29147 208749 29175
rect 208777 29147 208811 29175
rect 208839 29147 217625 29175
rect 217653 29147 217687 29175
rect 217715 29147 217749 29175
rect 217777 29147 217811 29175
rect 217839 29147 226625 29175
rect 226653 29147 226687 29175
rect 226715 29147 226749 29175
rect 226777 29147 226811 29175
rect 226839 29147 235625 29175
rect 235653 29147 235687 29175
rect 235715 29147 235749 29175
rect 235777 29147 235811 29175
rect 235839 29147 244625 29175
rect 244653 29147 244687 29175
rect 244715 29147 244749 29175
rect 244777 29147 244811 29175
rect 244839 29147 253625 29175
rect 253653 29147 253687 29175
rect 253715 29147 253749 29175
rect 253777 29147 253811 29175
rect 253839 29147 262625 29175
rect 262653 29147 262687 29175
rect 262715 29147 262749 29175
rect 262777 29147 262811 29175
rect 262839 29147 271625 29175
rect 271653 29147 271687 29175
rect 271715 29147 271749 29175
rect 271777 29147 271811 29175
rect 271839 29147 280625 29175
rect 280653 29147 280687 29175
rect 280715 29147 280749 29175
rect 280777 29147 280811 29175
rect 280839 29147 289625 29175
rect 289653 29147 289687 29175
rect 289715 29147 289749 29175
rect 289777 29147 289811 29175
rect 289839 29147 298248 29175
rect 298276 29147 298310 29175
rect 298338 29147 298372 29175
rect 298400 29147 298434 29175
rect 298462 29147 298990 29175
rect -958 29113 298990 29147
rect -958 29085 -430 29113
rect -402 29085 -368 29113
rect -340 29085 -306 29113
rect -278 29085 -244 29113
rect -216 29085 1625 29113
rect 1653 29085 1687 29113
rect 1715 29085 1749 29113
rect 1777 29085 1811 29113
rect 1839 29085 10625 29113
rect 10653 29085 10687 29113
rect 10715 29085 10749 29113
rect 10777 29085 10811 29113
rect 10839 29085 19625 29113
rect 19653 29085 19687 29113
rect 19715 29085 19749 29113
rect 19777 29085 19811 29113
rect 19839 29085 28625 29113
rect 28653 29085 28687 29113
rect 28715 29085 28749 29113
rect 28777 29085 28811 29113
rect 28839 29085 37625 29113
rect 37653 29085 37687 29113
rect 37715 29085 37749 29113
rect 37777 29085 37811 29113
rect 37839 29085 46625 29113
rect 46653 29085 46687 29113
rect 46715 29085 46749 29113
rect 46777 29085 46811 29113
rect 46839 29085 55625 29113
rect 55653 29085 55687 29113
rect 55715 29085 55749 29113
rect 55777 29085 55811 29113
rect 55839 29085 64625 29113
rect 64653 29085 64687 29113
rect 64715 29085 64749 29113
rect 64777 29085 64811 29113
rect 64839 29085 73625 29113
rect 73653 29085 73687 29113
rect 73715 29085 73749 29113
rect 73777 29085 73811 29113
rect 73839 29085 82625 29113
rect 82653 29085 82687 29113
rect 82715 29085 82749 29113
rect 82777 29085 82811 29113
rect 82839 29085 91625 29113
rect 91653 29085 91687 29113
rect 91715 29085 91749 29113
rect 91777 29085 91811 29113
rect 91839 29085 100625 29113
rect 100653 29085 100687 29113
rect 100715 29085 100749 29113
rect 100777 29085 100811 29113
rect 100839 29085 109625 29113
rect 109653 29085 109687 29113
rect 109715 29085 109749 29113
rect 109777 29085 109811 29113
rect 109839 29085 118625 29113
rect 118653 29085 118687 29113
rect 118715 29085 118749 29113
rect 118777 29085 118811 29113
rect 118839 29085 127625 29113
rect 127653 29085 127687 29113
rect 127715 29085 127749 29113
rect 127777 29085 127811 29113
rect 127839 29085 136625 29113
rect 136653 29085 136687 29113
rect 136715 29085 136749 29113
rect 136777 29085 136811 29113
rect 136839 29085 145625 29113
rect 145653 29085 145687 29113
rect 145715 29085 145749 29113
rect 145777 29085 145811 29113
rect 145839 29085 154625 29113
rect 154653 29085 154687 29113
rect 154715 29085 154749 29113
rect 154777 29085 154811 29113
rect 154839 29085 163625 29113
rect 163653 29085 163687 29113
rect 163715 29085 163749 29113
rect 163777 29085 163811 29113
rect 163839 29085 172625 29113
rect 172653 29085 172687 29113
rect 172715 29085 172749 29113
rect 172777 29085 172811 29113
rect 172839 29085 181625 29113
rect 181653 29085 181687 29113
rect 181715 29085 181749 29113
rect 181777 29085 181811 29113
rect 181839 29085 190625 29113
rect 190653 29085 190687 29113
rect 190715 29085 190749 29113
rect 190777 29085 190811 29113
rect 190839 29085 199625 29113
rect 199653 29085 199687 29113
rect 199715 29085 199749 29113
rect 199777 29085 199811 29113
rect 199839 29085 208625 29113
rect 208653 29085 208687 29113
rect 208715 29085 208749 29113
rect 208777 29085 208811 29113
rect 208839 29085 217625 29113
rect 217653 29085 217687 29113
rect 217715 29085 217749 29113
rect 217777 29085 217811 29113
rect 217839 29085 226625 29113
rect 226653 29085 226687 29113
rect 226715 29085 226749 29113
rect 226777 29085 226811 29113
rect 226839 29085 235625 29113
rect 235653 29085 235687 29113
rect 235715 29085 235749 29113
rect 235777 29085 235811 29113
rect 235839 29085 244625 29113
rect 244653 29085 244687 29113
rect 244715 29085 244749 29113
rect 244777 29085 244811 29113
rect 244839 29085 253625 29113
rect 253653 29085 253687 29113
rect 253715 29085 253749 29113
rect 253777 29085 253811 29113
rect 253839 29085 262625 29113
rect 262653 29085 262687 29113
rect 262715 29085 262749 29113
rect 262777 29085 262811 29113
rect 262839 29085 271625 29113
rect 271653 29085 271687 29113
rect 271715 29085 271749 29113
rect 271777 29085 271811 29113
rect 271839 29085 280625 29113
rect 280653 29085 280687 29113
rect 280715 29085 280749 29113
rect 280777 29085 280811 29113
rect 280839 29085 289625 29113
rect 289653 29085 289687 29113
rect 289715 29085 289749 29113
rect 289777 29085 289811 29113
rect 289839 29085 298248 29113
rect 298276 29085 298310 29113
rect 298338 29085 298372 29113
rect 298400 29085 298434 29113
rect 298462 29085 298990 29113
rect -958 29051 298990 29085
rect -958 29023 -430 29051
rect -402 29023 -368 29051
rect -340 29023 -306 29051
rect -278 29023 -244 29051
rect -216 29023 1625 29051
rect 1653 29023 1687 29051
rect 1715 29023 1749 29051
rect 1777 29023 1811 29051
rect 1839 29023 10625 29051
rect 10653 29023 10687 29051
rect 10715 29023 10749 29051
rect 10777 29023 10811 29051
rect 10839 29023 19625 29051
rect 19653 29023 19687 29051
rect 19715 29023 19749 29051
rect 19777 29023 19811 29051
rect 19839 29023 28625 29051
rect 28653 29023 28687 29051
rect 28715 29023 28749 29051
rect 28777 29023 28811 29051
rect 28839 29023 37625 29051
rect 37653 29023 37687 29051
rect 37715 29023 37749 29051
rect 37777 29023 37811 29051
rect 37839 29023 46625 29051
rect 46653 29023 46687 29051
rect 46715 29023 46749 29051
rect 46777 29023 46811 29051
rect 46839 29023 55625 29051
rect 55653 29023 55687 29051
rect 55715 29023 55749 29051
rect 55777 29023 55811 29051
rect 55839 29023 64625 29051
rect 64653 29023 64687 29051
rect 64715 29023 64749 29051
rect 64777 29023 64811 29051
rect 64839 29023 73625 29051
rect 73653 29023 73687 29051
rect 73715 29023 73749 29051
rect 73777 29023 73811 29051
rect 73839 29023 82625 29051
rect 82653 29023 82687 29051
rect 82715 29023 82749 29051
rect 82777 29023 82811 29051
rect 82839 29023 91625 29051
rect 91653 29023 91687 29051
rect 91715 29023 91749 29051
rect 91777 29023 91811 29051
rect 91839 29023 100625 29051
rect 100653 29023 100687 29051
rect 100715 29023 100749 29051
rect 100777 29023 100811 29051
rect 100839 29023 109625 29051
rect 109653 29023 109687 29051
rect 109715 29023 109749 29051
rect 109777 29023 109811 29051
rect 109839 29023 118625 29051
rect 118653 29023 118687 29051
rect 118715 29023 118749 29051
rect 118777 29023 118811 29051
rect 118839 29023 127625 29051
rect 127653 29023 127687 29051
rect 127715 29023 127749 29051
rect 127777 29023 127811 29051
rect 127839 29023 136625 29051
rect 136653 29023 136687 29051
rect 136715 29023 136749 29051
rect 136777 29023 136811 29051
rect 136839 29023 145625 29051
rect 145653 29023 145687 29051
rect 145715 29023 145749 29051
rect 145777 29023 145811 29051
rect 145839 29023 154625 29051
rect 154653 29023 154687 29051
rect 154715 29023 154749 29051
rect 154777 29023 154811 29051
rect 154839 29023 163625 29051
rect 163653 29023 163687 29051
rect 163715 29023 163749 29051
rect 163777 29023 163811 29051
rect 163839 29023 172625 29051
rect 172653 29023 172687 29051
rect 172715 29023 172749 29051
rect 172777 29023 172811 29051
rect 172839 29023 181625 29051
rect 181653 29023 181687 29051
rect 181715 29023 181749 29051
rect 181777 29023 181811 29051
rect 181839 29023 190625 29051
rect 190653 29023 190687 29051
rect 190715 29023 190749 29051
rect 190777 29023 190811 29051
rect 190839 29023 199625 29051
rect 199653 29023 199687 29051
rect 199715 29023 199749 29051
rect 199777 29023 199811 29051
rect 199839 29023 208625 29051
rect 208653 29023 208687 29051
rect 208715 29023 208749 29051
rect 208777 29023 208811 29051
rect 208839 29023 217625 29051
rect 217653 29023 217687 29051
rect 217715 29023 217749 29051
rect 217777 29023 217811 29051
rect 217839 29023 226625 29051
rect 226653 29023 226687 29051
rect 226715 29023 226749 29051
rect 226777 29023 226811 29051
rect 226839 29023 235625 29051
rect 235653 29023 235687 29051
rect 235715 29023 235749 29051
rect 235777 29023 235811 29051
rect 235839 29023 244625 29051
rect 244653 29023 244687 29051
rect 244715 29023 244749 29051
rect 244777 29023 244811 29051
rect 244839 29023 253625 29051
rect 253653 29023 253687 29051
rect 253715 29023 253749 29051
rect 253777 29023 253811 29051
rect 253839 29023 262625 29051
rect 262653 29023 262687 29051
rect 262715 29023 262749 29051
rect 262777 29023 262811 29051
rect 262839 29023 271625 29051
rect 271653 29023 271687 29051
rect 271715 29023 271749 29051
rect 271777 29023 271811 29051
rect 271839 29023 280625 29051
rect 280653 29023 280687 29051
rect 280715 29023 280749 29051
rect 280777 29023 280811 29051
rect 280839 29023 289625 29051
rect 289653 29023 289687 29051
rect 289715 29023 289749 29051
rect 289777 29023 289811 29051
rect 289839 29023 298248 29051
rect 298276 29023 298310 29051
rect 298338 29023 298372 29051
rect 298400 29023 298434 29051
rect 298462 29023 298990 29051
rect -958 28989 298990 29023
rect -958 28961 -430 28989
rect -402 28961 -368 28989
rect -340 28961 -306 28989
rect -278 28961 -244 28989
rect -216 28961 1625 28989
rect 1653 28961 1687 28989
rect 1715 28961 1749 28989
rect 1777 28961 1811 28989
rect 1839 28961 10625 28989
rect 10653 28961 10687 28989
rect 10715 28961 10749 28989
rect 10777 28961 10811 28989
rect 10839 28961 19625 28989
rect 19653 28961 19687 28989
rect 19715 28961 19749 28989
rect 19777 28961 19811 28989
rect 19839 28961 28625 28989
rect 28653 28961 28687 28989
rect 28715 28961 28749 28989
rect 28777 28961 28811 28989
rect 28839 28961 37625 28989
rect 37653 28961 37687 28989
rect 37715 28961 37749 28989
rect 37777 28961 37811 28989
rect 37839 28961 46625 28989
rect 46653 28961 46687 28989
rect 46715 28961 46749 28989
rect 46777 28961 46811 28989
rect 46839 28961 55625 28989
rect 55653 28961 55687 28989
rect 55715 28961 55749 28989
rect 55777 28961 55811 28989
rect 55839 28961 64625 28989
rect 64653 28961 64687 28989
rect 64715 28961 64749 28989
rect 64777 28961 64811 28989
rect 64839 28961 73625 28989
rect 73653 28961 73687 28989
rect 73715 28961 73749 28989
rect 73777 28961 73811 28989
rect 73839 28961 82625 28989
rect 82653 28961 82687 28989
rect 82715 28961 82749 28989
rect 82777 28961 82811 28989
rect 82839 28961 91625 28989
rect 91653 28961 91687 28989
rect 91715 28961 91749 28989
rect 91777 28961 91811 28989
rect 91839 28961 100625 28989
rect 100653 28961 100687 28989
rect 100715 28961 100749 28989
rect 100777 28961 100811 28989
rect 100839 28961 109625 28989
rect 109653 28961 109687 28989
rect 109715 28961 109749 28989
rect 109777 28961 109811 28989
rect 109839 28961 118625 28989
rect 118653 28961 118687 28989
rect 118715 28961 118749 28989
rect 118777 28961 118811 28989
rect 118839 28961 127625 28989
rect 127653 28961 127687 28989
rect 127715 28961 127749 28989
rect 127777 28961 127811 28989
rect 127839 28961 136625 28989
rect 136653 28961 136687 28989
rect 136715 28961 136749 28989
rect 136777 28961 136811 28989
rect 136839 28961 145625 28989
rect 145653 28961 145687 28989
rect 145715 28961 145749 28989
rect 145777 28961 145811 28989
rect 145839 28961 154625 28989
rect 154653 28961 154687 28989
rect 154715 28961 154749 28989
rect 154777 28961 154811 28989
rect 154839 28961 163625 28989
rect 163653 28961 163687 28989
rect 163715 28961 163749 28989
rect 163777 28961 163811 28989
rect 163839 28961 172625 28989
rect 172653 28961 172687 28989
rect 172715 28961 172749 28989
rect 172777 28961 172811 28989
rect 172839 28961 181625 28989
rect 181653 28961 181687 28989
rect 181715 28961 181749 28989
rect 181777 28961 181811 28989
rect 181839 28961 190625 28989
rect 190653 28961 190687 28989
rect 190715 28961 190749 28989
rect 190777 28961 190811 28989
rect 190839 28961 199625 28989
rect 199653 28961 199687 28989
rect 199715 28961 199749 28989
rect 199777 28961 199811 28989
rect 199839 28961 208625 28989
rect 208653 28961 208687 28989
rect 208715 28961 208749 28989
rect 208777 28961 208811 28989
rect 208839 28961 217625 28989
rect 217653 28961 217687 28989
rect 217715 28961 217749 28989
rect 217777 28961 217811 28989
rect 217839 28961 226625 28989
rect 226653 28961 226687 28989
rect 226715 28961 226749 28989
rect 226777 28961 226811 28989
rect 226839 28961 235625 28989
rect 235653 28961 235687 28989
rect 235715 28961 235749 28989
rect 235777 28961 235811 28989
rect 235839 28961 244625 28989
rect 244653 28961 244687 28989
rect 244715 28961 244749 28989
rect 244777 28961 244811 28989
rect 244839 28961 253625 28989
rect 253653 28961 253687 28989
rect 253715 28961 253749 28989
rect 253777 28961 253811 28989
rect 253839 28961 262625 28989
rect 262653 28961 262687 28989
rect 262715 28961 262749 28989
rect 262777 28961 262811 28989
rect 262839 28961 271625 28989
rect 271653 28961 271687 28989
rect 271715 28961 271749 28989
rect 271777 28961 271811 28989
rect 271839 28961 280625 28989
rect 280653 28961 280687 28989
rect 280715 28961 280749 28989
rect 280777 28961 280811 28989
rect 280839 28961 289625 28989
rect 289653 28961 289687 28989
rect 289715 28961 289749 28989
rect 289777 28961 289811 28989
rect 289839 28961 298248 28989
rect 298276 28961 298310 28989
rect 298338 28961 298372 28989
rect 298400 28961 298434 28989
rect 298462 28961 298990 28989
rect -958 28913 298990 28961
rect -958 23175 298990 23223
rect -958 23147 -910 23175
rect -882 23147 -848 23175
rect -820 23147 -786 23175
rect -758 23147 -724 23175
rect -696 23147 3485 23175
rect 3513 23147 3547 23175
rect 3575 23147 3609 23175
rect 3637 23147 3671 23175
rect 3699 23147 12485 23175
rect 12513 23147 12547 23175
rect 12575 23147 12609 23175
rect 12637 23147 12671 23175
rect 12699 23147 21485 23175
rect 21513 23147 21547 23175
rect 21575 23147 21609 23175
rect 21637 23147 21671 23175
rect 21699 23147 30485 23175
rect 30513 23147 30547 23175
rect 30575 23147 30609 23175
rect 30637 23147 30671 23175
rect 30699 23147 39485 23175
rect 39513 23147 39547 23175
rect 39575 23147 39609 23175
rect 39637 23147 39671 23175
rect 39699 23147 48485 23175
rect 48513 23147 48547 23175
rect 48575 23147 48609 23175
rect 48637 23147 48671 23175
rect 48699 23147 57485 23175
rect 57513 23147 57547 23175
rect 57575 23147 57609 23175
rect 57637 23147 57671 23175
rect 57699 23147 66485 23175
rect 66513 23147 66547 23175
rect 66575 23147 66609 23175
rect 66637 23147 66671 23175
rect 66699 23147 75485 23175
rect 75513 23147 75547 23175
rect 75575 23147 75609 23175
rect 75637 23147 75671 23175
rect 75699 23147 84485 23175
rect 84513 23147 84547 23175
rect 84575 23147 84609 23175
rect 84637 23147 84671 23175
rect 84699 23147 93485 23175
rect 93513 23147 93547 23175
rect 93575 23147 93609 23175
rect 93637 23147 93671 23175
rect 93699 23147 102485 23175
rect 102513 23147 102547 23175
rect 102575 23147 102609 23175
rect 102637 23147 102671 23175
rect 102699 23147 111485 23175
rect 111513 23147 111547 23175
rect 111575 23147 111609 23175
rect 111637 23147 111671 23175
rect 111699 23147 120485 23175
rect 120513 23147 120547 23175
rect 120575 23147 120609 23175
rect 120637 23147 120671 23175
rect 120699 23147 129485 23175
rect 129513 23147 129547 23175
rect 129575 23147 129609 23175
rect 129637 23147 129671 23175
rect 129699 23147 138485 23175
rect 138513 23147 138547 23175
rect 138575 23147 138609 23175
rect 138637 23147 138671 23175
rect 138699 23147 147485 23175
rect 147513 23147 147547 23175
rect 147575 23147 147609 23175
rect 147637 23147 147671 23175
rect 147699 23147 156485 23175
rect 156513 23147 156547 23175
rect 156575 23147 156609 23175
rect 156637 23147 156671 23175
rect 156699 23147 165485 23175
rect 165513 23147 165547 23175
rect 165575 23147 165609 23175
rect 165637 23147 165671 23175
rect 165699 23147 174485 23175
rect 174513 23147 174547 23175
rect 174575 23147 174609 23175
rect 174637 23147 174671 23175
rect 174699 23147 183485 23175
rect 183513 23147 183547 23175
rect 183575 23147 183609 23175
rect 183637 23147 183671 23175
rect 183699 23147 192485 23175
rect 192513 23147 192547 23175
rect 192575 23147 192609 23175
rect 192637 23147 192671 23175
rect 192699 23147 201485 23175
rect 201513 23147 201547 23175
rect 201575 23147 201609 23175
rect 201637 23147 201671 23175
rect 201699 23147 210485 23175
rect 210513 23147 210547 23175
rect 210575 23147 210609 23175
rect 210637 23147 210671 23175
rect 210699 23147 219485 23175
rect 219513 23147 219547 23175
rect 219575 23147 219609 23175
rect 219637 23147 219671 23175
rect 219699 23147 228485 23175
rect 228513 23147 228547 23175
rect 228575 23147 228609 23175
rect 228637 23147 228671 23175
rect 228699 23147 237485 23175
rect 237513 23147 237547 23175
rect 237575 23147 237609 23175
rect 237637 23147 237671 23175
rect 237699 23147 246485 23175
rect 246513 23147 246547 23175
rect 246575 23147 246609 23175
rect 246637 23147 246671 23175
rect 246699 23147 255485 23175
rect 255513 23147 255547 23175
rect 255575 23147 255609 23175
rect 255637 23147 255671 23175
rect 255699 23147 264485 23175
rect 264513 23147 264547 23175
rect 264575 23147 264609 23175
rect 264637 23147 264671 23175
rect 264699 23147 273485 23175
rect 273513 23147 273547 23175
rect 273575 23147 273609 23175
rect 273637 23147 273671 23175
rect 273699 23147 282485 23175
rect 282513 23147 282547 23175
rect 282575 23147 282609 23175
rect 282637 23147 282671 23175
rect 282699 23147 291485 23175
rect 291513 23147 291547 23175
rect 291575 23147 291609 23175
rect 291637 23147 291671 23175
rect 291699 23147 298728 23175
rect 298756 23147 298790 23175
rect 298818 23147 298852 23175
rect 298880 23147 298914 23175
rect 298942 23147 298990 23175
rect -958 23113 298990 23147
rect -958 23085 -910 23113
rect -882 23085 -848 23113
rect -820 23085 -786 23113
rect -758 23085 -724 23113
rect -696 23085 3485 23113
rect 3513 23085 3547 23113
rect 3575 23085 3609 23113
rect 3637 23085 3671 23113
rect 3699 23085 12485 23113
rect 12513 23085 12547 23113
rect 12575 23085 12609 23113
rect 12637 23085 12671 23113
rect 12699 23085 21485 23113
rect 21513 23085 21547 23113
rect 21575 23085 21609 23113
rect 21637 23085 21671 23113
rect 21699 23085 30485 23113
rect 30513 23085 30547 23113
rect 30575 23085 30609 23113
rect 30637 23085 30671 23113
rect 30699 23085 39485 23113
rect 39513 23085 39547 23113
rect 39575 23085 39609 23113
rect 39637 23085 39671 23113
rect 39699 23085 48485 23113
rect 48513 23085 48547 23113
rect 48575 23085 48609 23113
rect 48637 23085 48671 23113
rect 48699 23085 57485 23113
rect 57513 23085 57547 23113
rect 57575 23085 57609 23113
rect 57637 23085 57671 23113
rect 57699 23085 66485 23113
rect 66513 23085 66547 23113
rect 66575 23085 66609 23113
rect 66637 23085 66671 23113
rect 66699 23085 75485 23113
rect 75513 23085 75547 23113
rect 75575 23085 75609 23113
rect 75637 23085 75671 23113
rect 75699 23085 84485 23113
rect 84513 23085 84547 23113
rect 84575 23085 84609 23113
rect 84637 23085 84671 23113
rect 84699 23085 93485 23113
rect 93513 23085 93547 23113
rect 93575 23085 93609 23113
rect 93637 23085 93671 23113
rect 93699 23085 102485 23113
rect 102513 23085 102547 23113
rect 102575 23085 102609 23113
rect 102637 23085 102671 23113
rect 102699 23085 111485 23113
rect 111513 23085 111547 23113
rect 111575 23085 111609 23113
rect 111637 23085 111671 23113
rect 111699 23085 120485 23113
rect 120513 23085 120547 23113
rect 120575 23085 120609 23113
rect 120637 23085 120671 23113
rect 120699 23085 129485 23113
rect 129513 23085 129547 23113
rect 129575 23085 129609 23113
rect 129637 23085 129671 23113
rect 129699 23085 138485 23113
rect 138513 23085 138547 23113
rect 138575 23085 138609 23113
rect 138637 23085 138671 23113
rect 138699 23085 147485 23113
rect 147513 23085 147547 23113
rect 147575 23085 147609 23113
rect 147637 23085 147671 23113
rect 147699 23085 156485 23113
rect 156513 23085 156547 23113
rect 156575 23085 156609 23113
rect 156637 23085 156671 23113
rect 156699 23085 165485 23113
rect 165513 23085 165547 23113
rect 165575 23085 165609 23113
rect 165637 23085 165671 23113
rect 165699 23085 174485 23113
rect 174513 23085 174547 23113
rect 174575 23085 174609 23113
rect 174637 23085 174671 23113
rect 174699 23085 183485 23113
rect 183513 23085 183547 23113
rect 183575 23085 183609 23113
rect 183637 23085 183671 23113
rect 183699 23085 192485 23113
rect 192513 23085 192547 23113
rect 192575 23085 192609 23113
rect 192637 23085 192671 23113
rect 192699 23085 201485 23113
rect 201513 23085 201547 23113
rect 201575 23085 201609 23113
rect 201637 23085 201671 23113
rect 201699 23085 210485 23113
rect 210513 23085 210547 23113
rect 210575 23085 210609 23113
rect 210637 23085 210671 23113
rect 210699 23085 219485 23113
rect 219513 23085 219547 23113
rect 219575 23085 219609 23113
rect 219637 23085 219671 23113
rect 219699 23085 228485 23113
rect 228513 23085 228547 23113
rect 228575 23085 228609 23113
rect 228637 23085 228671 23113
rect 228699 23085 237485 23113
rect 237513 23085 237547 23113
rect 237575 23085 237609 23113
rect 237637 23085 237671 23113
rect 237699 23085 246485 23113
rect 246513 23085 246547 23113
rect 246575 23085 246609 23113
rect 246637 23085 246671 23113
rect 246699 23085 255485 23113
rect 255513 23085 255547 23113
rect 255575 23085 255609 23113
rect 255637 23085 255671 23113
rect 255699 23085 264485 23113
rect 264513 23085 264547 23113
rect 264575 23085 264609 23113
rect 264637 23085 264671 23113
rect 264699 23085 273485 23113
rect 273513 23085 273547 23113
rect 273575 23085 273609 23113
rect 273637 23085 273671 23113
rect 273699 23085 282485 23113
rect 282513 23085 282547 23113
rect 282575 23085 282609 23113
rect 282637 23085 282671 23113
rect 282699 23085 291485 23113
rect 291513 23085 291547 23113
rect 291575 23085 291609 23113
rect 291637 23085 291671 23113
rect 291699 23085 298728 23113
rect 298756 23085 298790 23113
rect 298818 23085 298852 23113
rect 298880 23085 298914 23113
rect 298942 23085 298990 23113
rect -958 23051 298990 23085
rect -958 23023 -910 23051
rect -882 23023 -848 23051
rect -820 23023 -786 23051
rect -758 23023 -724 23051
rect -696 23023 3485 23051
rect 3513 23023 3547 23051
rect 3575 23023 3609 23051
rect 3637 23023 3671 23051
rect 3699 23023 12485 23051
rect 12513 23023 12547 23051
rect 12575 23023 12609 23051
rect 12637 23023 12671 23051
rect 12699 23023 21485 23051
rect 21513 23023 21547 23051
rect 21575 23023 21609 23051
rect 21637 23023 21671 23051
rect 21699 23023 30485 23051
rect 30513 23023 30547 23051
rect 30575 23023 30609 23051
rect 30637 23023 30671 23051
rect 30699 23023 39485 23051
rect 39513 23023 39547 23051
rect 39575 23023 39609 23051
rect 39637 23023 39671 23051
rect 39699 23023 48485 23051
rect 48513 23023 48547 23051
rect 48575 23023 48609 23051
rect 48637 23023 48671 23051
rect 48699 23023 57485 23051
rect 57513 23023 57547 23051
rect 57575 23023 57609 23051
rect 57637 23023 57671 23051
rect 57699 23023 66485 23051
rect 66513 23023 66547 23051
rect 66575 23023 66609 23051
rect 66637 23023 66671 23051
rect 66699 23023 75485 23051
rect 75513 23023 75547 23051
rect 75575 23023 75609 23051
rect 75637 23023 75671 23051
rect 75699 23023 84485 23051
rect 84513 23023 84547 23051
rect 84575 23023 84609 23051
rect 84637 23023 84671 23051
rect 84699 23023 93485 23051
rect 93513 23023 93547 23051
rect 93575 23023 93609 23051
rect 93637 23023 93671 23051
rect 93699 23023 102485 23051
rect 102513 23023 102547 23051
rect 102575 23023 102609 23051
rect 102637 23023 102671 23051
rect 102699 23023 111485 23051
rect 111513 23023 111547 23051
rect 111575 23023 111609 23051
rect 111637 23023 111671 23051
rect 111699 23023 120485 23051
rect 120513 23023 120547 23051
rect 120575 23023 120609 23051
rect 120637 23023 120671 23051
rect 120699 23023 129485 23051
rect 129513 23023 129547 23051
rect 129575 23023 129609 23051
rect 129637 23023 129671 23051
rect 129699 23023 138485 23051
rect 138513 23023 138547 23051
rect 138575 23023 138609 23051
rect 138637 23023 138671 23051
rect 138699 23023 147485 23051
rect 147513 23023 147547 23051
rect 147575 23023 147609 23051
rect 147637 23023 147671 23051
rect 147699 23023 156485 23051
rect 156513 23023 156547 23051
rect 156575 23023 156609 23051
rect 156637 23023 156671 23051
rect 156699 23023 165485 23051
rect 165513 23023 165547 23051
rect 165575 23023 165609 23051
rect 165637 23023 165671 23051
rect 165699 23023 174485 23051
rect 174513 23023 174547 23051
rect 174575 23023 174609 23051
rect 174637 23023 174671 23051
rect 174699 23023 183485 23051
rect 183513 23023 183547 23051
rect 183575 23023 183609 23051
rect 183637 23023 183671 23051
rect 183699 23023 192485 23051
rect 192513 23023 192547 23051
rect 192575 23023 192609 23051
rect 192637 23023 192671 23051
rect 192699 23023 201485 23051
rect 201513 23023 201547 23051
rect 201575 23023 201609 23051
rect 201637 23023 201671 23051
rect 201699 23023 210485 23051
rect 210513 23023 210547 23051
rect 210575 23023 210609 23051
rect 210637 23023 210671 23051
rect 210699 23023 219485 23051
rect 219513 23023 219547 23051
rect 219575 23023 219609 23051
rect 219637 23023 219671 23051
rect 219699 23023 228485 23051
rect 228513 23023 228547 23051
rect 228575 23023 228609 23051
rect 228637 23023 228671 23051
rect 228699 23023 237485 23051
rect 237513 23023 237547 23051
rect 237575 23023 237609 23051
rect 237637 23023 237671 23051
rect 237699 23023 246485 23051
rect 246513 23023 246547 23051
rect 246575 23023 246609 23051
rect 246637 23023 246671 23051
rect 246699 23023 255485 23051
rect 255513 23023 255547 23051
rect 255575 23023 255609 23051
rect 255637 23023 255671 23051
rect 255699 23023 264485 23051
rect 264513 23023 264547 23051
rect 264575 23023 264609 23051
rect 264637 23023 264671 23051
rect 264699 23023 273485 23051
rect 273513 23023 273547 23051
rect 273575 23023 273609 23051
rect 273637 23023 273671 23051
rect 273699 23023 282485 23051
rect 282513 23023 282547 23051
rect 282575 23023 282609 23051
rect 282637 23023 282671 23051
rect 282699 23023 291485 23051
rect 291513 23023 291547 23051
rect 291575 23023 291609 23051
rect 291637 23023 291671 23051
rect 291699 23023 298728 23051
rect 298756 23023 298790 23051
rect 298818 23023 298852 23051
rect 298880 23023 298914 23051
rect 298942 23023 298990 23051
rect -958 22989 298990 23023
rect -958 22961 -910 22989
rect -882 22961 -848 22989
rect -820 22961 -786 22989
rect -758 22961 -724 22989
rect -696 22961 3485 22989
rect 3513 22961 3547 22989
rect 3575 22961 3609 22989
rect 3637 22961 3671 22989
rect 3699 22961 12485 22989
rect 12513 22961 12547 22989
rect 12575 22961 12609 22989
rect 12637 22961 12671 22989
rect 12699 22961 21485 22989
rect 21513 22961 21547 22989
rect 21575 22961 21609 22989
rect 21637 22961 21671 22989
rect 21699 22961 30485 22989
rect 30513 22961 30547 22989
rect 30575 22961 30609 22989
rect 30637 22961 30671 22989
rect 30699 22961 39485 22989
rect 39513 22961 39547 22989
rect 39575 22961 39609 22989
rect 39637 22961 39671 22989
rect 39699 22961 48485 22989
rect 48513 22961 48547 22989
rect 48575 22961 48609 22989
rect 48637 22961 48671 22989
rect 48699 22961 57485 22989
rect 57513 22961 57547 22989
rect 57575 22961 57609 22989
rect 57637 22961 57671 22989
rect 57699 22961 66485 22989
rect 66513 22961 66547 22989
rect 66575 22961 66609 22989
rect 66637 22961 66671 22989
rect 66699 22961 75485 22989
rect 75513 22961 75547 22989
rect 75575 22961 75609 22989
rect 75637 22961 75671 22989
rect 75699 22961 84485 22989
rect 84513 22961 84547 22989
rect 84575 22961 84609 22989
rect 84637 22961 84671 22989
rect 84699 22961 93485 22989
rect 93513 22961 93547 22989
rect 93575 22961 93609 22989
rect 93637 22961 93671 22989
rect 93699 22961 102485 22989
rect 102513 22961 102547 22989
rect 102575 22961 102609 22989
rect 102637 22961 102671 22989
rect 102699 22961 111485 22989
rect 111513 22961 111547 22989
rect 111575 22961 111609 22989
rect 111637 22961 111671 22989
rect 111699 22961 120485 22989
rect 120513 22961 120547 22989
rect 120575 22961 120609 22989
rect 120637 22961 120671 22989
rect 120699 22961 129485 22989
rect 129513 22961 129547 22989
rect 129575 22961 129609 22989
rect 129637 22961 129671 22989
rect 129699 22961 138485 22989
rect 138513 22961 138547 22989
rect 138575 22961 138609 22989
rect 138637 22961 138671 22989
rect 138699 22961 147485 22989
rect 147513 22961 147547 22989
rect 147575 22961 147609 22989
rect 147637 22961 147671 22989
rect 147699 22961 156485 22989
rect 156513 22961 156547 22989
rect 156575 22961 156609 22989
rect 156637 22961 156671 22989
rect 156699 22961 165485 22989
rect 165513 22961 165547 22989
rect 165575 22961 165609 22989
rect 165637 22961 165671 22989
rect 165699 22961 174485 22989
rect 174513 22961 174547 22989
rect 174575 22961 174609 22989
rect 174637 22961 174671 22989
rect 174699 22961 183485 22989
rect 183513 22961 183547 22989
rect 183575 22961 183609 22989
rect 183637 22961 183671 22989
rect 183699 22961 192485 22989
rect 192513 22961 192547 22989
rect 192575 22961 192609 22989
rect 192637 22961 192671 22989
rect 192699 22961 201485 22989
rect 201513 22961 201547 22989
rect 201575 22961 201609 22989
rect 201637 22961 201671 22989
rect 201699 22961 210485 22989
rect 210513 22961 210547 22989
rect 210575 22961 210609 22989
rect 210637 22961 210671 22989
rect 210699 22961 219485 22989
rect 219513 22961 219547 22989
rect 219575 22961 219609 22989
rect 219637 22961 219671 22989
rect 219699 22961 228485 22989
rect 228513 22961 228547 22989
rect 228575 22961 228609 22989
rect 228637 22961 228671 22989
rect 228699 22961 237485 22989
rect 237513 22961 237547 22989
rect 237575 22961 237609 22989
rect 237637 22961 237671 22989
rect 237699 22961 246485 22989
rect 246513 22961 246547 22989
rect 246575 22961 246609 22989
rect 246637 22961 246671 22989
rect 246699 22961 255485 22989
rect 255513 22961 255547 22989
rect 255575 22961 255609 22989
rect 255637 22961 255671 22989
rect 255699 22961 264485 22989
rect 264513 22961 264547 22989
rect 264575 22961 264609 22989
rect 264637 22961 264671 22989
rect 264699 22961 273485 22989
rect 273513 22961 273547 22989
rect 273575 22961 273609 22989
rect 273637 22961 273671 22989
rect 273699 22961 282485 22989
rect 282513 22961 282547 22989
rect 282575 22961 282609 22989
rect 282637 22961 282671 22989
rect 282699 22961 291485 22989
rect 291513 22961 291547 22989
rect 291575 22961 291609 22989
rect 291637 22961 291671 22989
rect 291699 22961 298728 22989
rect 298756 22961 298790 22989
rect 298818 22961 298852 22989
rect 298880 22961 298914 22989
rect 298942 22961 298990 22989
rect -958 22913 298990 22961
rect -958 20175 298990 20223
rect -958 20147 -430 20175
rect -402 20147 -368 20175
rect -340 20147 -306 20175
rect -278 20147 -244 20175
rect -216 20147 1625 20175
rect 1653 20147 1687 20175
rect 1715 20147 1749 20175
rect 1777 20147 1811 20175
rect 1839 20147 10625 20175
rect 10653 20147 10687 20175
rect 10715 20147 10749 20175
rect 10777 20147 10811 20175
rect 10839 20147 19625 20175
rect 19653 20147 19687 20175
rect 19715 20147 19749 20175
rect 19777 20147 19811 20175
rect 19839 20147 28625 20175
rect 28653 20147 28687 20175
rect 28715 20147 28749 20175
rect 28777 20147 28811 20175
rect 28839 20147 37625 20175
rect 37653 20147 37687 20175
rect 37715 20147 37749 20175
rect 37777 20147 37811 20175
rect 37839 20147 46625 20175
rect 46653 20147 46687 20175
rect 46715 20147 46749 20175
rect 46777 20147 46811 20175
rect 46839 20147 55625 20175
rect 55653 20147 55687 20175
rect 55715 20147 55749 20175
rect 55777 20147 55811 20175
rect 55839 20147 64625 20175
rect 64653 20147 64687 20175
rect 64715 20147 64749 20175
rect 64777 20147 64811 20175
rect 64839 20147 73625 20175
rect 73653 20147 73687 20175
rect 73715 20147 73749 20175
rect 73777 20147 73811 20175
rect 73839 20147 82625 20175
rect 82653 20147 82687 20175
rect 82715 20147 82749 20175
rect 82777 20147 82811 20175
rect 82839 20147 91625 20175
rect 91653 20147 91687 20175
rect 91715 20147 91749 20175
rect 91777 20147 91811 20175
rect 91839 20147 100625 20175
rect 100653 20147 100687 20175
rect 100715 20147 100749 20175
rect 100777 20147 100811 20175
rect 100839 20147 109625 20175
rect 109653 20147 109687 20175
rect 109715 20147 109749 20175
rect 109777 20147 109811 20175
rect 109839 20147 118625 20175
rect 118653 20147 118687 20175
rect 118715 20147 118749 20175
rect 118777 20147 118811 20175
rect 118839 20147 127625 20175
rect 127653 20147 127687 20175
rect 127715 20147 127749 20175
rect 127777 20147 127811 20175
rect 127839 20147 136625 20175
rect 136653 20147 136687 20175
rect 136715 20147 136749 20175
rect 136777 20147 136811 20175
rect 136839 20147 145625 20175
rect 145653 20147 145687 20175
rect 145715 20147 145749 20175
rect 145777 20147 145811 20175
rect 145839 20147 154625 20175
rect 154653 20147 154687 20175
rect 154715 20147 154749 20175
rect 154777 20147 154811 20175
rect 154839 20147 163625 20175
rect 163653 20147 163687 20175
rect 163715 20147 163749 20175
rect 163777 20147 163811 20175
rect 163839 20147 172625 20175
rect 172653 20147 172687 20175
rect 172715 20147 172749 20175
rect 172777 20147 172811 20175
rect 172839 20147 181625 20175
rect 181653 20147 181687 20175
rect 181715 20147 181749 20175
rect 181777 20147 181811 20175
rect 181839 20147 190625 20175
rect 190653 20147 190687 20175
rect 190715 20147 190749 20175
rect 190777 20147 190811 20175
rect 190839 20147 199625 20175
rect 199653 20147 199687 20175
rect 199715 20147 199749 20175
rect 199777 20147 199811 20175
rect 199839 20147 208625 20175
rect 208653 20147 208687 20175
rect 208715 20147 208749 20175
rect 208777 20147 208811 20175
rect 208839 20147 217625 20175
rect 217653 20147 217687 20175
rect 217715 20147 217749 20175
rect 217777 20147 217811 20175
rect 217839 20147 226625 20175
rect 226653 20147 226687 20175
rect 226715 20147 226749 20175
rect 226777 20147 226811 20175
rect 226839 20147 235625 20175
rect 235653 20147 235687 20175
rect 235715 20147 235749 20175
rect 235777 20147 235811 20175
rect 235839 20147 244625 20175
rect 244653 20147 244687 20175
rect 244715 20147 244749 20175
rect 244777 20147 244811 20175
rect 244839 20147 253625 20175
rect 253653 20147 253687 20175
rect 253715 20147 253749 20175
rect 253777 20147 253811 20175
rect 253839 20147 262625 20175
rect 262653 20147 262687 20175
rect 262715 20147 262749 20175
rect 262777 20147 262811 20175
rect 262839 20147 271625 20175
rect 271653 20147 271687 20175
rect 271715 20147 271749 20175
rect 271777 20147 271811 20175
rect 271839 20147 280625 20175
rect 280653 20147 280687 20175
rect 280715 20147 280749 20175
rect 280777 20147 280811 20175
rect 280839 20147 289625 20175
rect 289653 20147 289687 20175
rect 289715 20147 289749 20175
rect 289777 20147 289811 20175
rect 289839 20147 298248 20175
rect 298276 20147 298310 20175
rect 298338 20147 298372 20175
rect 298400 20147 298434 20175
rect 298462 20147 298990 20175
rect -958 20113 298990 20147
rect -958 20085 -430 20113
rect -402 20085 -368 20113
rect -340 20085 -306 20113
rect -278 20085 -244 20113
rect -216 20085 1625 20113
rect 1653 20085 1687 20113
rect 1715 20085 1749 20113
rect 1777 20085 1811 20113
rect 1839 20085 10625 20113
rect 10653 20085 10687 20113
rect 10715 20085 10749 20113
rect 10777 20085 10811 20113
rect 10839 20085 19625 20113
rect 19653 20085 19687 20113
rect 19715 20085 19749 20113
rect 19777 20085 19811 20113
rect 19839 20085 28625 20113
rect 28653 20085 28687 20113
rect 28715 20085 28749 20113
rect 28777 20085 28811 20113
rect 28839 20085 37625 20113
rect 37653 20085 37687 20113
rect 37715 20085 37749 20113
rect 37777 20085 37811 20113
rect 37839 20085 46625 20113
rect 46653 20085 46687 20113
rect 46715 20085 46749 20113
rect 46777 20085 46811 20113
rect 46839 20085 55625 20113
rect 55653 20085 55687 20113
rect 55715 20085 55749 20113
rect 55777 20085 55811 20113
rect 55839 20085 64625 20113
rect 64653 20085 64687 20113
rect 64715 20085 64749 20113
rect 64777 20085 64811 20113
rect 64839 20085 73625 20113
rect 73653 20085 73687 20113
rect 73715 20085 73749 20113
rect 73777 20085 73811 20113
rect 73839 20085 82625 20113
rect 82653 20085 82687 20113
rect 82715 20085 82749 20113
rect 82777 20085 82811 20113
rect 82839 20085 91625 20113
rect 91653 20085 91687 20113
rect 91715 20085 91749 20113
rect 91777 20085 91811 20113
rect 91839 20085 100625 20113
rect 100653 20085 100687 20113
rect 100715 20085 100749 20113
rect 100777 20085 100811 20113
rect 100839 20085 109625 20113
rect 109653 20085 109687 20113
rect 109715 20085 109749 20113
rect 109777 20085 109811 20113
rect 109839 20085 118625 20113
rect 118653 20085 118687 20113
rect 118715 20085 118749 20113
rect 118777 20085 118811 20113
rect 118839 20085 127625 20113
rect 127653 20085 127687 20113
rect 127715 20085 127749 20113
rect 127777 20085 127811 20113
rect 127839 20085 136625 20113
rect 136653 20085 136687 20113
rect 136715 20085 136749 20113
rect 136777 20085 136811 20113
rect 136839 20085 145625 20113
rect 145653 20085 145687 20113
rect 145715 20085 145749 20113
rect 145777 20085 145811 20113
rect 145839 20085 154625 20113
rect 154653 20085 154687 20113
rect 154715 20085 154749 20113
rect 154777 20085 154811 20113
rect 154839 20085 163625 20113
rect 163653 20085 163687 20113
rect 163715 20085 163749 20113
rect 163777 20085 163811 20113
rect 163839 20085 172625 20113
rect 172653 20085 172687 20113
rect 172715 20085 172749 20113
rect 172777 20085 172811 20113
rect 172839 20085 181625 20113
rect 181653 20085 181687 20113
rect 181715 20085 181749 20113
rect 181777 20085 181811 20113
rect 181839 20085 190625 20113
rect 190653 20085 190687 20113
rect 190715 20085 190749 20113
rect 190777 20085 190811 20113
rect 190839 20085 199625 20113
rect 199653 20085 199687 20113
rect 199715 20085 199749 20113
rect 199777 20085 199811 20113
rect 199839 20085 208625 20113
rect 208653 20085 208687 20113
rect 208715 20085 208749 20113
rect 208777 20085 208811 20113
rect 208839 20085 217625 20113
rect 217653 20085 217687 20113
rect 217715 20085 217749 20113
rect 217777 20085 217811 20113
rect 217839 20085 226625 20113
rect 226653 20085 226687 20113
rect 226715 20085 226749 20113
rect 226777 20085 226811 20113
rect 226839 20085 235625 20113
rect 235653 20085 235687 20113
rect 235715 20085 235749 20113
rect 235777 20085 235811 20113
rect 235839 20085 244625 20113
rect 244653 20085 244687 20113
rect 244715 20085 244749 20113
rect 244777 20085 244811 20113
rect 244839 20085 253625 20113
rect 253653 20085 253687 20113
rect 253715 20085 253749 20113
rect 253777 20085 253811 20113
rect 253839 20085 262625 20113
rect 262653 20085 262687 20113
rect 262715 20085 262749 20113
rect 262777 20085 262811 20113
rect 262839 20085 271625 20113
rect 271653 20085 271687 20113
rect 271715 20085 271749 20113
rect 271777 20085 271811 20113
rect 271839 20085 280625 20113
rect 280653 20085 280687 20113
rect 280715 20085 280749 20113
rect 280777 20085 280811 20113
rect 280839 20085 289625 20113
rect 289653 20085 289687 20113
rect 289715 20085 289749 20113
rect 289777 20085 289811 20113
rect 289839 20085 298248 20113
rect 298276 20085 298310 20113
rect 298338 20085 298372 20113
rect 298400 20085 298434 20113
rect 298462 20085 298990 20113
rect -958 20051 298990 20085
rect -958 20023 -430 20051
rect -402 20023 -368 20051
rect -340 20023 -306 20051
rect -278 20023 -244 20051
rect -216 20023 1625 20051
rect 1653 20023 1687 20051
rect 1715 20023 1749 20051
rect 1777 20023 1811 20051
rect 1839 20023 10625 20051
rect 10653 20023 10687 20051
rect 10715 20023 10749 20051
rect 10777 20023 10811 20051
rect 10839 20023 19625 20051
rect 19653 20023 19687 20051
rect 19715 20023 19749 20051
rect 19777 20023 19811 20051
rect 19839 20023 28625 20051
rect 28653 20023 28687 20051
rect 28715 20023 28749 20051
rect 28777 20023 28811 20051
rect 28839 20023 37625 20051
rect 37653 20023 37687 20051
rect 37715 20023 37749 20051
rect 37777 20023 37811 20051
rect 37839 20023 46625 20051
rect 46653 20023 46687 20051
rect 46715 20023 46749 20051
rect 46777 20023 46811 20051
rect 46839 20023 55625 20051
rect 55653 20023 55687 20051
rect 55715 20023 55749 20051
rect 55777 20023 55811 20051
rect 55839 20023 64625 20051
rect 64653 20023 64687 20051
rect 64715 20023 64749 20051
rect 64777 20023 64811 20051
rect 64839 20023 73625 20051
rect 73653 20023 73687 20051
rect 73715 20023 73749 20051
rect 73777 20023 73811 20051
rect 73839 20023 82625 20051
rect 82653 20023 82687 20051
rect 82715 20023 82749 20051
rect 82777 20023 82811 20051
rect 82839 20023 91625 20051
rect 91653 20023 91687 20051
rect 91715 20023 91749 20051
rect 91777 20023 91811 20051
rect 91839 20023 100625 20051
rect 100653 20023 100687 20051
rect 100715 20023 100749 20051
rect 100777 20023 100811 20051
rect 100839 20023 109625 20051
rect 109653 20023 109687 20051
rect 109715 20023 109749 20051
rect 109777 20023 109811 20051
rect 109839 20023 118625 20051
rect 118653 20023 118687 20051
rect 118715 20023 118749 20051
rect 118777 20023 118811 20051
rect 118839 20023 127625 20051
rect 127653 20023 127687 20051
rect 127715 20023 127749 20051
rect 127777 20023 127811 20051
rect 127839 20023 136625 20051
rect 136653 20023 136687 20051
rect 136715 20023 136749 20051
rect 136777 20023 136811 20051
rect 136839 20023 145625 20051
rect 145653 20023 145687 20051
rect 145715 20023 145749 20051
rect 145777 20023 145811 20051
rect 145839 20023 154625 20051
rect 154653 20023 154687 20051
rect 154715 20023 154749 20051
rect 154777 20023 154811 20051
rect 154839 20023 163625 20051
rect 163653 20023 163687 20051
rect 163715 20023 163749 20051
rect 163777 20023 163811 20051
rect 163839 20023 172625 20051
rect 172653 20023 172687 20051
rect 172715 20023 172749 20051
rect 172777 20023 172811 20051
rect 172839 20023 181625 20051
rect 181653 20023 181687 20051
rect 181715 20023 181749 20051
rect 181777 20023 181811 20051
rect 181839 20023 190625 20051
rect 190653 20023 190687 20051
rect 190715 20023 190749 20051
rect 190777 20023 190811 20051
rect 190839 20023 199625 20051
rect 199653 20023 199687 20051
rect 199715 20023 199749 20051
rect 199777 20023 199811 20051
rect 199839 20023 208625 20051
rect 208653 20023 208687 20051
rect 208715 20023 208749 20051
rect 208777 20023 208811 20051
rect 208839 20023 217625 20051
rect 217653 20023 217687 20051
rect 217715 20023 217749 20051
rect 217777 20023 217811 20051
rect 217839 20023 226625 20051
rect 226653 20023 226687 20051
rect 226715 20023 226749 20051
rect 226777 20023 226811 20051
rect 226839 20023 235625 20051
rect 235653 20023 235687 20051
rect 235715 20023 235749 20051
rect 235777 20023 235811 20051
rect 235839 20023 244625 20051
rect 244653 20023 244687 20051
rect 244715 20023 244749 20051
rect 244777 20023 244811 20051
rect 244839 20023 253625 20051
rect 253653 20023 253687 20051
rect 253715 20023 253749 20051
rect 253777 20023 253811 20051
rect 253839 20023 262625 20051
rect 262653 20023 262687 20051
rect 262715 20023 262749 20051
rect 262777 20023 262811 20051
rect 262839 20023 271625 20051
rect 271653 20023 271687 20051
rect 271715 20023 271749 20051
rect 271777 20023 271811 20051
rect 271839 20023 280625 20051
rect 280653 20023 280687 20051
rect 280715 20023 280749 20051
rect 280777 20023 280811 20051
rect 280839 20023 289625 20051
rect 289653 20023 289687 20051
rect 289715 20023 289749 20051
rect 289777 20023 289811 20051
rect 289839 20023 298248 20051
rect 298276 20023 298310 20051
rect 298338 20023 298372 20051
rect 298400 20023 298434 20051
rect 298462 20023 298990 20051
rect -958 19989 298990 20023
rect -958 19961 -430 19989
rect -402 19961 -368 19989
rect -340 19961 -306 19989
rect -278 19961 -244 19989
rect -216 19961 1625 19989
rect 1653 19961 1687 19989
rect 1715 19961 1749 19989
rect 1777 19961 1811 19989
rect 1839 19961 10625 19989
rect 10653 19961 10687 19989
rect 10715 19961 10749 19989
rect 10777 19961 10811 19989
rect 10839 19961 19625 19989
rect 19653 19961 19687 19989
rect 19715 19961 19749 19989
rect 19777 19961 19811 19989
rect 19839 19961 28625 19989
rect 28653 19961 28687 19989
rect 28715 19961 28749 19989
rect 28777 19961 28811 19989
rect 28839 19961 37625 19989
rect 37653 19961 37687 19989
rect 37715 19961 37749 19989
rect 37777 19961 37811 19989
rect 37839 19961 46625 19989
rect 46653 19961 46687 19989
rect 46715 19961 46749 19989
rect 46777 19961 46811 19989
rect 46839 19961 55625 19989
rect 55653 19961 55687 19989
rect 55715 19961 55749 19989
rect 55777 19961 55811 19989
rect 55839 19961 64625 19989
rect 64653 19961 64687 19989
rect 64715 19961 64749 19989
rect 64777 19961 64811 19989
rect 64839 19961 73625 19989
rect 73653 19961 73687 19989
rect 73715 19961 73749 19989
rect 73777 19961 73811 19989
rect 73839 19961 82625 19989
rect 82653 19961 82687 19989
rect 82715 19961 82749 19989
rect 82777 19961 82811 19989
rect 82839 19961 91625 19989
rect 91653 19961 91687 19989
rect 91715 19961 91749 19989
rect 91777 19961 91811 19989
rect 91839 19961 100625 19989
rect 100653 19961 100687 19989
rect 100715 19961 100749 19989
rect 100777 19961 100811 19989
rect 100839 19961 109625 19989
rect 109653 19961 109687 19989
rect 109715 19961 109749 19989
rect 109777 19961 109811 19989
rect 109839 19961 118625 19989
rect 118653 19961 118687 19989
rect 118715 19961 118749 19989
rect 118777 19961 118811 19989
rect 118839 19961 127625 19989
rect 127653 19961 127687 19989
rect 127715 19961 127749 19989
rect 127777 19961 127811 19989
rect 127839 19961 136625 19989
rect 136653 19961 136687 19989
rect 136715 19961 136749 19989
rect 136777 19961 136811 19989
rect 136839 19961 145625 19989
rect 145653 19961 145687 19989
rect 145715 19961 145749 19989
rect 145777 19961 145811 19989
rect 145839 19961 154625 19989
rect 154653 19961 154687 19989
rect 154715 19961 154749 19989
rect 154777 19961 154811 19989
rect 154839 19961 163625 19989
rect 163653 19961 163687 19989
rect 163715 19961 163749 19989
rect 163777 19961 163811 19989
rect 163839 19961 172625 19989
rect 172653 19961 172687 19989
rect 172715 19961 172749 19989
rect 172777 19961 172811 19989
rect 172839 19961 181625 19989
rect 181653 19961 181687 19989
rect 181715 19961 181749 19989
rect 181777 19961 181811 19989
rect 181839 19961 190625 19989
rect 190653 19961 190687 19989
rect 190715 19961 190749 19989
rect 190777 19961 190811 19989
rect 190839 19961 199625 19989
rect 199653 19961 199687 19989
rect 199715 19961 199749 19989
rect 199777 19961 199811 19989
rect 199839 19961 208625 19989
rect 208653 19961 208687 19989
rect 208715 19961 208749 19989
rect 208777 19961 208811 19989
rect 208839 19961 217625 19989
rect 217653 19961 217687 19989
rect 217715 19961 217749 19989
rect 217777 19961 217811 19989
rect 217839 19961 226625 19989
rect 226653 19961 226687 19989
rect 226715 19961 226749 19989
rect 226777 19961 226811 19989
rect 226839 19961 235625 19989
rect 235653 19961 235687 19989
rect 235715 19961 235749 19989
rect 235777 19961 235811 19989
rect 235839 19961 244625 19989
rect 244653 19961 244687 19989
rect 244715 19961 244749 19989
rect 244777 19961 244811 19989
rect 244839 19961 253625 19989
rect 253653 19961 253687 19989
rect 253715 19961 253749 19989
rect 253777 19961 253811 19989
rect 253839 19961 262625 19989
rect 262653 19961 262687 19989
rect 262715 19961 262749 19989
rect 262777 19961 262811 19989
rect 262839 19961 271625 19989
rect 271653 19961 271687 19989
rect 271715 19961 271749 19989
rect 271777 19961 271811 19989
rect 271839 19961 280625 19989
rect 280653 19961 280687 19989
rect 280715 19961 280749 19989
rect 280777 19961 280811 19989
rect 280839 19961 289625 19989
rect 289653 19961 289687 19989
rect 289715 19961 289749 19989
rect 289777 19961 289811 19989
rect 289839 19961 298248 19989
rect 298276 19961 298310 19989
rect 298338 19961 298372 19989
rect 298400 19961 298434 19989
rect 298462 19961 298990 19989
rect -958 19913 298990 19961
rect -958 14175 298990 14223
rect -958 14147 -910 14175
rect -882 14147 -848 14175
rect -820 14147 -786 14175
rect -758 14147 -724 14175
rect -696 14147 3485 14175
rect 3513 14147 3547 14175
rect 3575 14147 3609 14175
rect 3637 14147 3671 14175
rect 3699 14147 12485 14175
rect 12513 14147 12547 14175
rect 12575 14147 12609 14175
rect 12637 14147 12671 14175
rect 12699 14147 21485 14175
rect 21513 14147 21547 14175
rect 21575 14147 21609 14175
rect 21637 14147 21671 14175
rect 21699 14147 30485 14175
rect 30513 14147 30547 14175
rect 30575 14147 30609 14175
rect 30637 14147 30671 14175
rect 30699 14147 39485 14175
rect 39513 14147 39547 14175
rect 39575 14147 39609 14175
rect 39637 14147 39671 14175
rect 39699 14147 48485 14175
rect 48513 14147 48547 14175
rect 48575 14147 48609 14175
rect 48637 14147 48671 14175
rect 48699 14147 57485 14175
rect 57513 14147 57547 14175
rect 57575 14147 57609 14175
rect 57637 14147 57671 14175
rect 57699 14147 66485 14175
rect 66513 14147 66547 14175
rect 66575 14147 66609 14175
rect 66637 14147 66671 14175
rect 66699 14147 75485 14175
rect 75513 14147 75547 14175
rect 75575 14147 75609 14175
rect 75637 14147 75671 14175
rect 75699 14147 84485 14175
rect 84513 14147 84547 14175
rect 84575 14147 84609 14175
rect 84637 14147 84671 14175
rect 84699 14147 93485 14175
rect 93513 14147 93547 14175
rect 93575 14147 93609 14175
rect 93637 14147 93671 14175
rect 93699 14147 102485 14175
rect 102513 14147 102547 14175
rect 102575 14147 102609 14175
rect 102637 14147 102671 14175
rect 102699 14147 111485 14175
rect 111513 14147 111547 14175
rect 111575 14147 111609 14175
rect 111637 14147 111671 14175
rect 111699 14147 120485 14175
rect 120513 14147 120547 14175
rect 120575 14147 120609 14175
rect 120637 14147 120671 14175
rect 120699 14147 129485 14175
rect 129513 14147 129547 14175
rect 129575 14147 129609 14175
rect 129637 14147 129671 14175
rect 129699 14147 138485 14175
rect 138513 14147 138547 14175
rect 138575 14147 138609 14175
rect 138637 14147 138671 14175
rect 138699 14147 147485 14175
rect 147513 14147 147547 14175
rect 147575 14147 147609 14175
rect 147637 14147 147671 14175
rect 147699 14147 156485 14175
rect 156513 14147 156547 14175
rect 156575 14147 156609 14175
rect 156637 14147 156671 14175
rect 156699 14147 165485 14175
rect 165513 14147 165547 14175
rect 165575 14147 165609 14175
rect 165637 14147 165671 14175
rect 165699 14147 174485 14175
rect 174513 14147 174547 14175
rect 174575 14147 174609 14175
rect 174637 14147 174671 14175
rect 174699 14147 183485 14175
rect 183513 14147 183547 14175
rect 183575 14147 183609 14175
rect 183637 14147 183671 14175
rect 183699 14147 192485 14175
rect 192513 14147 192547 14175
rect 192575 14147 192609 14175
rect 192637 14147 192671 14175
rect 192699 14147 201485 14175
rect 201513 14147 201547 14175
rect 201575 14147 201609 14175
rect 201637 14147 201671 14175
rect 201699 14147 210485 14175
rect 210513 14147 210547 14175
rect 210575 14147 210609 14175
rect 210637 14147 210671 14175
rect 210699 14147 219485 14175
rect 219513 14147 219547 14175
rect 219575 14147 219609 14175
rect 219637 14147 219671 14175
rect 219699 14147 228485 14175
rect 228513 14147 228547 14175
rect 228575 14147 228609 14175
rect 228637 14147 228671 14175
rect 228699 14147 237485 14175
rect 237513 14147 237547 14175
rect 237575 14147 237609 14175
rect 237637 14147 237671 14175
rect 237699 14147 246485 14175
rect 246513 14147 246547 14175
rect 246575 14147 246609 14175
rect 246637 14147 246671 14175
rect 246699 14147 255485 14175
rect 255513 14147 255547 14175
rect 255575 14147 255609 14175
rect 255637 14147 255671 14175
rect 255699 14147 264485 14175
rect 264513 14147 264547 14175
rect 264575 14147 264609 14175
rect 264637 14147 264671 14175
rect 264699 14147 273485 14175
rect 273513 14147 273547 14175
rect 273575 14147 273609 14175
rect 273637 14147 273671 14175
rect 273699 14147 282485 14175
rect 282513 14147 282547 14175
rect 282575 14147 282609 14175
rect 282637 14147 282671 14175
rect 282699 14147 291485 14175
rect 291513 14147 291547 14175
rect 291575 14147 291609 14175
rect 291637 14147 291671 14175
rect 291699 14147 298728 14175
rect 298756 14147 298790 14175
rect 298818 14147 298852 14175
rect 298880 14147 298914 14175
rect 298942 14147 298990 14175
rect -958 14113 298990 14147
rect -958 14085 -910 14113
rect -882 14085 -848 14113
rect -820 14085 -786 14113
rect -758 14085 -724 14113
rect -696 14085 3485 14113
rect 3513 14085 3547 14113
rect 3575 14085 3609 14113
rect 3637 14085 3671 14113
rect 3699 14085 12485 14113
rect 12513 14085 12547 14113
rect 12575 14085 12609 14113
rect 12637 14085 12671 14113
rect 12699 14085 21485 14113
rect 21513 14085 21547 14113
rect 21575 14085 21609 14113
rect 21637 14085 21671 14113
rect 21699 14085 30485 14113
rect 30513 14085 30547 14113
rect 30575 14085 30609 14113
rect 30637 14085 30671 14113
rect 30699 14085 39485 14113
rect 39513 14085 39547 14113
rect 39575 14085 39609 14113
rect 39637 14085 39671 14113
rect 39699 14085 48485 14113
rect 48513 14085 48547 14113
rect 48575 14085 48609 14113
rect 48637 14085 48671 14113
rect 48699 14085 57485 14113
rect 57513 14085 57547 14113
rect 57575 14085 57609 14113
rect 57637 14085 57671 14113
rect 57699 14085 66485 14113
rect 66513 14085 66547 14113
rect 66575 14085 66609 14113
rect 66637 14085 66671 14113
rect 66699 14085 75485 14113
rect 75513 14085 75547 14113
rect 75575 14085 75609 14113
rect 75637 14085 75671 14113
rect 75699 14085 84485 14113
rect 84513 14085 84547 14113
rect 84575 14085 84609 14113
rect 84637 14085 84671 14113
rect 84699 14085 93485 14113
rect 93513 14085 93547 14113
rect 93575 14085 93609 14113
rect 93637 14085 93671 14113
rect 93699 14085 102485 14113
rect 102513 14085 102547 14113
rect 102575 14085 102609 14113
rect 102637 14085 102671 14113
rect 102699 14085 111485 14113
rect 111513 14085 111547 14113
rect 111575 14085 111609 14113
rect 111637 14085 111671 14113
rect 111699 14085 120485 14113
rect 120513 14085 120547 14113
rect 120575 14085 120609 14113
rect 120637 14085 120671 14113
rect 120699 14085 129485 14113
rect 129513 14085 129547 14113
rect 129575 14085 129609 14113
rect 129637 14085 129671 14113
rect 129699 14085 138485 14113
rect 138513 14085 138547 14113
rect 138575 14085 138609 14113
rect 138637 14085 138671 14113
rect 138699 14085 147485 14113
rect 147513 14085 147547 14113
rect 147575 14085 147609 14113
rect 147637 14085 147671 14113
rect 147699 14085 156485 14113
rect 156513 14085 156547 14113
rect 156575 14085 156609 14113
rect 156637 14085 156671 14113
rect 156699 14085 165485 14113
rect 165513 14085 165547 14113
rect 165575 14085 165609 14113
rect 165637 14085 165671 14113
rect 165699 14085 174485 14113
rect 174513 14085 174547 14113
rect 174575 14085 174609 14113
rect 174637 14085 174671 14113
rect 174699 14085 183485 14113
rect 183513 14085 183547 14113
rect 183575 14085 183609 14113
rect 183637 14085 183671 14113
rect 183699 14085 192485 14113
rect 192513 14085 192547 14113
rect 192575 14085 192609 14113
rect 192637 14085 192671 14113
rect 192699 14085 201485 14113
rect 201513 14085 201547 14113
rect 201575 14085 201609 14113
rect 201637 14085 201671 14113
rect 201699 14085 210485 14113
rect 210513 14085 210547 14113
rect 210575 14085 210609 14113
rect 210637 14085 210671 14113
rect 210699 14085 219485 14113
rect 219513 14085 219547 14113
rect 219575 14085 219609 14113
rect 219637 14085 219671 14113
rect 219699 14085 228485 14113
rect 228513 14085 228547 14113
rect 228575 14085 228609 14113
rect 228637 14085 228671 14113
rect 228699 14085 237485 14113
rect 237513 14085 237547 14113
rect 237575 14085 237609 14113
rect 237637 14085 237671 14113
rect 237699 14085 246485 14113
rect 246513 14085 246547 14113
rect 246575 14085 246609 14113
rect 246637 14085 246671 14113
rect 246699 14085 255485 14113
rect 255513 14085 255547 14113
rect 255575 14085 255609 14113
rect 255637 14085 255671 14113
rect 255699 14085 264485 14113
rect 264513 14085 264547 14113
rect 264575 14085 264609 14113
rect 264637 14085 264671 14113
rect 264699 14085 273485 14113
rect 273513 14085 273547 14113
rect 273575 14085 273609 14113
rect 273637 14085 273671 14113
rect 273699 14085 282485 14113
rect 282513 14085 282547 14113
rect 282575 14085 282609 14113
rect 282637 14085 282671 14113
rect 282699 14085 291485 14113
rect 291513 14085 291547 14113
rect 291575 14085 291609 14113
rect 291637 14085 291671 14113
rect 291699 14085 298728 14113
rect 298756 14085 298790 14113
rect 298818 14085 298852 14113
rect 298880 14085 298914 14113
rect 298942 14085 298990 14113
rect -958 14051 298990 14085
rect -958 14023 -910 14051
rect -882 14023 -848 14051
rect -820 14023 -786 14051
rect -758 14023 -724 14051
rect -696 14023 3485 14051
rect 3513 14023 3547 14051
rect 3575 14023 3609 14051
rect 3637 14023 3671 14051
rect 3699 14023 12485 14051
rect 12513 14023 12547 14051
rect 12575 14023 12609 14051
rect 12637 14023 12671 14051
rect 12699 14023 21485 14051
rect 21513 14023 21547 14051
rect 21575 14023 21609 14051
rect 21637 14023 21671 14051
rect 21699 14023 30485 14051
rect 30513 14023 30547 14051
rect 30575 14023 30609 14051
rect 30637 14023 30671 14051
rect 30699 14023 39485 14051
rect 39513 14023 39547 14051
rect 39575 14023 39609 14051
rect 39637 14023 39671 14051
rect 39699 14023 48485 14051
rect 48513 14023 48547 14051
rect 48575 14023 48609 14051
rect 48637 14023 48671 14051
rect 48699 14023 57485 14051
rect 57513 14023 57547 14051
rect 57575 14023 57609 14051
rect 57637 14023 57671 14051
rect 57699 14023 66485 14051
rect 66513 14023 66547 14051
rect 66575 14023 66609 14051
rect 66637 14023 66671 14051
rect 66699 14023 75485 14051
rect 75513 14023 75547 14051
rect 75575 14023 75609 14051
rect 75637 14023 75671 14051
rect 75699 14023 84485 14051
rect 84513 14023 84547 14051
rect 84575 14023 84609 14051
rect 84637 14023 84671 14051
rect 84699 14023 93485 14051
rect 93513 14023 93547 14051
rect 93575 14023 93609 14051
rect 93637 14023 93671 14051
rect 93699 14023 102485 14051
rect 102513 14023 102547 14051
rect 102575 14023 102609 14051
rect 102637 14023 102671 14051
rect 102699 14023 111485 14051
rect 111513 14023 111547 14051
rect 111575 14023 111609 14051
rect 111637 14023 111671 14051
rect 111699 14023 120485 14051
rect 120513 14023 120547 14051
rect 120575 14023 120609 14051
rect 120637 14023 120671 14051
rect 120699 14023 129485 14051
rect 129513 14023 129547 14051
rect 129575 14023 129609 14051
rect 129637 14023 129671 14051
rect 129699 14023 138485 14051
rect 138513 14023 138547 14051
rect 138575 14023 138609 14051
rect 138637 14023 138671 14051
rect 138699 14023 147485 14051
rect 147513 14023 147547 14051
rect 147575 14023 147609 14051
rect 147637 14023 147671 14051
rect 147699 14023 156485 14051
rect 156513 14023 156547 14051
rect 156575 14023 156609 14051
rect 156637 14023 156671 14051
rect 156699 14023 165485 14051
rect 165513 14023 165547 14051
rect 165575 14023 165609 14051
rect 165637 14023 165671 14051
rect 165699 14023 174485 14051
rect 174513 14023 174547 14051
rect 174575 14023 174609 14051
rect 174637 14023 174671 14051
rect 174699 14023 183485 14051
rect 183513 14023 183547 14051
rect 183575 14023 183609 14051
rect 183637 14023 183671 14051
rect 183699 14023 192485 14051
rect 192513 14023 192547 14051
rect 192575 14023 192609 14051
rect 192637 14023 192671 14051
rect 192699 14023 201485 14051
rect 201513 14023 201547 14051
rect 201575 14023 201609 14051
rect 201637 14023 201671 14051
rect 201699 14023 210485 14051
rect 210513 14023 210547 14051
rect 210575 14023 210609 14051
rect 210637 14023 210671 14051
rect 210699 14023 219485 14051
rect 219513 14023 219547 14051
rect 219575 14023 219609 14051
rect 219637 14023 219671 14051
rect 219699 14023 228485 14051
rect 228513 14023 228547 14051
rect 228575 14023 228609 14051
rect 228637 14023 228671 14051
rect 228699 14023 237485 14051
rect 237513 14023 237547 14051
rect 237575 14023 237609 14051
rect 237637 14023 237671 14051
rect 237699 14023 246485 14051
rect 246513 14023 246547 14051
rect 246575 14023 246609 14051
rect 246637 14023 246671 14051
rect 246699 14023 255485 14051
rect 255513 14023 255547 14051
rect 255575 14023 255609 14051
rect 255637 14023 255671 14051
rect 255699 14023 264485 14051
rect 264513 14023 264547 14051
rect 264575 14023 264609 14051
rect 264637 14023 264671 14051
rect 264699 14023 273485 14051
rect 273513 14023 273547 14051
rect 273575 14023 273609 14051
rect 273637 14023 273671 14051
rect 273699 14023 282485 14051
rect 282513 14023 282547 14051
rect 282575 14023 282609 14051
rect 282637 14023 282671 14051
rect 282699 14023 291485 14051
rect 291513 14023 291547 14051
rect 291575 14023 291609 14051
rect 291637 14023 291671 14051
rect 291699 14023 298728 14051
rect 298756 14023 298790 14051
rect 298818 14023 298852 14051
rect 298880 14023 298914 14051
rect 298942 14023 298990 14051
rect -958 13989 298990 14023
rect -958 13961 -910 13989
rect -882 13961 -848 13989
rect -820 13961 -786 13989
rect -758 13961 -724 13989
rect -696 13961 3485 13989
rect 3513 13961 3547 13989
rect 3575 13961 3609 13989
rect 3637 13961 3671 13989
rect 3699 13961 12485 13989
rect 12513 13961 12547 13989
rect 12575 13961 12609 13989
rect 12637 13961 12671 13989
rect 12699 13961 21485 13989
rect 21513 13961 21547 13989
rect 21575 13961 21609 13989
rect 21637 13961 21671 13989
rect 21699 13961 30485 13989
rect 30513 13961 30547 13989
rect 30575 13961 30609 13989
rect 30637 13961 30671 13989
rect 30699 13961 39485 13989
rect 39513 13961 39547 13989
rect 39575 13961 39609 13989
rect 39637 13961 39671 13989
rect 39699 13961 48485 13989
rect 48513 13961 48547 13989
rect 48575 13961 48609 13989
rect 48637 13961 48671 13989
rect 48699 13961 57485 13989
rect 57513 13961 57547 13989
rect 57575 13961 57609 13989
rect 57637 13961 57671 13989
rect 57699 13961 66485 13989
rect 66513 13961 66547 13989
rect 66575 13961 66609 13989
rect 66637 13961 66671 13989
rect 66699 13961 75485 13989
rect 75513 13961 75547 13989
rect 75575 13961 75609 13989
rect 75637 13961 75671 13989
rect 75699 13961 84485 13989
rect 84513 13961 84547 13989
rect 84575 13961 84609 13989
rect 84637 13961 84671 13989
rect 84699 13961 93485 13989
rect 93513 13961 93547 13989
rect 93575 13961 93609 13989
rect 93637 13961 93671 13989
rect 93699 13961 102485 13989
rect 102513 13961 102547 13989
rect 102575 13961 102609 13989
rect 102637 13961 102671 13989
rect 102699 13961 111485 13989
rect 111513 13961 111547 13989
rect 111575 13961 111609 13989
rect 111637 13961 111671 13989
rect 111699 13961 120485 13989
rect 120513 13961 120547 13989
rect 120575 13961 120609 13989
rect 120637 13961 120671 13989
rect 120699 13961 129485 13989
rect 129513 13961 129547 13989
rect 129575 13961 129609 13989
rect 129637 13961 129671 13989
rect 129699 13961 138485 13989
rect 138513 13961 138547 13989
rect 138575 13961 138609 13989
rect 138637 13961 138671 13989
rect 138699 13961 147485 13989
rect 147513 13961 147547 13989
rect 147575 13961 147609 13989
rect 147637 13961 147671 13989
rect 147699 13961 156485 13989
rect 156513 13961 156547 13989
rect 156575 13961 156609 13989
rect 156637 13961 156671 13989
rect 156699 13961 165485 13989
rect 165513 13961 165547 13989
rect 165575 13961 165609 13989
rect 165637 13961 165671 13989
rect 165699 13961 174485 13989
rect 174513 13961 174547 13989
rect 174575 13961 174609 13989
rect 174637 13961 174671 13989
rect 174699 13961 183485 13989
rect 183513 13961 183547 13989
rect 183575 13961 183609 13989
rect 183637 13961 183671 13989
rect 183699 13961 192485 13989
rect 192513 13961 192547 13989
rect 192575 13961 192609 13989
rect 192637 13961 192671 13989
rect 192699 13961 201485 13989
rect 201513 13961 201547 13989
rect 201575 13961 201609 13989
rect 201637 13961 201671 13989
rect 201699 13961 210485 13989
rect 210513 13961 210547 13989
rect 210575 13961 210609 13989
rect 210637 13961 210671 13989
rect 210699 13961 219485 13989
rect 219513 13961 219547 13989
rect 219575 13961 219609 13989
rect 219637 13961 219671 13989
rect 219699 13961 228485 13989
rect 228513 13961 228547 13989
rect 228575 13961 228609 13989
rect 228637 13961 228671 13989
rect 228699 13961 237485 13989
rect 237513 13961 237547 13989
rect 237575 13961 237609 13989
rect 237637 13961 237671 13989
rect 237699 13961 246485 13989
rect 246513 13961 246547 13989
rect 246575 13961 246609 13989
rect 246637 13961 246671 13989
rect 246699 13961 255485 13989
rect 255513 13961 255547 13989
rect 255575 13961 255609 13989
rect 255637 13961 255671 13989
rect 255699 13961 264485 13989
rect 264513 13961 264547 13989
rect 264575 13961 264609 13989
rect 264637 13961 264671 13989
rect 264699 13961 273485 13989
rect 273513 13961 273547 13989
rect 273575 13961 273609 13989
rect 273637 13961 273671 13989
rect 273699 13961 282485 13989
rect 282513 13961 282547 13989
rect 282575 13961 282609 13989
rect 282637 13961 282671 13989
rect 282699 13961 291485 13989
rect 291513 13961 291547 13989
rect 291575 13961 291609 13989
rect 291637 13961 291671 13989
rect 291699 13961 298728 13989
rect 298756 13961 298790 13989
rect 298818 13961 298852 13989
rect 298880 13961 298914 13989
rect 298942 13961 298990 13989
rect -958 13913 298990 13961
rect -958 11175 298990 11223
rect -958 11147 -430 11175
rect -402 11147 -368 11175
rect -340 11147 -306 11175
rect -278 11147 -244 11175
rect -216 11147 1625 11175
rect 1653 11147 1687 11175
rect 1715 11147 1749 11175
rect 1777 11147 1811 11175
rect 1839 11147 10625 11175
rect 10653 11147 10687 11175
rect 10715 11147 10749 11175
rect 10777 11147 10811 11175
rect 10839 11147 19625 11175
rect 19653 11147 19687 11175
rect 19715 11147 19749 11175
rect 19777 11147 19811 11175
rect 19839 11147 28625 11175
rect 28653 11147 28687 11175
rect 28715 11147 28749 11175
rect 28777 11147 28811 11175
rect 28839 11147 37625 11175
rect 37653 11147 37687 11175
rect 37715 11147 37749 11175
rect 37777 11147 37811 11175
rect 37839 11147 46625 11175
rect 46653 11147 46687 11175
rect 46715 11147 46749 11175
rect 46777 11147 46811 11175
rect 46839 11147 55625 11175
rect 55653 11147 55687 11175
rect 55715 11147 55749 11175
rect 55777 11147 55811 11175
rect 55839 11147 64625 11175
rect 64653 11147 64687 11175
rect 64715 11147 64749 11175
rect 64777 11147 64811 11175
rect 64839 11147 73625 11175
rect 73653 11147 73687 11175
rect 73715 11147 73749 11175
rect 73777 11147 73811 11175
rect 73839 11147 82625 11175
rect 82653 11147 82687 11175
rect 82715 11147 82749 11175
rect 82777 11147 82811 11175
rect 82839 11147 91625 11175
rect 91653 11147 91687 11175
rect 91715 11147 91749 11175
rect 91777 11147 91811 11175
rect 91839 11147 100625 11175
rect 100653 11147 100687 11175
rect 100715 11147 100749 11175
rect 100777 11147 100811 11175
rect 100839 11147 109625 11175
rect 109653 11147 109687 11175
rect 109715 11147 109749 11175
rect 109777 11147 109811 11175
rect 109839 11147 118625 11175
rect 118653 11147 118687 11175
rect 118715 11147 118749 11175
rect 118777 11147 118811 11175
rect 118839 11147 127625 11175
rect 127653 11147 127687 11175
rect 127715 11147 127749 11175
rect 127777 11147 127811 11175
rect 127839 11147 136625 11175
rect 136653 11147 136687 11175
rect 136715 11147 136749 11175
rect 136777 11147 136811 11175
rect 136839 11147 145625 11175
rect 145653 11147 145687 11175
rect 145715 11147 145749 11175
rect 145777 11147 145811 11175
rect 145839 11147 154625 11175
rect 154653 11147 154687 11175
rect 154715 11147 154749 11175
rect 154777 11147 154811 11175
rect 154839 11147 163625 11175
rect 163653 11147 163687 11175
rect 163715 11147 163749 11175
rect 163777 11147 163811 11175
rect 163839 11147 172625 11175
rect 172653 11147 172687 11175
rect 172715 11147 172749 11175
rect 172777 11147 172811 11175
rect 172839 11147 181625 11175
rect 181653 11147 181687 11175
rect 181715 11147 181749 11175
rect 181777 11147 181811 11175
rect 181839 11147 190625 11175
rect 190653 11147 190687 11175
rect 190715 11147 190749 11175
rect 190777 11147 190811 11175
rect 190839 11147 199625 11175
rect 199653 11147 199687 11175
rect 199715 11147 199749 11175
rect 199777 11147 199811 11175
rect 199839 11147 208625 11175
rect 208653 11147 208687 11175
rect 208715 11147 208749 11175
rect 208777 11147 208811 11175
rect 208839 11147 217625 11175
rect 217653 11147 217687 11175
rect 217715 11147 217749 11175
rect 217777 11147 217811 11175
rect 217839 11147 226625 11175
rect 226653 11147 226687 11175
rect 226715 11147 226749 11175
rect 226777 11147 226811 11175
rect 226839 11147 235625 11175
rect 235653 11147 235687 11175
rect 235715 11147 235749 11175
rect 235777 11147 235811 11175
rect 235839 11147 244625 11175
rect 244653 11147 244687 11175
rect 244715 11147 244749 11175
rect 244777 11147 244811 11175
rect 244839 11147 253625 11175
rect 253653 11147 253687 11175
rect 253715 11147 253749 11175
rect 253777 11147 253811 11175
rect 253839 11147 262625 11175
rect 262653 11147 262687 11175
rect 262715 11147 262749 11175
rect 262777 11147 262811 11175
rect 262839 11147 271625 11175
rect 271653 11147 271687 11175
rect 271715 11147 271749 11175
rect 271777 11147 271811 11175
rect 271839 11147 280625 11175
rect 280653 11147 280687 11175
rect 280715 11147 280749 11175
rect 280777 11147 280811 11175
rect 280839 11147 289625 11175
rect 289653 11147 289687 11175
rect 289715 11147 289749 11175
rect 289777 11147 289811 11175
rect 289839 11147 298248 11175
rect 298276 11147 298310 11175
rect 298338 11147 298372 11175
rect 298400 11147 298434 11175
rect 298462 11147 298990 11175
rect -958 11113 298990 11147
rect -958 11085 -430 11113
rect -402 11085 -368 11113
rect -340 11085 -306 11113
rect -278 11085 -244 11113
rect -216 11085 1625 11113
rect 1653 11085 1687 11113
rect 1715 11085 1749 11113
rect 1777 11085 1811 11113
rect 1839 11085 10625 11113
rect 10653 11085 10687 11113
rect 10715 11085 10749 11113
rect 10777 11085 10811 11113
rect 10839 11085 19625 11113
rect 19653 11085 19687 11113
rect 19715 11085 19749 11113
rect 19777 11085 19811 11113
rect 19839 11085 28625 11113
rect 28653 11085 28687 11113
rect 28715 11085 28749 11113
rect 28777 11085 28811 11113
rect 28839 11085 37625 11113
rect 37653 11085 37687 11113
rect 37715 11085 37749 11113
rect 37777 11085 37811 11113
rect 37839 11085 46625 11113
rect 46653 11085 46687 11113
rect 46715 11085 46749 11113
rect 46777 11085 46811 11113
rect 46839 11085 55625 11113
rect 55653 11085 55687 11113
rect 55715 11085 55749 11113
rect 55777 11085 55811 11113
rect 55839 11085 64625 11113
rect 64653 11085 64687 11113
rect 64715 11085 64749 11113
rect 64777 11085 64811 11113
rect 64839 11085 73625 11113
rect 73653 11085 73687 11113
rect 73715 11085 73749 11113
rect 73777 11085 73811 11113
rect 73839 11085 82625 11113
rect 82653 11085 82687 11113
rect 82715 11085 82749 11113
rect 82777 11085 82811 11113
rect 82839 11085 91625 11113
rect 91653 11085 91687 11113
rect 91715 11085 91749 11113
rect 91777 11085 91811 11113
rect 91839 11085 100625 11113
rect 100653 11085 100687 11113
rect 100715 11085 100749 11113
rect 100777 11085 100811 11113
rect 100839 11085 109625 11113
rect 109653 11085 109687 11113
rect 109715 11085 109749 11113
rect 109777 11085 109811 11113
rect 109839 11085 118625 11113
rect 118653 11085 118687 11113
rect 118715 11085 118749 11113
rect 118777 11085 118811 11113
rect 118839 11085 127625 11113
rect 127653 11085 127687 11113
rect 127715 11085 127749 11113
rect 127777 11085 127811 11113
rect 127839 11085 136625 11113
rect 136653 11085 136687 11113
rect 136715 11085 136749 11113
rect 136777 11085 136811 11113
rect 136839 11085 145625 11113
rect 145653 11085 145687 11113
rect 145715 11085 145749 11113
rect 145777 11085 145811 11113
rect 145839 11085 154625 11113
rect 154653 11085 154687 11113
rect 154715 11085 154749 11113
rect 154777 11085 154811 11113
rect 154839 11085 163625 11113
rect 163653 11085 163687 11113
rect 163715 11085 163749 11113
rect 163777 11085 163811 11113
rect 163839 11085 172625 11113
rect 172653 11085 172687 11113
rect 172715 11085 172749 11113
rect 172777 11085 172811 11113
rect 172839 11085 181625 11113
rect 181653 11085 181687 11113
rect 181715 11085 181749 11113
rect 181777 11085 181811 11113
rect 181839 11085 190625 11113
rect 190653 11085 190687 11113
rect 190715 11085 190749 11113
rect 190777 11085 190811 11113
rect 190839 11085 199625 11113
rect 199653 11085 199687 11113
rect 199715 11085 199749 11113
rect 199777 11085 199811 11113
rect 199839 11085 208625 11113
rect 208653 11085 208687 11113
rect 208715 11085 208749 11113
rect 208777 11085 208811 11113
rect 208839 11085 217625 11113
rect 217653 11085 217687 11113
rect 217715 11085 217749 11113
rect 217777 11085 217811 11113
rect 217839 11085 226625 11113
rect 226653 11085 226687 11113
rect 226715 11085 226749 11113
rect 226777 11085 226811 11113
rect 226839 11085 235625 11113
rect 235653 11085 235687 11113
rect 235715 11085 235749 11113
rect 235777 11085 235811 11113
rect 235839 11085 244625 11113
rect 244653 11085 244687 11113
rect 244715 11085 244749 11113
rect 244777 11085 244811 11113
rect 244839 11085 253625 11113
rect 253653 11085 253687 11113
rect 253715 11085 253749 11113
rect 253777 11085 253811 11113
rect 253839 11085 262625 11113
rect 262653 11085 262687 11113
rect 262715 11085 262749 11113
rect 262777 11085 262811 11113
rect 262839 11085 271625 11113
rect 271653 11085 271687 11113
rect 271715 11085 271749 11113
rect 271777 11085 271811 11113
rect 271839 11085 280625 11113
rect 280653 11085 280687 11113
rect 280715 11085 280749 11113
rect 280777 11085 280811 11113
rect 280839 11085 289625 11113
rect 289653 11085 289687 11113
rect 289715 11085 289749 11113
rect 289777 11085 289811 11113
rect 289839 11085 298248 11113
rect 298276 11085 298310 11113
rect 298338 11085 298372 11113
rect 298400 11085 298434 11113
rect 298462 11085 298990 11113
rect -958 11051 298990 11085
rect -958 11023 -430 11051
rect -402 11023 -368 11051
rect -340 11023 -306 11051
rect -278 11023 -244 11051
rect -216 11023 1625 11051
rect 1653 11023 1687 11051
rect 1715 11023 1749 11051
rect 1777 11023 1811 11051
rect 1839 11023 10625 11051
rect 10653 11023 10687 11051
rect 10715 11023 10749 11051
rect 10777 11023 10811 11051
rect 10839 11023 19625 11051
rect 19653 11023 19687 11051
rect 19715 11023 19749 11051
rect 19777 11023 19811 11051
rect 19839 11023 28625 11051
rect 28653 11023 28687 11051
rect 28715 11023 28749 11051
rect 28777 11023 28811 11051
rect 28839 11023 37625 11051
rect 37653 11023 37687 11051
rect 37715 11023 37749 11051
rect 37777 11023 37811 11051
rect 37839 11023 46625 11051
rect 46653 11023 46687 11051
rect 46715 11023 46749 11051
rect 46777 11023 46811 11051
rect 46839 11023 55625 11051
rect 55653 11023 55687 11051
rect 55715 11023 55749 11051
rect 55777 11023 55811 11051
rect 55839 11023 64625 11051
rect 64653 11023 64687 11051
rect 64715 11023 64749 11051
rect 64777 11023 64811 11051
rect 64839 11023 73625 11051
rect 73653 11023 73687 11051
rect 73715 11023 73749 11051
rect 73777 11023 73811 11051
rect 73839 11023 82625 11051
rect 82653 11023 82687 11051
rect 82715 11023 82749 11051
rect 82777 11023 82811 11051
rect 82839 11023 91625 11051
rect 91653 11023 91687 11051
rect 91715 11023 91749 11051
rect 91777 11023 91811 11051
rect 91839 11023 100625 11051
rect 100653 11023 100687 11051
rect 100715 11023 100749 11051
rect 100777 11023 100811 11051
rect 100839 11023 109625 11051
rect 109653 11023 109687 11051
rect 109715 11023 109749 11051
rect 109777 11023 109811 11051
rect 109839 11023 118625 11051
rect 118653 11023 118687 11051
rect 118715 11023 118749 11051
rect 118777 11023 118811 11051
rect 118839 11023 127625 11051
rect 127653 11023 127687 11051
rect 127715 11023 127749 11051
rect 127777 11023 127811 11051
rect 127839 11023 136625 11051
rect 136653 11023 136687 11051
rect 136715 11023 136749 11051
rect 136777 11023 136811 11051
rect 136839 11023 145625 11051
rect 145653 11023 145687 11051
rect 145715 11023 145749 11051
rect 145777 11023 145811 11051
rect 145839 11023 154625 11051
rect 154653 11023 154687 11051
rect 154715 11023 154749 11051
rect 154777 11023 154811 11051
rect 154839 11023 163625 11051
rect 163653 11023 163687 11051
rect 163715 11023 163749 11051
rect 163777 11023 163811 11051
rect 163839 11023 172625 11051
rect 172653 11023 172687 11051
rect 172715 11023 172749 11051
rect 172777 11023 172811 11051
rect 172839 11023 181625 11051
rect 181653 11023 181687 11051
rect 181715 11023 181749 11051
rect 181777 11023 181811 11051
rect 181839 11023 190625 11051
rect 190653 11023 190687 11051
rect 190715 11023 190749 11051
rect 190777 11023 190811 11051
rect 190839 11023 199625 11051
rect 199653 11023 199687 11051
rect 199715 11023 199749 11051
rect 199777 11023 199811 11051
rect 199839 11023 208625 11051
rect 208653 11023 208687 11051
rect 208715 11023 208749 11051
rect 208777 11023 208811 11051
rect 208839 11023 217625 11051
rect 217653 11023 217687 11051
rect 217715 11023 217749 11051
rect 217777 11023 217811 11051
rect 217839 11023 226625 11051
rect 226653 11023 226687 11051
rect 226715 11023 226749 11051
rect 226777 11023 226811 11051
rect 226839 11023 235625 11051
rect 235653 11023 235687 11051
rect 235715 11023 235749 11051
rect 235777 11023 235811 11051
rect 235839 11023 244625 11051
rect 244653 11023 244687 11051
rect 244715 11023 244749 11051
rect 244777 11023 244811 11051
rect 244839 11023 253625 11051
rect 253653 11023 253687 11051
rect 253715 11023 253749 11051
rect 253777 11023 253811 11051
rect 253839 11023 262625 11051
rect 262653 11023 262687 11051
rect 262715 11023 262749 11051
rect 262777 11023 262811 11051
rect 262839 11023 271625 11051
rect 271653 11023 271687 11051
rect 271715 11023 271749 11051
rect 271777 11023 271811 11051
rect 271839 11023 280625 11051
rect 280653 11023 280687 11051
rect 280715 11023 280749 11051
rect 280777 11023 280811 11051
rect 280839 11023 289625 11051
rect 289653 11023 289687 11051
rect 289715 11023 289749 11051
rect 289777 11023 289811 11051
rect 289839 11023 298248 11051
rect 298276 11023 298310 11051
rect 298338 11023 298372 11051
rect 298400 11023 298434 11051
rect 298462 11023 298990 11051
rect -958 10989 298990 11023
rect -958 10961 -430 10989
rect -402 10961 -368 10989
rect -340 10961 -306 10989
rect -278 10961 -244 10989
rect -216 10961 1625 10989
rect 1653 10961 1687 10989
rect 1715 10961 1749 10989
rect 1777 10961 1811 10989
rect 1839 10961 10625 10989
rect 10653 10961 10687 10989
rect 10715 10961 10749 10989
rect 10777 10961 10811 10989
rect 10839 10961 19625 10989
rect 19653 10961 19687 10989
rect 19715 10961 19749 10989
rect 19777 10961 19811 10989
rect 19839 10961 28625 10989
rect 28653 10961 28687 10989
rect 28715 10961 28749 10989
rect 28777 10961 28811 10989
rect 28839 10961 37625 10989
rect 37653 10961 37687 10989
rect 37715 10961 37749 10989
rect 37777 10961 37811 10989
rect 37839 10961 46625 10989
rect 46653 10961 46687 10989
rect 46715 10961 46749 10989
rect 46777 10961 46811 10989
rect 46839 10961 55625 10989
rect 55653 10961 55687 10989
rect 55715 10961 55749 10989
rect 55777 10961 55811 10989
rect 55839 10961 64625 10989
rect 64653 10961 64687 10989
rect 64715 10961 64749 10989
rect 64777 10961 64811 10989
rect 64839 10961 73625 10989
rect 73653 10961 73687 10989
rect 73715 10961 73749 10989
rect 73777 10961 73811 10989
rect 73839 10961 82625 10989
rect 82653 10961 82687 10989
rect 82715 10961 82749 10989
rect 82777 10961 82811 10989
rect 82839 10961 91625 10989
rect 91653 10961 91687 10989
rect 91715 10961 91749 10989
rect 91777 10961 91811 10989
rect 91839 10961 100625 10989
rect 100653 10961 100687 10989
rect 100715 10961 100749 10989
rect 100777 10961 100811 10989
rect 100839 10961 109625 10989
rect 109653 10961 109687 10989
rect 109715 10961 109749 10989
rect 109777 10961 109811 10989
rect 109839 10961 118625 10989
rect 118653 10961 118687 10989
rect 118715 10961 118749 10989
rect 118777 10961 118811 10989
rect 118839 10961 127625 10989
rect 127653 10961 127687 10989
rect 127715 10961 127749 10989
rect 127777 10961 127811 10989
rect 127839 10961 136625 10989
rect 136653 10961 136687 10989
rect 136715 10961 136749 10989
rect 136777 10961 136811 10989
rect 136839 10961 145625 10989
rect 145653 10961 145687 10989
rect 145715 10961 145749 10989
rect 145777 10961 145811 10989
rect 145839 10961 154625 10989
rect 154653 10961 154687 10989
rect 154715 10961 154749 10989
rect 154777 10961 154811 10989
rect 154839 10961 163625 10989
rect 163653 10961 163687 10989
rect 163715 10961 163749 10989
rect 163777 10961 163811 10989
rect 163839 10961 172625 10989
rect 172653 10961 172687 10989
rect 172715 10961 172749 10989
rect 172777 10961 172811 10989
rect 172839 10961 181625 10989
rect 181653 10961 181687 10989
rect 181715 10961 181749 10989
rect 181777 10961 181811 10989
rect 181839 10961 190625 10989
rect 190653 10961 190687 10989
rect 190715 10961 190749 10989
rect 190777 10961 190811 10989
rect 190839 10961 199625 10989
rect 199653 10961 199687 10989
rect 199715 10961 199749 10989
rect 199777 10961 199811 10989
rect 199839 10961 208625 10989
rect 208653 10961 208687 10989
rect 208715 10961 208749 10989
rect 208777 10961 208811 10989
rect 208839 10961 217625 10989
rect 217653 10961 217687 10989
rect 217715 10961 217749 10989
rect 217777 10961 217811 10989
rect 217839 10961 226625 10989
rect 226653 10961 226687 10989
rect 226715 10961 226749 10989
rect 226777 10961 226811 10989
rect 226839 10961 235625 10989
rect 235653 10961 235687 10989
rect 235715 10961 235749 10989
rect 235777 10961 235811 10989
rect 235839 10961 244625 10989
rect 244653 10961 244687 10989
rect 244715 10961 244749 10989
rect 244777 10961 244811 10989
rect 244839 10961 253625 10989
rect 253653 10961 253687 10989
rect 253715 10961 253749 10989
rect 253777 10961 253811 10989
rect 253839 10961 262625 10989
rect 262653 10961 262687 10989
rect 262715 10961 262749 10989
rect 262777 10961 262811 10989
rect 262839 10961 271625 10989
rect 271653 10961 271687 10989
rect 271715 10961 271749 10989
rect 271777 10961 271811 10989
rect 271839 10961 280625 10989
rect 280653 10961 280687 10989
rect 280715 10961 280749 10989
rect 280777 10961 280811 10989
rect 280839 10961 289625 10989
rect 289653 10961 289687 10989
rect 289715 10961 289749 10989
rect 289777 10961 289811 10989
rect 289839 10961 298248 10989
rect 298276 10961 298310 10989
rect 298338 10961 298372 10989
rect 298400 10961 298434 10989
rect 298462 10961 298990 10989
rect -958 10913 298990 10961
rect -958 5175 298990 5223
rect -958 5147 -910 5175
rect -882 5147 -848 5175
rect -820 5147 -786 5175
rect -758 5147 -724 5175
rect -696 5147 3485 5175
rect 3513 5147 3547 5175
rect 3575 5147 3609 5175
rect 3637 5147 3671 5175
rect 3699 5147 12485 5175
rect 12513 5147 12547 5175
rect 12575 5147 12609 5175
rect 12637 5147 12671 5175
rect 12699 5147 21485 5175
rect 21513 5147 21547 5175
rect 21575 5147 21609 5175
rect 21637 5147 21671 5175
rect 21699 5147 30485 5175
rect 30513 5147 30547 5175
rect 30575 5147 30609 5175
rect 30637 5147 30671 5175
rect 30699 5147 39485 5175
rect 39513 5147 39547 5175
rect 39575 5147 39609 5175
rect 39637 5147 39671 5175
rect 39699 5147 48485 5175
rect 48513 5147 48547 5175
rect 48575 5147 48609 5175
rect 48637 5147 48671 5175
rect 48699 5147 57485 5175
rect 57513 5147 57547 5175
rect 57575 5147 57609 5175
rect 57637 5147 57671 5175
rect 57699 5147 66485 5175
rect 66513 5147 66547 5175
rect 66575 5147 66609 5175
rect 66637 5147 66671 5175
rect 66699 5147 75485 5175
rect 75513 5147 75547 5175
rect 75575 5147 75609 5175
rect 75637 5147 75671 5175
rect 75699 5147 84485 5175
rect 84513 5147 84547 5175
rect 84575 5147 84609 5175
rect 84637 5147 84671 5175
rect 84699 5147 93485 5175
rect 93513 5147 93547 5175
rect 93575 5147 93609 5175
rect 93637 5147 93671 5175
rect 93699 5147 102485 5175
rect 102513 5147 102547 5175
rect 102575 5147 102609 5175
rect 102637 5147 102671 5175
rect 102699 5147 111485 5175
rect 111513 5147 111547 5175
rect 111575 5147 111609 5175
rect 111637 5147 111671 5175
rect 111699 5147 120485 5175
rect 120513 5147 120547 5175
rect 120575 5147 120609 5175
rect 120637 5147 120671 5175
rect 120699 5147 129485 5175
rect 129513 5147 129547 5175
rect 129575 5147 129609 5175
rect 129637 5147 129671 5175
rect 129699 5147 138485 5175
rect 138513 5147 138547 5175
rect 138575 5147 138609 5175
rect 138637 5147 138671 5175
rect 138699 5147 147485 5175
rect 147513 5147 147547 5175
rect 147575 5147 147609 5175
rect 147637 5147 147671 5175
rect 147699 5147 156485 5175
rect 156513 5147 156547 5175
rect 156575 5147 156609 5175
rect 156637 5147 156671 5175
rect 156699 5147 165485 5175
rect 165513 5147 165547 5175
rect 165575 5147 165609 5175
rect 165637 5147 165671 5175
rect 165699 5147 174485 5175
rect 174513 5147 174547 5175
rect 174575 5147 174609 5175
rect 174637 5147 174671 5175
rect 174699 5147 183485 5175
rect 183513 5147 183547 5175
rect 183575 5147 183609 5175
rect 183637 5147 183671 5175
rect 183699 5147 192485 5175
rect 192513 5147 192547 5175
rect 192575 5147 192609 5175
rect 192637 5147 192671 5175
rect 192699 5147 201485 5175
rect 201513 5147 201547 5175
rect 201575 5147 201609 5175
rect 201637 5147 201671 5175
rect 201699 5147 210485 5175
rect 210513 5147 210547 5175
rect 210575 5147 210609 5175
rect 210637 5147 210671 5175
rect 210699 5147 219485 5175
rect 219513 5147 219547 5175
rect 219575 5147 219609 5175
rect 219637 5147 219671 5175
rect 219699 5147 228485 5175
rect 228513 5147 228547 5175
rect 228575 5147 228609 5175
rect 228637 5147 228671 5175
rect 228699 5147 237485 5175
rect 237513 5147 237547 5175
rect 237575 5147 237609 5175
rect 237637 5147 237671 5175
rect 237699 5147 246485 5175
rect 246513 5147 246547 5175
rect 246575 5147 246609 5175
rect 246637 5147 246671 5175
rect 246699 5147 255485 5175
rect 255513 5147 255547 5175
rect 255575 5147 255609 5175
rect 255637 5147 255671 5175
rect 255699 5147 264485 5175
rect 264513 5147 264547 5175
rect 264575 5147 264609 5175
rect 264637 5147 264671 5175
rect 264699 5147 273485 5175
rect 273513 5147 273547 5175
rect 273575 5147 273609 5175
rect 273637 5147 273671 5175
rect 273699 5147 282485 5175
rect 282513 5147 282547 5175
rect 282575 5147 282609 5175
rect 282637 5147 282671 5175
rect 282699 5147 291485 5175
rect 291513 5147 291547 5175
rect 291575 5147 291609 5175
rect 291637 5147 291671 5175
rect 291699 5147 298728 5175
rect 298756 5147 298790 5175
rect 298818 5147 298852 5175
rect 298880 5147 298914 5175
rect 298942 5147 298990 5175
rect -958 5113 298990 5147
rect -958 5085 -910 5113
rect -882 5085 -848 5113
rect -820 5085 -786 5113
rect -758 5085 -724 5113
rect -696 5085 3485 5113
rect 3513 5085 3547 5113
rect 3575 5085 3609 5113
rect 3637 5085 3671 5113
rect 3699 5085 12485 5113
rect 12513 5085 12547 5113
rect 12575 5085 12609 5113
rect 12637 5085 12671 5113
rect 12699 5085 21485 5113
rect 21513 5085 21547 5113
rect 21575 5085 21609 5113
rect 21637 5085 21671 5113
rect 21699 5085 30485 5113
rect 30513 5085 30547 5113
rect 30575 5085 30609 5113
rect 30637 5085 30671 5113
rect 30699 5085 39485 5113
rect 39513 5085 39547 5113
rect 39575 5085 39609 5113
rect 39637 5085 39671 5113
rect 39699 5085 48485 5113
rect 48513 5085 48547 5113
rect 48575 5085 48609 5113
rect 48637 5085 48671 5113
rect 48699 5085 57485 5113
rect 57513 5085 57547 5113
rect 57575 5085 57609 5113
rect 57637 5085 57671 5113
rect 57699 5085 66485 5113
rect 66513 5085 66547 5113
rect 66575 5085 66609 5113
rect 66637 5085 66671 5113
rect 66699 5085 75485 5113
rect 75513 5085 75547 5113
rect 75575 5085 75609 5113
rect 75637 5085 75671 5113
rect 75699 5085 84485 5113
rect 84513 5085 84547 5113
rect 84575 5085 84609 5113
rect 84637 5085 84671 5113
rect 84699 5085 93485 5113
rect 93513 5085 93547 5113
rect 93575 5085 93609 5113
rect 93637 5085 93671 5113
rect 93699 5085 102485 5113
rect 102513 5085 102547 5113
rect 102575 5085 102609 5113
rect 102637 5085 102671 5113
rect 102699 5085 111485 5113
rect 111513 5085 111547 5113
rect 111575 5085 111609 5113
rect 111637 5085 111671 5113
rect 111699 5085 120485 5113
rect 120513 5085 120547 5113
rect 120575 5085 120609 5113
rect 120637 5085 120671 5113
rect 120699 5085 129485 5113
rect 129513 5085 129547 5113
rect 129575 5085 129609 5113
rect 129637 5085 129671 5113
rect 129699 5085 138485 5113
rect 138513 5085 138547 5113
rect 138575 5085 138609 5113
rect 138637 5085 138671 5113
rect 138699 5085 147485 5113
rect 147513 5085 147547 5113
rect 147575 5085 147609 5113
rect 147637 5085 147671 5113
rect 147699 5085 156485 5113
rect 156513 5085 156547 5113
rect 156575 5085 156609 5113
rect 156637 5085 156671 5113
rect 156699 5085 165485 5113
rect 165513 5085 165547 5113
rect 165575 5085 165609 5113
rect 165637 5085 165671 5113
rect 165699 5085 174485 5113
rect 174513 5085 174547 5113
rect 174575 5085 174609 5113
rect 174637 5085 174671 5113
rect 174699 5085 183485 5113
rect 183513 5085 183547 5113
rect 183575 5085 183609 5113
rect 183637 5085 183671 5113
rect 183699 5085 192485 5113
rect 192513 5085 192547 5113
rect 192575 5085 192609 5113
rect 192637 5085 192671 5113
rect 192699 5085 201485 5113
rect 201513 5085 201547 5113
rect 201575 5085 201609 5113
rect 201637 5085 201671 5113
rect 201699 5085 210485 5113
rect 210513 5085 210547 5113
rect 210575 5085 210609 5113
rect 210637 5085 210671 5113
rect 210699 5085 219485 5113
rect 219513 5085 219547 5113
rect 219575 5085 219609 5113
rect 219637 5085 219671 5113
rect 219699 5085 228485 5113
rect 228513 5085 228547 5113
rect 228575 5085 228609 5113
rect 228637 5085 228671 5113
rect 228699 5085 237485 5113
rect 237513 5085 237547 5113
rect 237575 5085 237609 5113
rect 237637 5085 237671 5113
rect 237699 5085 246485 5113
rect 246513 5085 246547 5113
rect 246575 5085 246609 5113
rect 246637 5085 246671 5113
rect 246699 5085 255485 5113
rect 255513 5085 255547 5113
rect 255575 5085 255609 5113
rect 255637 5085 255671 5113
rect 255699 5085 264485 5113
rect 264513 5085 264547 5113
rect 264575 5085 264609 5113
rect 264637 5085 264671 5113
rect 264699 5085 273485 5113
rect 273513 5085 273547 5113
rect 273575 5085 273609 5113
rect 273637 5085 273671 5113
rect 273699 5085 282485 5113
rect 282513 5085 282547 5113
rect 282575 5085 282609 5113
rect 282637 5085 282671 5113
rect 282699 5085 291485 5113
rect 291513 5085 291547 5113
rect 291575 5085 291609 5113
rect 291637 5085 291671 5113
rect 291699 5085 298728 5113
rect 298756 5085 298790 5113
rect 298818 5085 298852 5113
rect 298880 5085 298914 5113
rect 298942 5085 298990 5113
rect -958 5051 298990 5085
rect -958 5023 -910 5051
rect -882 5023 -848 5051
rect -820 5023 -786 5051
rect -758 5023 -724 5051
rect -696 5023 3485 5051
rect 3513 5023 3547 5051
rect 3575 5023 3609 5051
rect 3637 5023 3671 5051
rect 3699 5023 12485 5051
rect 12513 5023 12547 5051
rect 12575 5023 12609 5051
rect 12637 5023 12671 5051
rect 12699 5023 21485 5051
rect 21513 5023 21547 5051
rect 21575 5023 21609 5051
rect 21637 5023 21671 5051
rect 21699 5023 30485 5051
rect 30513 5023 30547 5051
rect 30575 5023 30609 5051
rect 30637 5023 30671 5051
rect 30699 5023 39485 5051
rect 39513 5023 39547 5051
rect 39575 5023 39609 5051
rect 39637 5023 39671 5051
rect 39699 5023 48485 5051
rect 48513 5023 48547 5051
rect 48575 5023 48609 5051
rect 48637 5023 48671 5051
rect 48699 5023 57485 5051
rect 57513 5023 57547 5051
rect 57575 5023 57609 5051
rect 57637 5023 57671 5051
rect 57699 5023 66485 5051
rect 66513 5023 66547 5051
rect 66575 5023 66609 5051
rect 66637 5023 66671 5051
rect 66699 5023 75485 5051
rect 75513 5023 75547 5051
rect 75575 5023 75609 5051
rect 75637 5023 75671 5051
rect 75699 5023 84485 5051
rect 84513 5023 84547 5051
rect 84575 5023 84609 5051
rect 84637 5023 84671 5051
rect 84699 5023 93485 5051
rect 93513 5023 93547 5051
rect 93575 5023 93609 5051
rect 93637 5023 93671 5051
rect 93699 5023 102485 5051
rect 102513 5023 102547 5051
rect 102575 5023 102609 5051
rect 102637 5023 102671 5051
rect 102699 5023 111485 5051
rect 111513 5023 111547 5051
rect 111575 5023 111609 5051
rect 111637 5023 111671 5051
rect 111699 5023 120485 5051
rect 120513 5023 120547 5051
rect 120575 5023 120609 5051
rect 120637 5023 120671 5051
rect 120699 5023 129485 5051
rect 129513 5023 129547 5051
rect 129575 5023 129609 5051
rect 129637 5023 129671 5051
rect 129699 5023 138485 5051
rect 138513 5023 138547 5051
rect 138575 5023 138609 5051
rect 138637 5023 138671 5051
rect 138699 5023 147485 5051
rect 147513 5023 147547 5051
rect 147575 5023 147609 5051
rect 147637 5023 147671 5051
rect 147699 5023 156485 5051
rect 156513 5023 156547 5051
rect 156575 5023 156609 5051
rect 156637 5023 156671 5051
rect 156699 5023 165485 5051
rect 165513 5023 165547 5051
rect 165575 5023 165609 5051
rect 165637 5023 165671 5051
rect 165699 5023 174485 5051
rect 174513 5023 174547 5051
rect 174575 5023 174609 5051
rect 174637 5023 174671 5051
rect 174699 5023 183485 5051
rect 183513 5023 183547 5051
rect 183575 5023 183609 5051
rect 183637 5023 183671 5051
rect 183699 5023 192485 5051
rect 192513 5023 192547 5051
rect 192575 5023 192609 5051
rect 192637 5023 192671 5051
rect 192699 5023 201485 5051
rect 201513 5023 201547 5051
rect 201575 5023 201609 5051
rect 201637 5023 201671 5051
rect 201699 5023 210485 5051
rect 210513 5023 210547 5051
rect 210575 5023 210609 5051
rect 210637 5023 210671 5051
rect 210699 5023 219485 5051
rect 219513 5023 219547 5051
rect 219575 5023 219609 5051
rect 219637 5023 219671 5051
rect 219699 5023 228485 5051
rect 228513 5023 228547 5051
rect 228575 5023 228609 5051
rect 228637 5023 228671 5051
rect 228699 5023 237485 5051
rect 237513 5023 237547 5051
rect 237575 5023 237609 5051
rect 237637 5023 237671 5051
rect 237699 5023 246485 5051
rect 246513 5023 246547 5051
rect 246575 5023 246609 5051
rect 246637 5023 246671 5051
rect 246699 5023 255485 5051
rect 255513 5023 255547 5051
rect 255575 5023 255609 5051
rect 255637 5023 255671 5051
rect 255699 5023 264485 5051
rect 264513 5023 264547 5051
rect 264575 5023 264609 5051
rect 264637 5023 264671 5051
rect 264699 5023 273485 5051
rect 273513 5023 273547 5051
rect 273575 5023 273609 5051
rect 273637 5023 273671 5051
rect 273699 5023 282485 5051
rect 282513 5023 282547 5051
rect 282575 5023 282609 5051
rect 282637 5023 282671 5051
rect 282699 5023 291485 5051
rect 291513 5023 291547 5051
rect 291575 5023 291609 5051
rect 291637 5023 291671 5051
rect 291699 5023 298728 5051
rect 298756 5023 298790 5051
rect 298818 5023 298852 5051
rect 298880 5023 298914 5051
rect 298942 5023 298990 5051
rect -958 4989 298990 5023
rect -958 4961 -910 4989
rect -882 4961 -848 4989
rect -820 4961 -786 4989
rect -758 4961 -724 4989
rect -696 4961 3485 4989
rect 3513 4961 3547 4989
rect 3575 4961 3609 4989
rect 3637 4961 3671 4989
rect 3699 4961 12485 4989
rect 12513 4961 12547 4989
rect 12575 4961 12609 4989
rect 12637 4961 12671 4989
rect 12699 4961 21485 4989
rect 21513 4961 21547 4989
rect 21575 4961 21609 4989
rect 21637 4961 21671 4989
rect 21699 4961 30485 4989
rect 30513 4961 30547 4989
rect 30575 4961 30609 4989
rect 30637 4961 30671 4989
rect 30699 4961 39485 4989
rect 39513 4961 39547 4989
rect 39575 4961 39609 4989
rect 39637 4961 39671 4989
rect 39699 4961 48485 4989
rect 48513 4961 48547 4989
rect 48575 4961 48609 4989
rect 48637 4961 48671 4989
rect 48699 4961 57485 4989
rect 57513 4961 57547 4989
rect 57575 4961 57609 4989
rect 57637 4961 57671 4989
rect 57699 4961 66485 4989
rect 66513 4961 66547 4989
rect 66575 4961 66609 4989
rect 66637 4961 66671 4989
rect 66699 4961 75485 4989
rect 75513 4961 75547 4989
rect 75575 4961 75609 4989
rect 75637 4961 75671 4989
rect 75699 4961 84485 4989
rect 84513 4961 84547 4989
rect 84575 4961 84609 4989
rect 84637 4961 84671 4989
rect 84699 4961 93485 4989
rect 93513 4961 93547 4989
rect 93575 4961 93609 4989
rect 93637 4961 93671 4989
rect 93699 4961 102485 4989
rect 102513 4961 102547 4989
rect 102575 4961 102609 4989
rect 102637 4961 102671 4989
rect 102699 4961 111485 4989
rect 111513 4961 111547 4989
rect 111575 4961 111609 4989
rect 111637 4961 111671 4989
rect 111699 4961 120485 4989
rect 120513 4961 120547 4989
rect 120575 4961 120609 4989
rect 120637 4961 120671 4989
rect 120699 4961 129485 4989
rect 129513 4961 129547 4989
rect 129575 4961 129609 4989
rect 129637 4961 129671 4989
rect 129699 4961 138485 4989
rect 138513 4961 138547 4989
rect 138575 4961 138609 4989
rect 138637 4961 138671 4989
rect 138699 4961 147485 4989
rect 147513 4961 147547 4989
rect 147575 4961 147609 4989
rect 147637 4961 147671 4989
rect 147699 4961 156485 4989
rect 156513 4961 156547 4989
rect 156575 4961 156609 4989
rect 156637 4961 156671 4989
rect 156699 4961 165485 4989
rect 165513 4961 165547 4989
rect 165575 4961 165609 4989
rect 165637 4961 165671 4989
rect 165699 4961 174485 4989
rect 174513 4961 174547 4989
rect 174575 4961 174609 4989
rect 174637 4961 174671 4989
rect 174699 4961 183485 4989
rect 183513 4961 183547 4989
rect 183575 4961 183609 4989
rect 183637 4961 183671 4989
rect 183699 4961 192485 4989
rect 192513 4961 192547 4989
rect 192575 4961 192609 4989
rect 192637 4961 192671 4989
rect 192699 4961 201485 4989
rect 201513 4961 201547 4989
rect 201575 4961 201609 4989
rect 201637 4961 201671 4989
rect 201699 4961 210485 4989
rect 210513 4961 210547 4989
rect 210575 4961 210609 4989
rect 210637 4961 210671 4989
rect 210699 4961 219485 4989
rect 219513 4961 219547 4989
rect 219575 4961 219609 4989
rect 219637 4961 219671 4989
rect 219699 4961 228485 4989
rect 228513 4961 228547 4989
rect 228575 4961 228609 4989
rect 228637 4961 228671 4989
rect 228699 4961 237485 4989
rect 237513 4961 237547 4989
rect 237575 4961 237609 4989
rect 237637 4961 237671 4989
rect 237699 4961 246485 4989
rect 246513 4961 246547 4989
rect 246575 4961 246609 4989
rect 246637 4961 246671 4989
rect 246699 4961 255485 4989
rect 255513 4961 255547 4989
rect 255575 4961 255609 4989
rect 255637 4961 255671 4989
rect 255699 4961 264485 4989
rect 264513 4961 264547 4989
rect 264575 4961 264609 4989
rect 264637 4961 264671 4989
rect 264699 4961 273485 4989
rect 273513 4961 273547 4989
rect 273575 4961 273609 4989
rect 273637 4961 273671 4989
rect 273699 4961 282485 4989
rect 282513 4961 282547 4989
rect 282575 4961 282609 4989
rect 282637 4961 282671 4989
rect 282699 4961 291485 4989
rect 291513 4961 291547 4989
rect 291575 4961 291609 4989
rect 291637 4961 291671 4989
rect 291699 4961 298728 4989
rect 298756 4961 298790 4989
rect 298818 4961 298852 4989
rect 298880 4961 298914 4989
rect 298942 4961 298990 4989
rect -958 4913 298990 4961
rect -958 2175 298990 2223
rect -958 2147 -430 2175
rect -402 2147 -368 2175
rect -340 2147 -306 2175
rect -278 2147 -244 2175
rect -216 2147 1625 2175
rect 1653 2147 1687 2175
rect 1715 2147 1749 2175
rect 1777 2147 1811 2175
rect 1839 2147 10625 2175
rect 10653 2147 10687 2175
rect 10715 2147 10749 2175
rect 10777 2147 10811 2175
rect 10839 2147 19625 2175
rect 19653 2147 19687 2175
rect 19715 2147 19749 2175
rect 19777 2147 19811 2175
rect 19839 2147 28625 2175
rect 28653 2147 28687 2175
rect 28715 2147 28749 2175
rect 28777 2147 28811 2175
rect 28839 2147 37625 2175
rect 37653 2147 37687 2175
rect 37715 2147 37749 2175
rect 37777 2147 37811 2175
rect 37839 2147 46625 2175
rect 46653 2147 46687 2175
rect 46715 2147 46749 2175
rect 46777 2147 46811 2175
rect 46839 2147 55625 2175
rect 55653 2147 55687 2175
rect 55715 2147 55749 2175
rect 55777 2147 55811 2175
rect 55839 2147 64625 2175
rect 64653 2147 64687 2175
rect 64715 2147 64749 2175
rect 64777 2147 64811 2175
rect 64839 2147 73625 2175
rect 73653 2147 73687 2175
rect 73715 2147 73749 2175
rect 73777 2147 73811 2175
rect 73839 2147 82625 2175
rect 82653 2147 82687 2175
rect 82715 2147 82749 2175
rect 82777 2147 82811 2175
rect 82839 2147 91625 2175
rect 91653 2147 91687 2175
rect 91715 2147 91749 2175
rect 91777 2147 91811 2175
rect 91839 2147 100625 2175
rect 100653 2147 100687 2175
rect 100715 2147 100749 2175
rect 100777 2147 100811 2175
rect 100839 2147 109625 2175
rect 109653 2147 109687 2175
rect 109715 2147 109749 2175
rect 109777 2147 109811 2175
rect 109839 2147 118625 2175
rect 118653 2147 118687 2175
rect 118715 2147 118749 2175
rect 118777 2147 118811 2175
rect 118839 2147 127625 2175
rect 127653 2147 127687 2175
rect 127715 2147 127749 2175
rect 127777 2147 127811 2175
rect 127839 2147 136625 2175
rect 136653 2147 136687 2175
rect 136715 2147 136749 2175
rect 136777 2147 136811 2175
rect 136839 2147 145625 2175
rect 145653 2147 145687 2175
rect 145715 2147 145749 2175
rect 145777 2147 145811 2175
rect 145839 2147 154625 2175
rect 154653 2147 154687 2175
rect 154715 2147 154749 2175
rect 154777 2147 154811 2175
rect 154839 2147 163625 2175
rect 163653 2147 163687 2175
rect 163715 2147 163749 2175
rect 163777 2147 163811 2175
rect 163839 2147 172625 2175
rect 172653 2147 172687 2175
rect 172715 2147 172749 2175
rect 172777 2147 172811 2175
rect 172839 2147 181625 2175
rect 181653 2147 181687 2175
rect 181715 2147 181749 2175
rect 181777 2147 181811 2175
rect 181839 2147 190625 2175
rect 190653 2147 190687 2175
rect 190715 2147 190749 2175
rect 190777 2147 190811 2175
rect 190839 2147 199625 2175
rect 199653 2147 199687 2175
rect 199715 2147 199749 2175
rect 199777 2147 199811 2175
rect 199839 2147 208625 2175
rect 208653 2147 208687 2175
rect 208715 2147 208749 2175
rect 208777 2147 208811 2175
rect 208839 2147 217625 2175
rect 217653 2147 217687 2175
rect 217715 2147 217749 2175
rect 217777 2147 217811 2175
rect 217839 2147 226625 2175
rect 226653 2147 226687 2175
rect 226715 2147 226749 2175
rect 226777 2147 226811 2175
rect 226839 2147 235625 2175
rect 235653 2147 235687 2175
rect 235715 2147 235749 2175
rect 235777 2147 235811 2175
rect 235839 2147 244625 2175
rect 244653 2147 244687 2175
rect 244715 2147 244749 2175
rect 244777 2147 244811 2175
rect 244839 2147 253625 2175
rect 253653 2147 253687 2175
rect 253715 2147 253749 2175
rect 253777 2147 253811 2175
rect 253839 2147 262625 2175
rect 262653 2147 262687 2175
rect 262715 2147 262749 2175
rect 262777 2147 262811 2175
rect 262839 2147 271625 2175
rect 271653 2147 271687 2175
rect 271715 2147 271749 2175
rect 271777 2147 271811 2175
rect 271839 2147 280625 2175
rect 280653 2147 280687 2175
rect 280715 2147 280749 2175
rect 280777 2147 280811 2175
rect 280839 2147 289625 2175
rect 289653 2147 289687 2175
rect 289715 2147 289749 2175
rect 289777 2147 289811 2175
rect 289839 2147 298248 2175
rect 298276 2147 298310 2175
rect 298338 2147 298372 2175
rect 298400 2147 298434 2175
rect 298462 2147 298990 2175
rect -958 2113 298990 2147
rect -958 2085 -430 2113
rect -402 2085 -368 2113
rect -340 2085 -306 2113
rect -278 2085 -244 2113
rect -216 2085 1625 2113
rect 1653 2085 1687 2113
rect 1715 2085 1749 2113
rect 1777 2085 1811 2113
rect 1839 2085 10625 2113
rect 10653 2085 10687 2113
rect 10715 2085 10749 2113
rect 10777 2085 10811 2113
rect 10839 2085 19625 2113
rect 19653 2085 19687 2113
rect 19715 2085 19749 2113
rect 19777 2085 19811 2113
rect 19839 2085 28625 2113
rect 28653 2085 28687 2113
rect 28715 2085 28749 2113
rect 28777 2085 28811 2113
rect 28839 2085 37625 2113
rect 37653 2085 37687 2113
rect 37715 2085 37749 2113
rect 37777 2085 37811 2113
rect 37839 2085 46625 2113
rect 46653 2085 46687 2113
rect 46715 2085 46749 2113
rect 46777 2085 46811 2113
rect 46839 2085 55625 2113
rect 55653 2085 55687 2113
rect 55715 2085 55749 2113
rect 55777 2085 55811 2113
rect 55839 2085 64625 2113
rect 64653 2085 64687 2113
rect 64715 2085 64749 2113
rect 64777 2085 64811 2113
rect 64839 2085 73625 2113
rect 73653 2085 73687 2113
rect 73715 2085 73749 2113
rect 73777 2085 73811 2113
rect 73839 2085 82625 2113
rect 82653 2085 82687 2113
rect 82715 2085 82749 2113
rect 82777 2085 82811 2113
rect 82839 2085 91625 2113
rect 91653 2085 91687 2113
rect 91715 2085 91749 2113
rect 91777 2085 91811 2113
rect 91839 2085 100625 2113
rect 100653 2085 100687 2113
rect 100715 2085 100749 2113
rect 100777 2085 100811 2113
rect 100839 2085 109625 2113
rect 109653 2085 109687 2113
rect 109715 2085 109749 2113
rect 109777 2085 109811 2113
rect 109839 2085 118625 2113
rect 118653 2085 118687 2113
rect 118715 2085 118749 2113
rect 118777 2085 118811 2113
rect 118839 2085 127625 2113
rect 127653 2085 127687 2113
rect 127715 2085 127749 2113
rect 127777 2085 127811 2113
rect 127839 2085 136625 2113
rect 136653 2085 136687 2113
rect 136715 2085 136749 2113
rect 136777 2085 136811 2113
rect 136839 2085 145625 2113
rect 145653 2085 145687 2113
rect 145715 2085 145749 2113
rect 145777 2085 145811 2113
rect 145839 2085 154625 2113
rect 154653 2085 154687 2113
rect 154715 2085 154749 2113
rect 154777 2085 154811 2113
rect 154839 2085 163625 2113
rect 163653 2085 163687 2113
rect 163715 2085 163749 2113
rect 163777 2085 163811 2113
rect 163839 2085 172625 2113
rect 172653 2085 172687 2113
rect 172715 2085 172749 2113
rect 172777 2085 172811 2113
rect 172839 2085 181625 2113
rect 181653 2085 181687 2113
rect 181715 2085 181749 2113
rect 181777 2085 181811 2113
rect 181839 2085 190625 2113
rect 190653 2085 190687 2113
rect 190715 2085 190749 2113
rect 190777 2085 190811 2113
rect 190839 2085 199625 2113
rect 199653 2085 199687 2113
rect 199715 2085 199749 2113
rect 199777 2085 199811 2113
rect 199839 2085 208625 2113
rect 208653 2085 208687 2113
rect 208715 2085 208749 2113
rect 208777 2085 208811 2113
rect 208839 2085 217625 2113
rect 217653 2085 217687 2113
rect 217715 2085 217749 2113
rect 217777 2085 217811 2113
rect 217839 2085 226625 2113
rect 226653 2085 226687 2113
rect 226715 2085 226749 2113
rect 226777 2085 226811 2113
rect 226839 2085 235625 2113
rect 235653 2085 235687 2113
rect 235715 2085 235749 2113
rect 235777 2085 235811 2113
rect 235839 2085 244625 2113
rect 244653 2085 244687 2113
rect 244715 2085 244749 2113
rect 244777 2085 244811 2113
rect 244839 2085 253625 2113
rect 253653 2085 253687 2113
rect 253715 2085 253749 2113
rect 253777 2085 253811 2113
rect 253839 2085 262625 2113
rect 262653 2085 262687 2113
rect 262715 2085 262749 2113
rect 262777 2085 262811 2113
rect 262839 2085 271625 2113
rect 271653 2085 271687 2113
rect 271715 2085 271749 2113
rect 271777 2085 271811 2113
rect 271839 2085 280625 2113
rect 280653 2085 280687 2113
rect 280715 2085 280749 2113
rect 280777 2085 280811 2113
rect 280839 2085 289625 2113
rect 289653 2085 289687 2113
rect 289715 2085 289749 2113
rect 289777 2085 289811 2113
rect 289839 2085 298248 2113
rect 298276 2085 298310 2113
rect 298338 2085 298372 2113
rect 298400 2085 298434 2113
rect 298462 2085 298990 2113
rect -958 2051 298990 2085
rect -958 2023 -430 2051
rect -402 2023 -368 2051
rect -340 2023 -306 2051
rect -278 2023 -244 2051
rect -216 2023 1625 2051
rect 1653 2023 1687 2051
rect 1715 2023 1749 2051
rect 1777 2023 1811 2051
rect 1839 2023 10625 2051
rect 10653 2023 10687 2051
rect 10715 2023 10749 2051
rect 10777 2023 10811 2051
rect 10839 2023 19625 2051
rect 19653 2023 19687 2051
rect 19715 2023 19749 2051
rect 19777 2023 19811 2051
rect 19839 2023 28625 2051
rect 28653 2023 28687 2051
rect 28715 2023 28749 2051
rect 28777 2023 28811 2051
rect 28839 2023 37625 2051
rect 37653 2023 37687 2051
rect 37715 2023 37749 2051
rect 37777 2023 37811 2051
rect 37839 2023 46625 2051
rect 46653 2023 46687 2051
rect 46715 2023 46749 2051
rect 46777 2023 46811 2051
rect 46839 2023 55625 2051
rect 55653 2023 55687 2051
rect 55715 2023 55749 2051
rect 55777 2023 55811 2051
rect 55839 2023 64625 2051
rect 64653 2023 64687 2051
rect 64715 2023 64749 2051
rect 64777 2023 64811 2051
rect 64839 2023 73625 2051
rect 73653 2023 73687 2051
rect 73715 2023 73749 2051
rect 73777 2023 73811 2051
rect 73839 2023 82625 2051
rect 82653 2023 82687 2051
rect 82715 2023 82749 2051
rect 82777 2023 82811 2051
rect 82839 2023 91625 2051
rect 91653 2023 91687 2051
rect 91715 2023 91749 2051
rect 91777 2023 91811 2051
rect 91839 2023 100625 2051
rect 100653 2023 100687 2051
rect 100715 2023 100749 2051
rect 100777 2023 100811 2051
rect 100839 2023 109625 2051
rect 109653 2023 109687 2051
rect 109715 2023 109749 2051
rect 109777 2023 109811 2051
rect 109839 2023 118625 2051
rect 118653 2023 118687 2051
rect 118715 2023 118749 2051
rect 118777 2023 118811 2051
rect 118839 2023 127625 2051
rect 127653 2023 127687 2051
rect 127715 2023 127749 2051
rect 127777 2023 127811 2051
rect 127839 2023 136625 2051
rect 136653 2023 136687 2051
rect 136715 2023 136749 2051
rect 136777 2023 136811 2051
rect 136839 2023 145625 2051
rect 145653 2023 145687 2051
rect 145715 2023 145749 2051
rect 145777 2023 145811 2051
rect 145839 2023 154625 2051
rect 154653 2023 154687 2051
rect 154715 2023 154749 2051
rect 154777 2023 154811 2051
rect 154839 2023 163625 2051
rect 163653 2023 163687 2051
rect 163715 2023 163749 2051
rect 163777 2023 163811 2051
rect 163839 2023 172625 2051
rect 172653 2023 172687 2051
rect 172715 2023 172749 2051
rect 172777 2023 172811 2051
rect 172839 2023 181625 2051
rect 181653 2023 181687 2051
rect 181715 2023 181749 2051
rect 181777 2023 181811 2051
rect 181839 2023 190625 2051
rect 190653 2023 190687 2051
rect 190715 2023 190749 2051
rect 190777 2023 190811 2051
rect 190839 2023 199625 2051
rect 199653 2023 199687 2051
rect 199715 2023 199749 2051
rect 199777 2023 199811 2051
rect 199839 2023 208625 2051
rect 208653 2023 208687 2051
rect 208715 2023 208749 2051
rect 208777 2023 208811 2051
rect 208839 2023 217625 2051
rect 217653 2023 217687 2051
rect 217715 2023 217749 2051
rect 217777 2023 217811 2051
rect 217839 2023 226625 2051
rect 226653 2023 226687 2051
rect 226715 2023 226749 2051
rect 226777 2023 226811 2051
rect 226839 2023 235625 2051
rect 235653 2023 235687 2051
rect 235715 2023 235749 2051
rect 235777 2023 235811 2051
rect 235839 2023 244625 2051
rect 244653 2023 244687 2051
rect 244715 2023 244749 2051
rect 244777 2023 244811 2051
rect 244839 2023 253625 2051
rect 253653 2023 253687 2051
rect 253715 2023 253749 2051
rect 253777 2023 253811 2051
rect 253839 2023 262625 2051
rect 262653 2023 262687 2051
rect 262715 2023 262749 2051
rect 262777 2023 262811 2051
rect 262839 2023 271625 2051
rect 271653 2023 271687 2051
rect 271715 2023 271749 2051
rect 271777 2023 271811 2051
rect 271839 2023 280625 2051
rect 280653 2023 280687 2051
rect 280715 2023 280749 2051
rect 280777 2023 280811 2051
rect 280839 2023 289625 2051
rect 289653 2023 289687 2051
rect 289715 2023 289749 2051
rect 289777 2023 289811 2051
rect 289839 2023 298248 2051
rect 298276 2023 298310 2051
rect 298338 2023 298372 2051
rect 298400 2023 298434 2051
rect 298462 2023 298990 2051
rect -958 1989 298990 2023
rect -958 1961 -430 1989
rect -402 1961 -368 1989
rect -340 1961 -306 1989
rect -278 1961 -244 1989
rect -216 1961 1625 1989
rect 1653 1961 1687 1989
rect 1715 1961 1749 1989
rect 1777 1961 1811 1989
rect 1839 1961 10625 1989
rect 10653 1961 10687 1989
rect 10715 1961 10749 1989
rect 10777 1961 10811 1989
rect 10839 1961 19625 1989
rect 19653 1961 19687 1989
rect 19715 1961 19749 1989
rect 19777 1961 19811 1989
rect 19839 1961 28625 1989
rect 28653 1961 28687 1989
rect 28715 1961 28749 1989
rect 28777 1961 28811 1989
rect 28839 1961 37625 1989
rect 37653 1961 37687 1989
rect 37715 1961 37749 1989
rect 37777 1961 37811 1989
rect 37839 1961 46625 1989
rect 46653 1961 46687 1989
rect 46715 1961 46749 1989
rect 46777 1961 46811 1989
rect 46839 1961 55625 1989
rect 55653 1961 55687 1989
rect 55715 1961 55749 1989
rect 55777 1961 55811 1989
rect 55839 1961 64625 1989
rect 64653 1961 64687 1989
rect 64715 1961 64749 1989
rect 64777 1961 64811 1989
rect 64839 1961 73625 1989
rect 73653 1961 73687 1989
rect 73715 1961 73749 1989
rect 73777 1961 73811 1989
rect 73839 1961 82625 1989
rect 82653 1961 82687 1989
rect 82715 1961 82749 1989
rect 82777 1961 82811 1989
rect 82839 1961 91625 1989
rect 91653 1961 91687 1989
rect 91715 1961 91749 1989
rect 91777 1961 91811 1989
rect 91839 1961 100625 1989
rect 100653 1961 100687 1989
rect 100715 1961 100749 1989
rect 100777 1961 100811 1989
rect 100839 1961 109625 1989
rect 109653 1961 109687 1989
rect 109715 1961 109749 1989
rect 109777 1961 109811 1989
rect 109839 1961 118625 1989
rect 118653 1961 118687 1989
rect 118715 1961 118749 1989
rect 118777 1961 118811 1989
rect 118839 1961 127625 1989
rect 127653 1961 127687 1989
rect 127715 1961 127749 1989
rect 127777 1961 127811 1989
rect 127839 1961 136625 1989
rect 136653 1961 136687 1989
rect 136715 1961 136749 1989
rect 136777 1961 136811 1989
rect 136839 1961 145625 1989
rect 145653 1961 145687 1989
rect 145715 1961 145749 1989
rect 145777 1961 145811 1989
rect 145839 1961 154625 1989
rect 154653 1961 154687 1989
rect 154715 1961 154749 1989
rect 154777 1961 154811 1989
rect 154839 1961 163625 1989
rect 163653 1961 163687 1989
rect 163715 1961 163749 1989
rect 163777 1961 163811 1989
rect 163839 1961 172625 1989
rect 172653 1961 172687 1989
rect 172715 1961 172749 1989
rect 172777 1961 172811 1989
rect 172839 1961 181625 1989
rect 181653 1961 181687 1989
rect 181715 1961 181749 1989
rect 181777 1961 181811 1989
rect 181839 1961 190625 1989
rect 190653 1961 190687 1989
rect 190715 1961 190749 1989
rect 190777 1961 190811 1989
rect 190839 1961 199625 1989
rect 199653 1961 199687 1989
rect 199715 1961 199749 1989
rect 199777 1961 199811 1989
rect 199839 1961 208625 1989
rect 208653 1961 208687 1989
rect 208715 1961 208749 1989
rect 208777 1961 208811 1989
rect 208839 1961 217625 1989
rect 217653 1961 217687 1989
rect 217715 1961 217749 1989
rect 217777 1961 217811 1989
rect 217839 1961 226625 1989
rect 226653 1961 226687 1989
rect 226715 1961 226749 1989
rect 226777 1961 226811 1989
rect 226839 1961 235625 1989
rect 235653 1961 235687 1989
rect 235715 1961 235749 1989
rect 235777 1961 235811 1989
rect 235839 1961 244625 1989
rect 244653 1961 244687 1989
rect 244715 1961 244749 1989
rect 244777 1961 244811 1989
rect 244839 1961 253625 1989
rect 253653 1961 253687 1989
rect 253715 1961 253749 1989
rect 253777 1961 253811 1989
rect 253839 1961 262625 1989
rect 262653 1961 262687 1989
rect 262715 1961 262749 1989
rect 262777 1961 262811 1989
rect 262839 1961 271625 1989
rect 271653 1961 271687 1989
rect 271715 1961 271749 1989
rect 271777 1961 271811 1989
rect 271839 1961 280625 1989
rect 280653 1961 280687 1989
rect 280715 1961 280749 1989
rect 280777 1961 280811 1989
rect 280839 1961 289625 1989
rect 289653 1961 289687 1989
rect 289715 1961 289749 1989
rect 289777 1961 289811 1989
rect 289839 1961 298248 1989
rect 298276 1961 298310 1989
rect 298338 1961 298372 1989
rect 298400 1961 298434 1989
rect 298462 1961 298990 1989
rect -958 1913 298990 1961
rect -478 -80 298510 -32
rect -478 -108 -430 -80
rect -402 -108 -368 -80
rect -340 -108 -306 -80
rect -278 -108 -244 -80
rect -216 -108 1625 -80
rect 1653 -108 1687 -80
rect 1715 -108 1749 -80
rect 1777 -108 1811 -80
rect 1839 -108 10625 -80
rect 10653 -108 10687 -80
rect 10715 -108 10749 -80
rect 10777 -108 10811 -80
rect 10839 -108 19625 -80
rect 19653 -108 19687 -80
rect 19715 -108 19749 -80
rect 19777 -108 19811 -80
rect 19839 -108 28625 -80
rect 28653 -108 28687 -80
rect 28715 -108 28749 -80
rect 28777 -108 28811 -80
rect 28839 -108 37625 -80
rect 37653 -108 37687 -80
rect 37715 -108 37749 -80
rect 37777 -108 37811 -80
rect 37839 -108 46625 -80
rect 46653 -108 46687 -80
rect 46715 -108 46749 -80
rect 46777 -108 46811 -80
rect 46839 -108 55625 -80
rect 55653 -108 55687 -80
rect 55715 -108 55749 -80
rect 55777 -108 55811 -80
rect 55839 -108 64625 -80
rect 64653 -108 64687 -80
rect 64715 -108 64749 -80
rect 64777 -108 64811 -80
rect 64839 -108 73625 -80
rect 73653 -108 73687 -80
rect 73715 -108 73749 -80
rect 73777 -108 73811 -80
rect 73839 -108 82625 -80
rect 82653 -108 82687 -80
rect 82715 -108 82749 -80
rect 82777 -108 82811 -80
rect 82839 -108 91625 -80
rect 91653 -108 91687 -80
rect 91715 -108 91749 -80
rect 91777 -108 91811 -80
rect 91839 -108 100625 -80
rect 100653 -108 100687 -80
rect 100715 -108 100749 -80
rect 100777 -108 100811 -80
rect 100839 -108 109625 -80
rect 109653 -108 109687 -80
rect 109715 -108 109749 -80
rect 109777 -108 109811 -80
rect 109839 -108 118625 -80
rect 118653 -108 118687 -80
rect 118715 -108 118749 -80
rect 118777 -108 118811 -80
rect 118839 -108 127625 -80
rect 127653 -108 127687 -80
rect 127715 -108 127749 -80
rect 127777 -108 127811 -80
rect 127839 -108 136625 -80
rect 136653 -108 136687 -80
rect 136715 -108 136749 -80
rect 136777 -108 136811 -80
rect 136839 -108 145625 -80
rect 145653 -108 145687 -80
rect 145715 -108 145749 -80
rect 145777 -108 145811 -80
rect 145839 -108 154625 -80
rect 154653 -108 154687 -80
rect 154715 -108 154749 -80
rect 154777 -108 154811 -80
rect 154839 -108 163625 -80
rect 163653 -108 163687 -80
rect 163715 -108 163749 -80
rect 163777 -108 163811 -80
rect 163839 -108 172625 -80
rect 172653 -108 172687 -80
rect 172715 -108 172749 -80
rect 172777 -108 172811 -80
rect 172839 -108 181625 -80
rect 181653 -108 181687 -80
rect 181715 -108 181749 -80
rect 181777 -108 181811 -80
rect 181839 -108 190625 -80
rect 190653 -108 190687 -80
rect 190715 -108 190749 -80
rect 190777 -108 190811 -80
rect 190839 -108 199625 -80
rect 199653 -108 199687 -80
rect 199715 -108 199749 -80
rect 199777 -108 199811 -80
rect 199839 -108 208625 -80
rect 208653 -108 208687 -80
rect 208715 -108 208749 -80
rect 208777 -108 208811 -80
rect 208839 -108 217625 -80
rect 217653 -108 217687 -80
rect 217715 -108 217749 -80
rect 217777 -108 217811 -80
rect 217839 -108 226625 -80
rect 226653 -108 226687 -80
rect 226715 -108 226749 -80
rect 226777 -108 226811 -80
rect 226839 -108 235625 -80
rect 235653 -108 235687 -80
rect 235715 -108 235749 -80
rect 235777 -108 235811 -80
rect 235839 -108 244625 -80
rect 244653 -108 244687 -80
rect 244715 -108 244749 -80
rect 244777 -108 244811 -80
rect 244839 -108 253625 -80
rect 253653 -108 253687 -80
rect 253715 -108 253749 -80
rect 253777 -108 253811 -80
rect 253839 -108 262625 -80
rect 262653 -108 262687 -80
rect 262715 -108 262749 -80
rect 262777 -108 262811 -80
rect 262839 -108 271625 -80
rect 271653 -108 271687 -80
rect 271715 -108 271749 -80
rect 271777 -108 271811 -80
rect 271839 -108 280625 -80
rect 280653 -108 280687 -80
rect 280715 -108 280749 -80
rect 280777 -108 280811 -80
rect 280839 -108 289625 -80
rect 289653 -108 289687 -80
rect 289715 -108 289749 -80
rect 289777 -108 289811 -80
rect 289839 -108 298248 -80
rect 298276 -108 298310 -80
rect 298338 -108 298372 -80
rect 298400 -108 298434 -80
rect 298462 -108 298510 -80
rect -478 -142 298510 -108
rect -478 -170 -430 -142
rect -402 -170 -368 -142
rect -340 -170 -306 -142
rect -278 -170 -244 -142
rect -216 -170 1625 -142
rect 1653 -170 1687 -142
rect 1715 -170 1749 -142
rect 1777 -170 1811 -142
rect 1839 -170 10625 -142
rect 10653 -170 10687 -142
rect 10715 -170 10749 -142
rect 10777 -170 10811 -142
rect 10839 -170 19625 -142
rect 19653 -170 19687 -142
rect 19715 -170 19749 -142
rect 19777 -170 19811 -142
rect 19839 -170 28625 -142
rect 28653 -170 28687 -142
rect 28715 -170 28749 -142
rect 28777 -170 28811 -142
rect 28839 -170 37625 -142
rect 37653 -170 37687 -142
rect 37715 -170 37749 -142
rect 37777 -170 37811 -142
rect 37839 -170 46625 -142
rect 46653 -170 46687 -142
rect 46715 -170 46749 -142
rect 46777 -170 46811 -142
rect 46839 -170 55625 -142
rect 55653 -170 55687 -142
rect 55715 -170 55749 -142
rect 55777 -170 55811 -142
rect 55839 -170 64625 -142
rect 64653 -170 64687 -142
rect 64715 -170 64749 -142
rect 64777 -170 64811 -142
rect 64839 -170 73625 -142
rect 73653 -170 73687 -142
rect 73715 -170 73749 -142
rect 73777 -170 73811 -142
rect 73839 -170 82625 -142
rect 82653 -170 82687 -142
rect 82715 -170 82749 -142
rect 82777 -170 82811 -142
rect 82839 -170 91625 -142
rect 91653 -170 91687 -142
rect 91715 -170 91749 -142
rect 91777 -170 91811 -142
rect 91839 -170 100625 -142
rect 100653 -170 100687 -142
rect 100715 -170 100749 -142
rect 100777 -170 100811 -142
rect 100839 -170 109625 -142
rect 109653 -170 109687 -142
rect 109715 -170 109749 -142
rect 109777 -170 109811 -142
rect 109839 -170 118625 -142
rect 118653 -170 118687 -142
rect 118715 -170 118749 -142
rect 118777 -170 118811 -142
rect 118839 -170 127625 -142
rect 127653 -170 127687 -142
rect 127715 -170 127749 -142
rect 127777 -170 127811 -142
rect 127839 -170 136625 -142
rect 136653 -170 136687 -142
rect 136715 -170 136749 -142
rect 136777 -170 136811 -142
rect 136839 -170 145625 -142
rect 145653 -170 145687 -142
rect 145715 -170 145749 -142
rect 145777 -170 145811 -142
rect 145839 -170 154625 -142
rect 154653 -170 154687 -142
rect 154715 -170 154749 -142
rect 154777 -170 154811 -142
rect 154839 -170 163625 -142
rect 163653 -170 163687 -142
rect 163715 -170 163749 -142
rect 163777 -170 163811 -142
rect 163839 -170 172625 -142
rect 172653 -170 172687 -142
rect 172715 -170 172749 -142
rect 172777 -170 172811 -142
rect 172839 -170 181625 -142
rect 181653 -170 181687 -142
rect 181715 -170 181749 -142
rect 181777 -170 181811 -142
rect 181839 -170 190625 -142
rect 190653 -170 190687 -142
rect 190715 -170 190749 -142
rect 190777 -170 190811 -142
rect 190839 -170 199625 -142
rect 199653 -170 199687 -142
rect 199715 -170 199749 -142
rect 199777 -170 199811 -142
rect 199839 -170 208625 -142
rect 208653 -170 208687 -142
rect 208715 -170 208749 -142
rect 208777 -170 208811 -142
rect 208839 -170 217625 -142
rect 217653 -170 217687 -142
rect 217715 -170 217749 -142
rect 217777 -170 217811 -142
rect 217839 -170 226625 -142
rect 226653 -170 226687 -142
rect 226715 -170 226749 -142
rect 226777 -170 226811 -142
rect 226839 -170 235625 -142
rect 235653 -170 235687 -142
rect 235715 -170 235749 -142
rect 235777 -170 235811 -142
rect 235839 -170 244625 -142
rect 244653 -170 244687 -142
rect 244715 -170 244749 -142
rect 244777 -170 244811 -142
rect 244839 -170 253625 -142
rect 253653 -170 253687 -142
rect 253715 -170 253749 -142
rect 253777 -170 253811 -142
rect 253839 -170 262625 -142
rect 262653 -170 262687 -142
rect 262715 -170 262749 -142
rect 262777 -170 262811 -142
rect 262839 -170 271625 -142
rect 271653 -170 271687 -142
rect 271715 -170 271749 -142
rect 271777 -170 271811 -142
rect 271839 -170 280625 -142
rect 280653 -170 280687 -142
rect 280715 -170 280749 -142
rect 280777 -170 280811 -142
rect 280839 -170 289625 -142
rect 289653 -170 289687 -142
rect 289715 -170 289749 -142
rect 289777 -170 289811 -142
rect 289839 -170 298248 -142
rect 298276 -170 298310 -142
rect 298338 -170 298372 -142
rect 298400 -170 298434 -142
rect 298462 -170 298510 -142
rect -478 -204 298510 -170
rect -478 -232 -430 -204
rect -402 -232 -368 -204
rect -340 -232 -306 -204
rect -278 -232 -244 -204
rect -216 -232 1625 -204
rect 1653 -232 1687 -204
rect 1715 -232 1749 -204
rect 1777 -232 1811 -204
rect 1839 -232 10625 -204
rect 10653 -232 10687 -204
rect 10715 -232 10749 -204
rect 10777 -232 10811 -204
rect 10839 -232 19625 -204
rect 19653 -232 19687 -204
rect 19715 -232 19749 -204
rect 19777 -232 19811 -204
rect 19839 -232 28625 -204
rect 28653 -232 28687 -204
rect 28715 -232 28749 -204
rect 28777 -232 28811 -204
rect 28839 -232 37625 -204
rect 37653 -232 37687 -204
rect 37715 -232 37749 -204
rect 37777 -232 37811 -204
rect 37839 -232 46625 -204
rect 46653 -232 46687 -204
rect 46715 -232 46749 -204
rect 46777 -232 46811 -204
rect 46839 -232 55625 -204
rect 55653 -232 55687 -204
rect 55715 -232 55749 -204
rect 55777 -232 55811 -204
rect 55839 -232 64625 -204
rect 64653 -232 64687 -204
rect 64715 -232 64749 -204
rect 64777 -232 64811 -204
rect 64839 -232 73625 -204
rect 73653 -232 73687 -204
rect 73715 -232 73749 -204
rect 73777 -232 73811 -204
rect 73839 -232 82625 -204
rect 82653 -232 82687 -204
rect 82715 -232 82749 -204
rect 82777 -232 82811 -204
rect 82839 -232 91625 -204
rect 91653 -232 91687 -204
rect 91715 -232 91749 -204
rect 91777 -232 91811 -204
rect 91839 -232 100625 -204
rect 100653 -232 100687 -204
rect 100715 -232 100749 -204
rect 100777 -232 100811 -204
rect 100839 -232 109625 -204
rect 109653 -232 109687 -204
rect 109715 -232 109749 -204
rect 109777 -232 109811 -204
rect 109839 -232 118625 -204
rect 118653 -232 118687 -204
rect 118715 -232 118749 -204
rect 118777 -232 118811 -204
rect 118839 -232 127625 -204
rect 127653 -232 127687 -204
rect 127715 -232 127749 -204
rect 127777 -232 127811 -204
rect 127839 -232 136625 -204
rect 136653 -232 136687 -204
rect 136715 -232 136749 -204
rect 136777 -232 136811 -204
rect 136839 -232 145625 -204
rect 145653 -232 145687 -204
rect 145715 -232 145749 -204
rect 145777 -232 145811 -204
rect 145839 -232 154625 -204
rect 154653 -232 154687 -204
rect 154715 -232 154749 -204
rect 154777 -232 154811 -204
rect 154839 -232 163625 -204
rect 163653 -232 163687 -204
rect 163715 -232 163749 -204
rect 163777 -232 163811 -204
rect 163839 -232 172625 -204
rect 172653 -232 172687 -204
rect 172715 -232 172749 -204
rect 172777 -232 172811 -204
rect 172839 -232 181625 -204
rect 181653 -232 181687 -204
rect 181715 -232 181749 -204
rect 181777 -232 181811 -204
rect 181839 -232 190625 -204
rect 190653 -232 190687 -204
rect 190715 -232 190749 -204
rect 190777 -232 190811 -204
rect 190839 -232 199625 -204
rect 199653 -232 199687 -204
rect 199715 -232 199749 -204
rect 199777 -232 199811 -204
rect 199839 -232 208625 -204
rect 208653 -232 208687 -204
rect 208715 -232 208749 -204
rect 208777 -232 208811 -204
rect 208839 -232 217625 -204
rect 217653 -232 217687 -204
rect 217715 -232 217749 -204
rect 217777 -232 217811 -204
rect 217839 -232 226625 -204
rect 226653 -232 226687 -204
rect 226715 -232 226749 -204
rect 226777 -232 226811 -204
rect 226839 -232 235625 -204
rect 235653 -232 235687 -204
rect 235715 -232 235749 -204
rect 235777 -232 235811 -204
rect 235839 -232 244625 -204
rect 244653 -232 244687 -204
rect 244715 -232 244749 -204
rect 244777 -232 244811 -204
rect 244839 -232 253625 -204
rect 253653 -232 253687 -204
rect 253715 -232 253749 -204
rect 253777 -232 253811 -204
rect 253839 -232 262625 -204
rect 262653 -232 262687 -204
rect 262715 -232 262749 -204
rect 262777 -232 262811 -204
rect 262839 -232 271625 -204
rect 271653 -232 271687 -204
rect 271715 -232 271749 -204
rect 271777 -232 271811 -204
rect 271839 -232 280625 -204
rect 280653 -232 280687 -204
rect 280715 -232 280749 -204
rect 280777 -232 280811 -204
rect 280839 -232 289625 -204
rect 289653 -232 289687 -204
rect 289715 -232 289749 -204
rect 289777 -232 289811 -204
rect 289839 -232 298248 -204
rect 298276 -232 298310 -204
rect 298338 -232 298372 -204
rect 298400 -232 298434 -204
rect 298462 -232 298510 -204
rect -478 -266 298510 -232
rect -478 -294 -430 -266
rect -402 -294 -368 -266
rect -340 -294 -306 -266
rect -278 -294 -244 -266
rect -216 -294 1625 -266
rect 1653 -294 1687 -266
rect 1715 -294 1749 -266
rect 1777 -294 1811 -266
rect 1839 -294 10625 -266
rect 10653 -294 10687 -266
rect 10715 -294 10749 -266
rect 10777 -294 10811 -266
rect 10839 -294 19625 -266
rect 19653 -294 19687 -266
rect 19715 -294 19749 -266
rect 19777 -294 19811 -266
rect 19839 -294 28625 -266
rect 28653 -294 28687 -266
rect 28715 -294 28749 -266
rect 28777 -294 28811 -266
rect 28839 -294 37625 -266
rect 37653 -294 37687 -266
rect 37715 -294 37749 -266
rect 37777 -294 37811 -266
rect 37839 -294 46625 -266
rect 46653 -294 46687 -266
rect 46715 -294 46749 -266
rect 46777 -294 46811 -266
rect 46839 -294 55625 -266
rect 55653 -294 55687 -266
rect 55715 -294 55749 -266
rect 55777 -294 55811 -266
rect 55839 -294 64625 -266
rect 64653 -294 64687 -266
rect 64715 -294 64749 -266
rect 64777 -294 64811 -266
rect 64839 -294 73625 -266
rect 73653 -294 73687 -266
rect 73715 -294 73749 -266
rect 73777 -294 73811 -266
rect 73839 -294 82625 -266
rect 82653 -294 82687 -266
rect 82715 -294 82749 -266
rect 82777 -294 82811 -266
rect 82839 -294 91625 -266
rect 91653 -294 91687 -266
rect 91715 -294 91749 -266
rect 91777 -294 91811 -266
rect 91839 -294 100625 -266
rect 100653 -294 100687 -266
rect 100715 -294 100749 -266
rect 100777 -294 100811 -266
rect 100839 -294 109625 -266
rect 109653 -294 109687 -266
rect 109715 -294 109749 -266
rect 109777 -294 109811 -266
rect 109839 -294 118625 -266
rect 118653 -294 118687 -266
rect 118715 -294 118749 -266
rect 118777 -294 118811 -266
rect 118839 -294 127625 -266
rect 127653 -294 127687 -266
rect 127715 -294 127749 -266
rect 127777 -294 127811 -266
rect 127839 -294 136625 -266
rect 136653 -294 136687 -266
rect 136715 -294 136749 -266
rect 136777 -294 136811 -266
rect 136839 -294 145625 -266
rect 145653 -294 145687 -266
rect 145715 -294 145749 -266
rect 145777 -294 145811 -266
rect 145839 -294 154625 -266
rect 154653 -294 154687 -266
rect 154715 -294 154749 -266
rect 154777 -294 154811 -266
rect 154839 -294 163625 -266
rect 163653 -294 163687 -266
rect 163715 -294 163749 -266
rect 163777 -294 163811 -266
rect 163839 -294 172625 -266
rect 172653 -294 172687 -266
rect 172715 -294 172749 -266
rect 172777 -294 172811 -266
rect 172839 -294 181625 -266
rect 181653 -294 181687 -266
rect 181715 -294 181749 -266
rect 181777 -294 181811 -266
rect 181839 -294 190625 -266
rect 190653 -294 190687 -266
rect 190715 -294 190749 -266
rect 190777 -294 190811 -266
rect 190839 -294 199625 -266
rect 199653 -294 199687 -266
rect 199715 -294 199749 -266
rect 199777 -294 199811 -266
rect 199839 -294 208625 -266
rect 208653 -294 208687 -266
rect 208715 -294 208749 -266
rect 208777 -294 208811 -266
rect 208839 -294 217625 -266
rect 217653 -294 217687 -266
rect 217715 -294 217749 -266
rect 217777 -294 217811 -266
rect 217839 -294 226625 -266
rect 226653 -294 226687 -266
rect 226715 -294 226749 -266
rect 226777 -294 226811 -266
rect 226839 -294 235625 -266
rect 235653 -294 235687 -266
rect 235715 -294 235749 -266
rect 235777 -294 235811 -266
rect 235839 -294 244625 -266
rect 244653 -294 244687 -266
rect 244715 -294 244749 -266
rect 244777 -294 244811 -266
rect 244839 -294 253625 -266
rect 253653 -294 253687 -266
rect 253715 -294 253749 -266
rect 253777 -294 253811 -266
rect 253839 -294 262625 -266
rect 262653 -294 262687 -266
rect 262715 -294 262749 -266
rect 262777 -294 262811 -266
rect 262839 -294 271625 -266
rect 271653 -294 271687 -266
rect 271715 -294 271749 -266
rect 271777 -294 271811 -266
rect 271839 -294 280625 -266
rect 280653 -294 280687 -266
rect 280715 -294 280749 -266
rect 280777 -294 280811 -266
rect 280839 -294 289625 -266
rect 289653 -294 289687 -266
rect 289715 -294 289749 -266
rect 289777 -294 289811 -266
rect 289839 -294 298248 -266
rect 298276 -294 298310 -266
rect 298338 -294 298372 -266
rect 298400 -294 298434 -266
rect 298462 -294 298510 -266
rect -478 -342 298510 -294
rect -958 -560 298990 -512
rect -958 -588 -910 -560
rect -882 -588 -848 -560
rect -820 -588 -786 -560
rect -758 -588 -724 -560
rect -696 -588 3485 -560
rect 3513 -588 3547 -560
rect 3575 -588 3609 -560
rect 3637 -588 3671 -560
rect 3699 -588 12485 -560
rect 12513 -588 12547 -560
rect 12575 -588 12609 -560
rect 12637 -588 12671 -560
rect 12699 -588 21485 -560
rect 21513 -588 21547 -560
rect 21575 -588 21609 -560
rect 21637 -588 21671 -560
rect 21699 -588 30485 -560
rect 30513 -588 30547 -560
rect 30575 -588 30609 -560
rect 30637 -588 30671 -560
rect 30699 -588 39485 -560
rect 39513 -588 39547 -560
rect 39575 -588 39609 -560
rect 39637 -588 39671 -560
rect 39699 -588 48485 -560
rect 48513 -588 48547 -560
rect 48575 -588 48609 -560
rect 48637 -588 48671 -560
rect 48699 -588 57485 -560
rect 57513 -588 57547 -560
rect 57575 -588 57609 -560
rect 57637 -588 57671 -560
rect 57699 -588 66485 -560
rect 66513 -588 66547 -560
rect 66575 -588 66609 -560
rect 66637 -588 66671 -560
rect 66699 -588 75485 -560
rect 75513 -588 75547 -560
rect 75575 -588 75609 -560
rect 75637 -588 75671 -560
rect 75699 -588 84485 -560
rect 84513 -588 84547 -560
rect 84575 -588 84609 -560
rect 84637 -588 84671 -560
rect 84699 -588 93485 -560
rect 93513 -588 93547 -560
rect 93575 -588 93609 -560
rect 93637 -588 93671 -560
rect 93699 -588 102485 -560
rect 102513 -588 102547 -560
rect 102575 -588 102609 -560
rect 102637 -588 102671 -560
rect 102699 -588 111485 -560
rect 111513 -588 111547 -560
rect 111575 -588 111609 -560
rect 111637 -588 111671 -560
rect 111699 -588 120485 -560
rect 120513 -588 120547 -560
rect 120575 -588 120609 -560
rect 120637 -588 120671 -560
rect 120699 -588 129485 -560
rect 129513 -588 129547 -560
rect 129575 -588 129609 -560
rect 129637 -588 129671 -560
rect 129699 -588 138485 -560
rect 138513 -588 138547 -560
rect 138575 -588 138609 -560
rect 138637 -588 138671 -560
rect 138699 -588 147485 -560
rect 147513 -588 147547 -560
rect 147575 -588 147609 -560
rect 147637 -588 147671 -560
rect 147699 -588 156485 -560
rect 156513 -588 156547 -560
rect 156575 -588 156609 -560
rect 156637 -588 156671 -560
rect 156699 -588 165485 -560
rect 165513 -588 165547 -560
rect 165575 -588 165609 -560
rect 165637 -588 165671 -560
rect 165699 -588 174485 -560
rect 174513 -588 174547 -560
rect 174575 -588 174609 -560
rect 174637 -588 174671 -560
rect 174699 -588 183485 -560
rect 183513 -588 183547 -560
rect 183575 -588 183609 -560
rect 183637 -588 183671 -560
rect 183699 -588 192485 -560
rect 192513 -588 192547 -560
rect 192575 -588 192609 -560
rect 192637 -588 192671 -560
rect 192699 -588 201485 -560
rect 201513 -588 201547 -560
rect 201575 -588 201609 -560
rect 201637 -588 201671 -560
rect 201699 -588 210485 -560
rect 210513 -588 210547 -560
rect 210575 -588 210609 -560
rect 210637 -588 210671 -560
rect 210699 -588 219485 -560
rect 219513 -588 219547 -560
rect 219575 -588 219609 -560
rect 219637 -588 219671 -560
rect 219699 -588 228485 -560
rect 228513 -588 228547 -560
rect 228575 -588 228609 -560
rect 228637 -588 228671 -560
rect 228699 -588 237485 -560
rect 237513 -588 237547 -560
rect 237575 -588 237609 -560
rect 237637 -588 237671 -560
rect 237699 -588 246485 -560
rect 246513 -588 246547 -560
rect 246575 -588 246609 -560
rect 246637 -588 246671 -560
rect 246699 -588 255485 -560
rect 255513 -588 255547 -560
rect 255575 -588 255609 -560
rect 255637 -588 255671 -560
rect 255699 -588 264485 -560
rect 264513 -588 264547 -560
rect 264575 -588 264609 -560
rect 264637 -588 264671 -560
rect 264699 -588 273485 -560
rect 273513 -588 273547 -560
rect 273575 -588 273609 -560
rect 273637 -588 273671 -560
rect 273699 -588 282485 -560
rect 282513 -588 282547 -560
rect 282575 -588 282609 -560
rect 282637 -588 282671 -560
rect 282699 -588 291485 -560
rect 291513 -588 291547 -560
rect 291575 -588 291609 -560
rect 291637 -588 291671 -560
rect 291699 -588 298728 -560
rect 298756 -588 298790 -560
rect 298818 -588 298852 -560
rect 298880 -588 298914 -560
rect 298942 -588 298990 -560
rect -958 -622 298990 -588
rect -958 -650 -910 -622
rect -882 -650 -848 -622
rect -820 -650 -786 -622
rect -758 -650 -724 -622
rect -696 -650 3485 -622
rect 3513 -650 3547 -622
rect 3575 -650 3609 -622
rect 3637 -650 3671 -622
rect 3699 -650 12485 -622
rect 12513 -650 12547 -622
rect 12575 -650 12609 -622
rect 12637 -650 12671 -622
rect 12699 -650 21485 -622
rect 21513 -650 21547 -622
rect 21575 -650 21609 -622
rect 21637 -650 21671 -622
rect 21699 -650 30485 -622
rect 30513 -650 30547 -622
rect 30575 -650 30609 -622
rect 30637 -650 30671 -622
rect 30699 -650 39485 -622
rect 39513 -650 39547 -622
rect 39575 -650 39609 -622
rect 39637 -650 39671 -622
rect 39699 -650 48485 -622
rect 48513 -650 48547 -622
rect 48575 -650 48609 -622
rect 48637 -650 48671 -622
rect 48699 -650 57485 -622
rect 57513 -650 57547 -622
rect 57575 -650 57609 -622
rect 57637 -650 57671 -622
rect 57699 -650 66485 -622
rect 66513 -650 66547 -622
rect 66575 -650 66609 -622
rect 66637 -650 66671 -622
rect 66699 -650 75485 -622
rect 75513 -650 75547 -622
rect 75575 -650 75609 -622
rect 75637 -650 75671 -622
rect 75699 -650 84485 -622
rect 84513 -650 84547 -622
rect 84575 -650 84609 -622
rect 84637 -650 84671 -622
rect 84699 -650 93485 -622
rect 93513 -650 93547 -622
rect 93575 -650 93609 -622
rect 93637 -650 93671 -622
rect 93699 -650 102485 -622
rect 102513 -650 102547 -622
rect 102575 -650 102609 -622
rect 102637 -650 102671 -622
rect 102699 -650 111485 -622
rect 111513 -650 111547 -622
rect 111575 -650 111609 -622
rect 111637 -650 111671 -622
rect 111699 -650 120485 -622
rect 120513 -650 120547 -622
rect 120575 -650 120609 -622
rect 120637 -650 120671 -622
rect 120699 -650 129485 -622
rect 129513 -650 129547 -622
rect 129575 -650 129609 -622
rect 129637 -650 129671 -622
rect 129699 -650 138485 -622
rect 138513 -650 138547 -622
rect 138575 -650 138609 -622
rect 138637 -650 138671 -622
rect 138699 -650 147485 -622
rect 147513 -650 147547 -622
rect 147575 -650 147609 -622
rect 147637 -650 147671 -622
rect 147699 -650 156485 -622
rect 156513 -650 156547 -622
rect 156575 -650 156609 -622
rect 156637 -650 156671 -622
rect 156699 -650 165485 -622
rect 165513 -650 165547 -622
rect 165575 -650 165609 -622
rect 165637 -650 165671 -622
rect 165699 -650 174485 -622
rect 174513 -650 174547 -622
rect 174575 -650 174609 -622
rect 174637 -650 174671 -622
rect 174699 -650 183485 -622
rect 183513 -650 183547 -622
rect 183575 -650 183609 -622
rect 183637 -650 183671 -622
rect 183699 -650 192485 -622
rect 192513 -650 192547 -622
rect 192575 -650 192609 -622
rect 192637 -650 192671 -622
rect 192699 -650 201485 -622
rect 201513 -650 201547 -622
rect 201575 -650 201609 -622
rect 201637 -650 201671 -622
rect 201699 -650 210485 -622
rect 210513 -650 210547 -622
rect 210575 -650 210609 -622
rect 210637 -650 210671 -622
rect 210699 -650 219485 -622
rect 219513 -650 219547 -622
rect 219575 -650 219609 -622
rect 219637 -650 219671 -622
rect 219699 -650 228485 -622
rect 228513 -650 228547 -622
rect 228575 -650 228609 -622
rect 228637 -650 228671 -622
rect 228699 -650 237485 -622
rect 237513 -650 237547 -622
rect 237575 -650 237609 -622
rect 237637 -650 237671 -622
rect 237699 -650 246485 -622
rect 246513 -650 246547 -622
rect 246575 -650 246609 -622
rect 246637 -650 246671 -622
rect 246699 -650 255485 -622
rect 255513 -650 255547 -622
rect 255575 -650 255609 -622
rect 255637 -650 255671 -622
rect 255699 -650 264485 -622
rect 264513 -650 264547 -622
rect 264575 -650 264609 -622
rect 264637 -650 264671 -622
rect 264699 -650 273485 -622
rect 273513 -650 273547 -622
rect 273575 -650 273609 -622
rect 273637 -650 273671 -622
rect 273699 -650 282485 -622
rect 282513 -650 282547 -622
rect 282575 -650 282609 -622
rect 282637 -650 282671 -622
rect 282699 -650 291485 -622
rect 291513 -650 291547 -622
rect 291575 -650 291609 -622
rect 291637 -650 291671 -622
rect 291699 -650 298728 -622
rect 298756 -650 298790 -622
rect 298818 -650 298852 -622
rect 298880 -650 298914 -622
rect 298942 -650 298990 -622
rect -958 -684 298990 -650
rect -958 -712 -910 -684
rect -882 -712 -848 -684
rect -820 -712 -786 -684
rect -758 -712 -724 -684
rect -696 -712 3485 -684
rect 3513 -712 3547 -684
rect 3575 -712 3609 -684
rect 3637 -712 3671 -684
rect 3699 -712 12485 -684
rect 12513 -712 12547 -684
rect 12575 -712 12609 -684
rect 12637 -712 12671 -684
rect 12699 -712 21485 -684
rect 21513 -712 21547 -684
rect 21575 -712 21609 -684
rect 21637 -712 21671 -684
rect 21699 -712 30485 -684
rect 30513 -712 30547 -684
rect 30575 -712 30609 -684
rect 30637 -712 30671 -684
rect 30699 -712 39485 -684
rect 39513 -712 39547 -684
rect 39575 -712 39609 -684
rect 39637 -712 39671 -684
rect 39699 -712 48485 -684
rect 48513 -712 48547 -684
rect 48575 -712 48609 -684
rect 48637 -712 48671 -684
rect 48699 -712 57485 -684
rect 57513 -712 57547 -684
rect 57575 -712 57609 -684
rect 57637 -712 57671 -684
rect 57699 -712 66485 -684
rect 66513 -712 66547 -684
rect 66575 -712 66609 -684
rect 66637 -712 66671 -684
rect 66699 -712 75485 -684
rect 75513 -712 75547 -684
rect 75575 -712 75609 -684
rect 75637 -712 75671 -684
rect 75699 -712 84485 -684
rect 84513 -712 84547 -684
rect 84575 -712 84609 -684
rect 84637 -712 84671 -684
rect 84699 -712 93485 -684
rect 93513 -712 93547 -684
rect 93575 -712 93609 -684
rect 93637 -712 93671 -684
rect 93699 -712 102485 -684
rect 102513 -712 102547 -684
rect 102575 -712 102609 -684
rect 102637 -712 102671 -684
rect 102699 -712 111485 -684
rect 111513 -712 111547 -684
rect 111575 -712 111609 -684
rect 111637 -712 111671 -684
rect 111699 -712 120485 -684
rect 120513 -712 120547 -684
rect 120575 -712 120609 -684
rect 120637 -712 120671 -684
rect 120699 -712 129485 -684
rect 129513 -712 129547 -684
rect 129575 -712 129609 -684
rect 129637 -712 129671 -684
rect 129699 -712 138485 -684
rect 138513 -712 138547 -684
rect 138575 -712 138609 -684
rect 138637 -712 138671 -684
rect 138699 -712 147485 -684
rect 147513 -712 147547 -684
rect 147575 -712 147609 -684
rect 147637 -712 147671 -684
rect 147699 -712 156485 -684
rect 156513 -712 156547 -684
rect 156575 -712 156609 -684
rect 156637 -712 156671 -684
rect 156699 -712 165485 -684
rect 165513 -712 165547 -684
rect 165575 -712 165609 -684
rect 165637 -712 165671 -684
rect 165699 -712 174485 -684
rect 174513 -712 174547 -684
rect 174575 -712 174609 -684
rect 174637 -712 174671 -684
rect 174699 -712 183485 -684
rect 183513 -712 183547 -684
rect 183575 -712 183609 -684
rect 183637 -712 183671 -684
rect 183699 -712 192485 -684
rect 192513 -712 192547 -684
rect 192575 -712 192609 -684
rect 192637 -712 192671 -684
rect 192699 -712 201485 -684
rect 201513 -712 201547 -684
rect 201575 -712 201609 -684
rect 201637 -712 201671 -684
rect 201699 -712 210485 -684
rect 210513 -712 210547 -684
rect 210575 -712 210609 -684
rect 210637 -712 210671 -684
rect 210699 -712 219485 -684
rect 219513 -712 219547 -684
rect 219575 -712 219609 -684
rect 219637 -712 219671 -684
rect 219699 -712 228485 -684
rect 228513 -712 228547 -684
rect 228575 -712 228609 -684
rect 228637 -712 228671 -684
rect 228699 -712 237485 -684
rect 237513 -712 237547 -684
rect 237575 -712 237609 -684
rect 237637 -712 237671 -684
rect 237699 -712 246485 -684
rect 246513 -712 246547 -684
rect 246575 -712 246609 -684
rect 246637 -712 246671 -684
rect 246699 -712 255485 -684
rect 255513 -712 255547 -684
rect 255575 -712 255609 -684
rect 255637 -712 255671 -684
rect 255699 -712 264485 -684
rect 264513 -712 264547 -684
rect 264575 -712 264609 -684
rect 264637 -712 264671 -684
rect 264699 -712 273485 -684
rect 273513 -712 273547 -684
rect 273575 -712 273609 -684
rect 273637 -712 273671 -684
rect 273699 -712 282485 -684
rect 282513 -712 282547 -684
rect 282575 -712 282609 -684
rect 282637 -712 282671 -684
rect 282699 -712 291485 -684
rect 291513 -712 291547 -684
rect 291575 -712 291609 -684
rect 291637 -712 291671 -684
rect 291699 -712 298728 -684
rect 298756 -712 298790 -684
rect 298818 -712 298852 -684
rect 298880 -712 298914 -684
rect 298942 -712 298990 -684
rect -958 -746 298990 -712
rect -958 -774 -910 -746
rect -882 -774 -848 -746
rect -820 -774 -786 -746
rect -758 -774 -724 -746
rect -696 -774 3485 -746
rect 3513 -774 3547 -746
rect 3575 -774 3609 -746
rect 3637 -774 3671 -746
rect 3699 -774 12485 -746
rect 12513 -774 12547 -746
rect 12575 -774 12609 -746
rect 12637 -774 12671 -746
rect 12699 -774 21485 -746
rect 21513 -774 21547 -746
rect 21575 -774 21609 -746
rect 21637 -774 21671 -746
rect 21699 -774 30485 -746
rect 30513 -774 30547 -746
rect 30575 -774 30609 -746
rect 30637 -774 30671 -746
rect 30699 -774 39485 -746
rect 39513 -774 39547 -746
rect 39575 -774 39609 -746
rect 39637 -774 39671 -746
rect 39699 -774 48485 -746
rect 48513 -774 48547 -746
rect 48575 -774 48609 -746
rect 48637 -774 48671 -746
rect 48699 -774 57485 -746
rect 57513 -774 57547 -746
rect 57575 -774 57609 -746
rect 57637 -774 57671 -746
rect 57699 -774 66485 -746
rect 66513 -774 66547 -746
rect 66575 -774 66609 -746
rect 66637 -774 66671 -746
rect 66699 -774 75485 -746
rect 75513 -774 75547 -746
rect 75575 -774 75609 -746
rect 75637 -774 75671 -746
rect 75699 -774 84485 -746
rect 84513 -774 84547 -746
rect 84575 -774 84609 -746
rect 84637 -774 84671 -746
rect 84699 -774 93485 -746
rect 93513 -774 93547 -746
rect 93575 -774 93609 -746
rect 93637 -774 93671 -746
rect 93699 -774 102485 -746
rect 102513 -774 102547 -746
rect 102575 -774 102609 -746
rect 102637 -774 102671 -746
rect 102699 -774 111485 -746
rect 111513 -774 111547 -746
rect 111575 -774 111609 -746
rect 111637 -774 111671 -746
rect 111699 -774 120485 -746
rect 120513 -774 120547 -746
rect 120575 -774 120609 -746
rect 120637 -774 120671 -746
rect 120699 -774 129485 -746
rect 129513 -774 129547 -746
rect 129575 -774 129609 -746
rect 129637 -774 129671 -746
rect 129699 -774 138485 -746
rect 138513 -774 138547 -746
rect 138575 -774 138609 -746
rect 138637 -774 138671 -746
rect 138699 -774 147485 -746
rect 147513 -774 147547 -746
rect 147575 -774 147609 -746
rect 147637 -774 147671 -746
rect 147699 -774 156485 -746
rect 156513 -774 156547 -746
rect 156575 -774 156609 -746
rect 156637 -774 156671 -746
rect 156699 -774 165485 -746
rect 165513 -774 165547 -746
rect 165575 -774 165609 -746
rect 165637 -774 165671 -746
rect 165699 -774 174485 -746
rect 174513 -774 174547 -746
rect 174575 -774 174609 -746
rect 174637 -774 174671 -746
rect 174699 -774 183485 -746
rect 183513 -774 183547 -746
rect 183575 -774 183609 -746
rect 183637 -774 183671 -746
rect 183699 -774 192485 -746
rect 192513 -774 192547 -746
rect 192575 -774 192609 -746
rect 192637 -774 192671 -746
rect 192699 -774 201485 -746
rect 201513 -774 201547 -746
rect 201575 -774 201609 -746
rect 201637 -774 201671 -746
rect 201699 -774 210485 -746
rect 210513 -774 210547 -746
rect 210575 -774 210609 -746
rect 210637 -774 210671 -746
rect 210699 -774 219485 -746
rect 219513 -774 219547 -746
rect 219575 -774 219609 -746
rect 219637 -774 219671 -746
rect 219699 -774 228485 -746
rect 228513 -774 228547 -746
rect 228575 -774 228609 -746
rect 228637 -774 228671 -746
rect 228699 -774 237485 -746
rect 237513 -774 237547 -746
rect 237575 -774 237609 -746
rect 237637 -774 237671 -746
rect 237699 -774 246485 -746
rect 246513 -774 246547 -746
rect 246575 -774 246609 -746
rect 246637 -774 246671 -746
rect 246699 -774 255485 -746
rect 255513 -774 255547 -746
rect 255575 -774 255609 -746
rect 255637 -774 255671 -746
rect 255699 -774 264485 -746
rect 264513 -774 264547 -746
rect 264575 -774 264609 -746
rect 264637 -774 264671 -746
rect 264699 -774 273485 -746
rect 273513 -774 273547 -746
rect 273575 -774 273609 -746
rect 273637 -774 273671 -746
rect 273699 -774 282485 -746
rect 282513 -774 282547 -746
rect 282575 -774 282609 -746
rect 282637 -774 282671 -746
rect 282699 -774 291485 -746
rect 291513 -774 291547 -746
rect 291575 -774 291609 -746
rect 291637 -774 291671 -746
rect 291699 -774 298728 -746
rect 298756 -774 298790 -746
rect 298818 -774 298852 -746
rect 298880 -774 298914 -746
rect 298942 -774 298990 -746
rect -958 -822 298990 -774
use serv_0  u_serv_0
timestamp 0
transform 1 0 50000 0 1 50000
box 672 345 70000 58438
use serv_1  u_serv_1
timestamp 0
transform 1 0 50000 0 1 125000
box 672 233 100000 58438
use serv_2  u_serv_2
timestamp 0
transform 1 0 50000 0 1 200000
box 672 233 100000 59575
<< labels >>
flabel metal3 s 297780 3556 298500 3668 0 FreeSans 448 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 297780 201796 298500 201908 0 FreeSans 448 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 297780 221620 298500 221732 0 FreeSans 448 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 297780 241444 298500 241556 0 FreeSans 448 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 297780 261268 298500 261380 0 FreeSans 448 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 297780 281092 298500 281204 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 292348 297780 292460 298500 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 259252 297780 259364 298500 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 226156 297780 226268 298500 0 FreeSans 448 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 193060 297780 193172 298500 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 159964 297780 160076 298500 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 297780 23380 298500 23492 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 126868 297780 126980 298500 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 93772 297780 93884 298500 0 FreeSans 448 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 60676 297780 60788 298500 0 FreeSans 448 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 27580 297780 27692 298500 0 FreeSans 448 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -480 293580 240 293692 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -480 272412 240 272524 0 FreeSans 448 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -480 251244 240 251356 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -480 230076 240 230188 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -480 208908 240 209020 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -480 187740 240 187852 0 FreeSans 448 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 297780 43204 298500 43316 0 FreeSans 448 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -480 166572 240 166684 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -480 145404 240 145516 0 FreeSans 448 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -480 124236 240 124348 0 FreeSans 448 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -480 103068 240 103180 0 FreeSans 448 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -480 81900 240 82012 0 FreeSans 448 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -480 60732 240 60844 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -480 39564 240 39676 0 FreeSans 448 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -480 18396 240 18508 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 297780 63028 298500 63140 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 297780 82852 298500 82964 0 FreeSans 448 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 297780 102676 298500 102788 0 FreeSans 448 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 297780 122500 298500 122612 0 FreeSans 448 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 297780 142324 298500 142436 0 FreeSans 448 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 297780 162148 298500 162260 0 FreeSans 448 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 297780 181972 298500 182084 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 297780 16772 298500 16884 0 FreeSans 448 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 297780 215012 298500 215124 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 297780 234836 298500 234948 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 297780 254660 298500 254772 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 297780 274484 298500 274596 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 297780 294308 298500 294420 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 270284 297780 270396 298500 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 237188 297780 237300 298500 0 FreeSans 448 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 204092 297780 204204 298500 0 FreeSans 448 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 170996 297780 171108 298500 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 137900 297780 138012 298500 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 297780 36596 298500 36708 0 FreeSans 448 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 104804 297780 104916 298500 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 71708 297780 71820 298500 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 38612 297780 38724 298500 0 FreeSans 448 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 5516 297780 5628 298500 0 FreeSans 448 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -480 279468 240 279580 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -480 258300 240 258412 0 FreeSans 448 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -480 237132 240 237244 0 FreeSans 448 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -480 215964 240 216076 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -480 194796 240 194908 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -480 173628 240 173740 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 297780 56420 298500 56532 0 FreeSans 448 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -480 152460 240 152572 0 FreeSans 448 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -480 131292 240 131404 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -480 110124 240 110236 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -480 88956 240 89068 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -480 67788 240 67900 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -480 46620 240 46732 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -480 25452 240 25564 0 FreeSans 448 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -480 4284 240 4396 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 297780 76244 298500 76356 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 297780 96068 298500 96180 0 FreeSans 448 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 297780 115892 298500 116004 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 297780 135716 298500 135828 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 297780 155540 298500 155652 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 297780 175364 298500 175476 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 297780 195188 298500 195300 0 FreeSans 448 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 297780 10164 298500 10276 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 297780 208404 298500 208516 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 297780 228228 298500 228340 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 297780 248052 298500 248164 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 297780 267876 298500 267988 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 297780 287700 298500 287812 0 FreeSans 448 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 281316 297780 281428 298500 0 FreeSans 448 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 248220 297780 248332 298500 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 215124 297780 215236 298500 0 FreeSans 448 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 182028 297780 182140 298500 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 148932 297780 149044 298500 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 297780 29988 298500 30100 0 FreeSans 448 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 115836 297780 115948 298500 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 82740 297780 82852 298500 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 49644 297780 49756 298500 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 16548 297780 16660 298500 0 FreeSans 448 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -480 286524 240 286636 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -480 265356 240 265468 0 FreeSans 448 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -480 244188 240 244300 0 FreeSans 448 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -480 223020 240 223132 0 FreeSans 448 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -480 201852 240 201964 0 FreeSans 448 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -480 180684 240 180796 0 FreeSans 448 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 297780 49812 298500 49924 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -480 159516 240 159628 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -480 138348 240 138460 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -480 117180 240 117292 0 FreeSans 448 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -480 96012 240 96124 0 FreeSans 448 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -480 74844 240 74956 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -480 53676 240 53788 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -480 32508 240 32620 0 FreeSans 448 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -480 11340 240 11452 0 FreeSans 448 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 297780 69636 298500 69748 0 FreeSans 448 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 297780 89460 298500 89572 0 FreeSans 448 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 297780 109284 298500 109396 0 FreeSans 448 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 297780 129108 298500 129220 0 FreeSans 448 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 297780 148932 298500 149044 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 297780 168756 298500 168868 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 297780 188580 298500 188692 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 106596 -480 106708 240 0 FreeSans 448 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 135156 -480 135268 240 0 FreeSans 448 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 138012 -480 138124 240 0 FreeSans 448 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 140868 -480 140980 240 0 FreeSans 448 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 143724 -480 143836 240 0 FreeSans 448 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 146580 -480 146692 240 0 FreeSans 448 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 149436 -480 149548 240 0 FreeSans 448 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 152292 -480 152404 240 0 FreeSans 448 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 155148 -480 155260 240 0 FreeSans 448 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 158004 -480 158116 240 0 FreeSans 448 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 160860 -480 160972 240 0 FreeSans 448 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 109452 -480 109564 240 0 FreeSans 448 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 163716 -480 163828 240 0 FreeSans 448 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 166572 -480 166684 240 0 FreeSans 448 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 169428 -480 169540 240 0 FreeSans 448 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 172284 -480 172396 240 0 FreeSans 448 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 175140 -480 175252 240 0 FreeSans 448 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 177996 -480 178108 240 0 FreeSans 448 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 180852 -480 180964 240 0 FreeSans 448 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 183708 -480 183820 240 0 FreeSans 448 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 186564 -480 186676 240 0 FreeSans 448 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 189420 -480 189532 240 0 FreeSans 448 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 112308 -480 112420 240 0 FreeSans 448 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 192276 -480 192388 240 0 FreeSans 448 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 195132 -480 195244 240 0 FreeSans 448 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 197988 -480 198100 240 0 FreeSans 448 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 200844 -480 200956 240 0 FreeSans 448 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 203700 -480 203812 240 0 FreeSans 448 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 206556 -480 206668 240 0 FreeSans 448 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 209412 -480 209524 240 0 FreeSans 448 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 212268 -480 212380 240 0 FreeSans 448 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 215124 -480 215236 240 0 FreeSans 448 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 217980 -480 218092 240 0 FreeSans 448 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 115164 -480 115276 240 0 FreeSans 448 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 220836 -480 220948 240 0 FreeSans 448 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 223692 -480 223804 240 0 FreeSans 448 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 226548 -480 226660 240 0 FreeSans 448 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 229404 -480 229516 240 0 FreeSans 448 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 232260 -480 232372 240 0 FreeSans 448 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 235116 -480 235228 240 0 FreeSans 448 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 237972 -480 238084 240 0 FreeSans 448 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 240828 -480 240940 240 0 FreeSans 448 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 243684 -480 243796 240 0 FreeSans 448 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 246540 -480 246652 240 0 FreeSans 448 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 118020 -480 118132 240 0 FreeSans 448 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 249396 -480 249508 240 0 FreeSans 448 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 252252 -480 252364 240 0 FreeSans 448 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 255108 -480 255220 240 0 FreeSans 448 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 257964 -480 258076 240 0 FreeSans 448 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 260820 -480 260932 240 0 FreeSans 448 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 263676 -480 263788 240 0 FreeSans 448 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 266532 -480 266644 240 0 FreeSans 448 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 269388 -480 269500 240 0 FreeSans 448 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 272244 -480 272356 240 0 FreeSans 448 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 275100 -480 275212 240 0 FreeSans 448 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 120876 -480 120988 240 0 FreeSans 448 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 277956 -480 278068 240 0 FreeSans 448 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 280812 -480 280924 240 0 FreeSans 448 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 283668 -480 283780 240 0 FreeSans 448 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 286524 -480 286636 240 0 FreeSans 448 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 123732 -480 123844 240 0 FreeSans 448 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 126588 -480 126700 240 0 FreeSans 448 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 129444 -480 129556 240 0 FreeSans 448 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 132300 -480 132412 240 0 FreeSans 448 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 107548 -480 107660 240 0 FreeSans 448 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 136108 -480 136220 240 0 FreeSans 448 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 138964 -480 139076 240 0 FreeSans 448 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 141820 -480 141932 240 0 FreeSans 448 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 144676 -480 144788 240 0 FreeSans 448 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 147532 -480 147644 240 0 FreeSans 448 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 150388 -480 150500 240 0 FreeSans 448 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 153244 -480 153356 240 0 FreeSans 448 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 156100 -480 156212 240 0 FreeSans 448 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 158956 -480 159068 240 0 FreeSans 448 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 161812 -480 161924 240 0 FreeSans 448 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 110404 -480 110516 240 0 FreeSans 448 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 164668 -480 164780 240 0 FreeSans 448 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 167524 -480 167636 240 0 FreeSans 448 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 170380 -480 170492 240 0 FreeSans 448 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 173236 -480 173348 240 0 FreeSans 448 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 176092 -480 176204 240 0 FreeSans 448 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 178948 -480 179060 240 0 FreeSans 448 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 181804 -480 181916 240 0 FreeSans 448 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 184660 -480 184772 240 0 FreeSans 448 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 187516 -480 187628 240 0 FreeSans 448 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 190372 -480 190484 240 0 FreeSans 448 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 113260 -480 113372 240 0 FreeSans 448 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 193228 -480 193340 240 0 FreeSans 448 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 196084 -480 196196 240 0 FreeSans 448 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 198940 -480 199052 240 0 FreeSans 448 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 201796 -480 201908 240 0 FreeSans 448 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 204652 -480 204764 240 0 FreeSans 448 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 207508 -480 207620 240 0 FreeSans 448 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 210364 -480 210476 240 0 FreeSans 448 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 213220 -480 213332 240 0 FreeSans 448 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 216076 -480 216188 240 0 FreeSans 448 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 218932 -480 219044 240 0 FreeSans 448 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 116116 -480 116228 240 0 FreeSans 448 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 221788 -480 221900 240 0 FreeSans 448 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 224644 -480 224756 240 0 FreeSans 448 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 227500 -480 227612 240 0 FreeSans 448 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 230356 -480 230468 240 0 FreeSans 448 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 233212 -480 233324 240 0 FreeSans 448 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 236068 -480 236180 240 0 FreeSans 448 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 238924 -480 239036 240 0 FreeSans 448 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 241780 -480 241892 240 0 FreeSans 448 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 244636 -480 244748 240 0 FreeSans 448 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 247492 -480 247604 240 0 FreeSans 448 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 118972 -480 119084 240 0 FreeSans 448 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 250348 -480 250460 240 0 FreeSans 448 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 253204 -480 253316 240 0 FreeSans 448 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 256060 -480 256172 240 0 FreeSans 448 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 258916 -480 259028 240 0 FreeSans 448 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 261772 -480 261884 240 0 FreeSans 448 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 264628 -480 264740 240 0 FreeSans 448 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 267484 -480 267596 240 0 FreeSans 448 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 270340 -480 270452 240 0 FreeSans 448 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 273196 -480 273308 240 0 FreeSans 448 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 276052 -480 276164 240 0 FreeSans 448 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 121828 -480 121940 240 0 FreeSans 448 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 278908 -480 279020 240 0 FreeSans 448 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 281764 -480 281876 240 0 FreeSans 448 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 284620 -480 284732 240 0 FreeSans 448 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 287476 -480 287588 240 0 FreeSans 448 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 124684 -480 124796 240 0 FreeSans 448 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 127540 -480 127652 240 0 FreeSans 448 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 130396 -480 130508 240 0 FreeSans 448 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 133252 -480 133364 240 0 FreeSans 448 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 108500 -480 108612 240 0 FreeSans 448 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 137060 -480 137172 240 0 FreeSans 448 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 139916 -480 140028 240 0 FreeSans 448 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 142772 -480 142884 240 0 FreeSans 448 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 145628 -480 145740 240 0 FreeSans 448 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 148484 -480 148596 240 0 FreeSans 448 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 151340 -480 151452 240 0 FreeSans 448 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 154196 -480 154308 240 0 FreeSans 448 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 157052 -480 157164 240 0 FreeSans 448 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 159908 -480 160020 240 0 FreeSans 448 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 162764 -480 162876 240 0 FreeSans 448 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 111356 -480 111468 240 0 FreeSans 448 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 165620 -480 165732 240 0 FreeSans 448 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 168476 -480 168588 240 0 FreeSans 448 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 171332 -480 171444 240 0 FreeSans 448 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 174188 -480 174300 240 0 FreeSans 448 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 177044 -480 177156 240 0 FreeSans 448 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 179900 -480 180012 240 0 FreeSans 448 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 182756 -480 182868 240 0 FreeSans 448 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 185612 -480 185724 240 0 FreeSans 448 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 188468 -480 188580 240 0 FreeSans 448 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 191324 -480 191436 240 0 FreeSans 448 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 114212 -480 114324 240 0 FreeSans 448 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 194180 -480 194292 240 0 FreeSans 448 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 197036 -480 197148 240 0 FreeSans 448 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 199892 -480 200004 240 0 FreeSans 448 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 202748 -480 202860 240 0 FreeSans 448 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 205604 -480 205716 240 0 FreeSans 448 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 208460 -480 208572 240 0 FreeSans 448 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 211316 -480 211428 240 0 FreeSans 448 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 214172 -480 214284 240 0 FreeSans 448 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 217028 -480 217140 240 0 FreeSans 448 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 219884 -480 219996 240 0 FreeSans 448 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 117068 -480 117180 240 0 FreeSans 448 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 222740 -480 222852 240 0 FreeSans 448 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 225596 -480 225708 240 0 FreeSans 448 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 228452 -480 228564 240 0 FreeSans 448 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 231308 -480 231420 240 0 FreeSans 448 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 234164 -480 234276 240 0 FreeSans 448 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 237020 -480 237132 240 0 FreeSans 448 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 239876 -480 239988 240 0 FreeSans 448 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 242732 -480 242844 240 0 FreeSans 448 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 245588 -480 245700 240 0 FreeSans 448 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 248444 -480 248556 240 0 FreeSans 448 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 119924 -480 120036 240 0 FreeSans 448 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 251300 -480 251412 240 0 FreeSans 448 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 254156 -480 254268 240 0 FreeSans 448 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 257012 -480 257124 240 0 FreeSans 448 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 259868 -480 259980 240 0 FreeSans 448 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 262724 -480 262836 240 0 FreeSans 448 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 265580 -480 265692 240 0 FreeSans 448 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 268436 -480 268548 240 0 FreeSans 448 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 271292 -480 271404 240 0 FreeSans 448 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 274148 -480 274260 240 0 FreeSans 448 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 277004 -480 277116 240 0 FreeSans 448 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 122780 -480 122892 240 0 FreeSans 448 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 279860 -480 279972 240 0 FreeSans 448 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 282716 -480 282828 240 0 FreeSans 448 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 285572 -480 285684 240 0 FreeSans 448 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 288428 -480 288540 240 0 FreeSans 448 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 125636 -480 125748 240 0 FreeSans 448 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 128492 -480 128604 240 0 FreeSans 448 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 131348 -480 131460 240 0 FreeSans 448 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 134204 -480 134316 240 0 FreeSans 448 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 289380 -480 289492 240 0 FreeSans 448 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 290332 -480 290444 240 0 FreeSans 448 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 291284 -480 291396 240 0 FreeSans 448 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 292236 -480 292348 240 0 FreeSans 448 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -478 -342 -168 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 -342 298510 -32 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -478 298344 298510 298654 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 298200 -342 298510 298654 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 1577 -822 1887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 10577 -822 10887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 19577 -822 19887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 28577 -822 28887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 37577 -822 37887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 46577 -822 46887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 55577 -822 55887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 55577 260603 55887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64577 -822 64887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 64577 260603 64887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 73577 -822 73887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 73577 260603 73887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 82577 -822 82887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 82577 260603 82887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 91577 -822 91887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 91577 260603 91887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 100577 -822 100887 49317 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 100577 100635 100887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 100577 260603 100887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 109577 -822 109887 49317 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 109577 100635 109887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 109577 260603 109887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 118577 -822 118887 49317 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 118577 100635 118887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 118577 260603 118887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 127577 -822 127887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 127577 260603 127887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 136577 -822 136887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 136577 260603 136887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 145577 -822 145887 124261 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 145577 260603 145887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 154577 -822 154887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 163577 -822 163887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 172577 -822 172887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 181577 -822 181887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 190577 -822 190887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 199577 -822 199887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 208577 -822 208887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 217577 -822 217887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 226577 -822 226887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 235577 -822 235887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 244577 -822 244887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 253577 -822 253887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 262577 -822 262887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 271577 -822 271887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 280577 -822 280887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 289577 -822 289887 299134 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 1913 298990 2223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 10913 298990 11223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 19913 298990 20223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 28913 298990 29223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 37913 298990 38223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 46913 298990 47223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 55913 298990 56223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 64913 298990 65223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 73913 298990 74223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 82913 298990 83223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 91913 298990 92223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 100913 298990 101223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 109913 298990 110223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 118913 298990 119223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 127913 298990 128223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 136913 298990 137223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 145913 298990 146223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 154913 298990 155223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 163913 298990 164223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 172913 298990 173223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 181913 298990 182223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 190913 298990 191223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 199913 298990 200223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 208913 298990 209223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 217913 298990 218223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 226913 298990 227223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 235913 298990 236223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 244913 298990 245223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 253913 298990 254223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 262913 298990 263223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 271913 298990 272223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 280913 298990 281223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -958 289913 298990 290223 0 FreeSans 2304 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -958 -822 -648 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 -822 298990 -512 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 298824 298990 299134 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 298680 -822 298990 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 3437 -822 3747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 12437 -822 12747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 21437 -822 21747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 30437 -822 30747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39437 -822 39747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 48437 -822 48747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 57437 -822 57747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 57437 182635 57747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 57437 260603 57747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66437 -822 66747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66437 182635 66747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 66437 260603 66747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 75437 -822 75747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 75437 184466 75747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 75437 260603 75747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 84437 -822 84747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 84437 182635 84747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 84437 260603 84747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 93437 -822 93747 49317 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 93437 100635 93747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 93437 182635 93747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 93437 260603 93747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 102437 -822 102747 49317 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 102437 100635 102747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 102437 182635 102747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 102437 260603 102747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 111437 -822 111747 49317 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 111437 100635 111747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 111437 182635 111747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 111437 260603 111747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 120437 -822 120747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 120437 182635 120747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 120437 260603 120747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 129437 -822 129747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 129437 182635 129747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 129437 260603 129747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 138437 -822 138747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 138437 182635 138747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 138437 260603 138747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 147437 -822 147747 124261 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 147437 182635 147747 199205 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 147437 260603 147747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 156437 -822 156747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 165437 -822 165747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 174437 -822 174747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 183437 -822 183747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 192437 -822 192747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 201437 -822 201747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 210437 -822 210747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 219437 -822 219747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 228437 -822 228747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 237437 -822 237747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 246437 -822 246747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 255437 -822 255747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 264437 -822 264747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 273437 -822 273747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 282437 -822 282747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 291437 -822 291747 299134 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 4913 298990 5223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 13913 298990 14223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 22913 298990 23223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 31913 298990 32223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 40913 298990 41223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 49913 298990 50223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 58913 298990 59223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 67913 298990 68223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 76913 298990 77223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 85913 298990 86223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 94913 298990 95223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 103913 298990 104223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 112913 298990 113223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 121913 298990 122223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 130913 298990 131223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 139913 298990 140223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 148913 298990 149223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 157913 298990 158223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 166913 298990 167223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 175913 298990 176223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 184913 298990 185223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 193913 298990 194223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 202913 298990 203223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 211913 298990 212223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 220913 298990 221223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 229913 298990 230223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 238913 298990 239223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 247913 298990 248223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 256913 298990 257223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 265913 298990 266223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 274913 298990 275223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 283913 298990 284223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -958 292913 298990 293223 0 FreeSans 2304 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 5684 -480 5796 240 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6636 -480 6748 240 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 7588 -480 7700 240 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 11396 -480 11508 240 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 43764 -480 43876 240 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 46620 -480 46732 240 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 49476 -480 49588 240 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 52332 -480 52444 240 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 55188 -480 55300 240 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 58044 -480 58156 240 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 60900 -480 61012 240 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 63756 -480 63868 240 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 66612 -480 66724 240 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 69468 -480 69580 240 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 15204 -480 15316 240 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 72324 -480 72436 240 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 75180 -480 75292 240 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 78036 -480 78148 240 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 80892 -480 81004 240 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 83748 -480 83860 240 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 86604 -480 86716 240 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 89460 -480 89572 240 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 92316 -480 92428 240 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 95172 -480 95284 240 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 98028 -480 98140 240 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 19012 -480 19124 240 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 100884 -480 100996 240 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 103740 -480 103852 240 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 22820 -480 22932 240 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 26628 -480 26740 240 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 29484 -480 29596 240 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 32340 -480 32452 240 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 35196 -480 35308 240 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 38052 -480 38164 240 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 40908 -480 41020 240 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 8540 -480 8652 240 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 12348 -480 12460 240 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 44716 -480 44828 240 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 47572 -480 47684 240 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 50428 -480 50540 240 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 53284 -480 53396 240 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 56140 -480 56252 240 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 58996 -480 59108 240 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 61852 -480 61964 240 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 64708 -480 64820 240 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 67564 -480 67676 240 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 70420 -480 70532 240 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 16156 -480 16268 240 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 73276 -480 73388 240 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 76132 -480 76244 240 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 78988 -480 79100 240 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 81844 -480 81956 240 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 84700 -480 84812 240 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 87556 -480 87668 240 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 90412 -480 90524 240 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 93268 -480 93380 240 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 96124 -480 96236 240 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 98980 -480 99092 240 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 19964 -480 20076 240 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 101836 -480 101948 240 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 104692 -480 104804 240 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 23772 -480 23884 240 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 27580 -480 27692 240 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 30436 -480 30548 240 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 33292 -480 33404 240 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 36148 -480 36260 240 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 39004 -480 39116 240 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 41860 -480 41972 240 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 13300 -480 13412 240 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 45668 -480 45780 240 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 48524 -480 48636 240 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 51380 -480 51492 240 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 54236 -480 54348 240 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 57092 -480 57204 240 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 59948 -480 60060 240 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 62804 -480 62916 240 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 65660 -480 65772 240 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 68516 -480 68628 240 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 71372 -480 71484 240 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 17108 -480 17220 240 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 74228 -480 74340 240 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 77084 -480 77196 240 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 79940 -480 80052 240 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 82796 -480 82908 240 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 85652 -480 85764 240 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 88508 -480 88620 240 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 91364 -480 91476 240 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 94220 -480 94332 240 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 97076 -480 97188 240 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 99932 -480 100044 240 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 20916 -480 21028 240 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 102788 -480 102900 240 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 105644 -480 105756 240 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 24724 -480 24836 240 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 28532 -480 28644 240 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 31388 -480 31500 240 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 34244 -480 34356 240 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 37100 -480 37212 240 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 39956 -480 40068 240 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 42812 -480 42924 240 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 14252 -480 14364 240 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 18060 -480 18172 240 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 21868 -480 21980 240 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 25676 -480 25788 240 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 9492 -480 9604 240 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 10444 -480 10556 240 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 144495 254161 144495 254161 0 vdd
rlabel via4 136815 257161 136815 257161 0 vss
rlabel metal3 296541 241444 296541 241444 0 io_in[12]
rlabel metal2 250740 196168 250740 196168 0 io_in[13]
rlabel metal3 297836 280812 297836 280812 0 io_in[14]
rlabel metal2 292348 218225 292348 218225 0 io_in[15]
rlabel metal2 258972 297836 258972 297836 0 io_in[16]
rlabel metal3 149940 201929 149940 201929 0 io_in[19]
rlabel metal2 151228 233240 151228 233240 0 io_in[20]
rlabel metal2 93884 296541 93884 296541 0 io_in[21]
rlabel metal2 60508 273238 60508 273238 0 io_in[22]
rlabel metal2 27216 297836 27216 297836 0 io_in[23]
rlabel metal3 296541 102676 296541 102676 0 io_in[5]
rlabel metal2 166740 88984 166740 88984 0 io_in[6]
rlabel metal3 297836 142128 297836 142128 0 io_in[7]
rlabel metal2 151620 113120 151620 113120 0 io_in[8]
rlabel metal2 152460 124768 152460 124768 0 io_in[9]
rlabel metal2 153300 153496 153300 153496 0 io_oeb[10]
rlabel metal3 297836 234584 297836 234584 0 io_oeb[11]
rlabel metal2 151340 168084 151340 168084 0 io_oeb[17]
rlabel metal2 151620 175532 151620 175532 0 io_oeb[18]
rlabel metal3 196 279160 196 279160 0 io_oeb[24]
rlabel metal3 1155 258412 1155 258412 0 io_oeb[25]
rlabel metal2 154140 140196 154140 140196 0 io_out[10]
rlabel metal2 155820 151844 155820 151844 0 io_out[11]
rlabel metal2 215124 296541 215124 296541 0 io_out[17]
rlabel metal2 176820 222852 176820 222852 0 io_out[18]
rlabel metal2 152068 254240 152068 254240 0 io_out[24]
rlabel metal3 196 264964 196 264964 0 io_out[25]
<< properties >>
string FIXED_BBOX 0 0 298020 298020
<< end >>
