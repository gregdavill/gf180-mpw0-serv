* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1343__B _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2106_ _0098_ net4 mod.cpu.bufreg2.i_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2037_ _0022_ net4 mod.cpu.bufreg2.i_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1270_ _0816_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1684__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1389__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A2 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1039__I1 mod.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1338__B _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1606_ mod.cpu.bufreg2.i_dat\[4\] _0323_ _0325_ _0819_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1537_ _0269_ _0680_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1468_ mod.cpu.ctrl.o_ibus_adr\[29\] _0972_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1399_ mod.cpu.bufreg.data\[15\] _0913_ _0917_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2052__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1197__A3 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1873__S _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1322_ mod.cpu.ctrl.o_ibus_adr\[0\] _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1253_ _0818_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1657__A1 mod.cpu.bufreg2.dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1184_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2075__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1693__S _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1706__B _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1940_ _0535_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1811__A1 mod.cpu.bufreg2.i_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1871_ _0510_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1305_ _0652_ mod.u_scanchain_local.module_data_in\[57\] _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1236_ _0805_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1167_ mod.cpu.immdec.imm11_7\[2\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2098__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1098_ mod.cpu.branch_op _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1577__I _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1436__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2070_ _0058_ net4 mod.u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1021_ mod.cpu.decode.opcode\[0\] _0616_ mod.cpu.decode.opcode\[2\] _0617_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ mod.cpu.ctrl.o_ibus_adr\[5\] _0540_ _0543_ mod.cpu.ctrl.o_ibus_adr\[6\] _0545_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1854_ _0495_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1785_ mod.cpu.immdec.imm19_12_20\[2\] _0397_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1012__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1219_ _0780_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1079__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2199_ _0190_ net3 mod.cpu.bufreg.data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2113__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1945__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1570_ _0775_ _0284_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _0113_ net3 mod.cpu.bufreg2.dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2053_ _0039_ net4 mod.u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2136__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1906_ _0533_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1837_ _0491_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1768_ mod.cpu.immdec.imm7 _0986_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1699_ _0759_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput7 net7 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2159__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1622_ mod.cpu.bufreg2.i_dat\[8\] _0336_ _0328_ mod.cpu.bufreg2.dat\[8\] _0337_ mod.cpu.bufreg2.dat\[9\]
+ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1553_ _0269_ mod.cpu.state.o_cnt_r\[0\] _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1484_ mod.cpu.bufreg.c_r _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1151__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2105_ _0097_ net4 mod.cpu.bufreg2.i_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2036_ _0021_ net4 mod.cpu.bufreg2.i_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1669__C1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1605_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1536_ _0756_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1467_ mod.u_scanchain_local.module_data_in\[92\] _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1398_ mod.cpu.ctrl.o_ibus_adr\[15\] _0907_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2019_ _0074_ net4 mod.cpu.bufreg2.i_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1115__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1321_ _0857_ mod.u_scanchain_local.module_data_in\[63\] _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1252_ mod.cpu.bufreg2.i_dat\[29\] mod.cpu.bufreg2.dat\[3\] _0817_ _0818_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1183_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1657__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1863__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1519_ _0252_ _0254_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1811__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1870_ mod.cpu.bufreg.data\[21\] mod.cpu.bufreg.data\[22\] _0506_ _0510_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1327__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1304_ mod.cpu.bufreg2.dat\[26\] _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1235_ _0722_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1166_ _0746_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1097_ _0674_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1802__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1999_ _0747_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1318__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2042__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2192__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1020_ mod.cpu.decode.opcode\[1\] _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1879__S _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1922_ _0544_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1853_ _0500_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1784_ _0438_ _0450_ _0454_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2065__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1218_ mod.cpu.bufreg2.i_dat\[21\] _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1079__A3 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2198_ _0189_ net3 mod.cpu.bufreg.data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1149_ _0731_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1711__A1 mod.cpu.bufreg2.i_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2088__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _0112_ net3 mod.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2052_ _0038_ net4 mod.u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1769__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1905_ _0806_ _0532_ _0529_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1836_ mod.cpu.bufreg.data\[6\] mod.cpu.bufreg.data\[7\] _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1767_ _0698_ _0729_ _0435_ _0437_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1698_ _0654_ _0762_ _0386_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2230__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1160__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1621_ _0320_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1552_ _0253_ _0278_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1691__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1483_ _0634_ _0985_ _0986_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2104_ _0096_ net4 mod.cpu.bufreg2.i_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2103__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2035_ _0020_ net4 mod.cpu.bufreg2.i_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1819_ mod.cpu.immdec.imm31 mod.cpu.bufreg2.i_dat\[31\] _0383_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1307__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1534__C _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1678__B1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__B1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1016__I mod.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1604_ _0294_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1535_ _0257_ _0268_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1466_ _0959_ _0971_ _0973_ _0974_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1397_ mod.u_scanchain_local.module_data_in\[78\] _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2018_ _0063_ net4 mod.cpu.bufreg2.i_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2149__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1320_ _0651_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1251_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1182_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1518_ _0253_ _0612_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1449_ mod.cpu.ctrl.o_ibus_adr\[25\] _0956_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1033__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1024__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1303_ _0846_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1234_ _0797_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1165_ mod.cpu.bufreg2.i_dat\[14\] mod.cpu.immdec.imm11_7\[1\] _0643_ _0746_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1204__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1096_ _0679_ _0680_ _0602_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1998_ _0588_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1114__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1050__S _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1006__A1 mod.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1557__A2 mod.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ mod.cpu.ctrl.o_ibus_adr\[4\] _0540_ _0543_ mod.cpu.ctrl.o_ibus_adr\[5\] _0544_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1852_ mod.cpu.bufreg.data\[13\] mod.cpu.bufreg.data\[14\] _0496_ _0500_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1783_ _0451_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1217_ _0791_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2197_ _0188_ net3 mod.cpu.bufreg.data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1148_ mod.cpu.ctrl.pc_plus_4_cy_r mod.cpu.ctrl.o_ibus_adr\[0\] _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1079_ _0657_ _0661_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1779__I _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2120_ _0111_ net3 mod.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2051_ _0037_ net4 mod.u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1769__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1904_ _0524_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _0484_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2032__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1766_ _0438_ _0437_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1697_ _0703_ _0759_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2182__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2249_ _0237_ net3 mod.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1209__A1 mod.cpu.bufreg2.i_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2055__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _0776_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1551_ _0266_ _0679_ mod.cpu.i_rf_ready _0783_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1482_ _0634_ mod.cpu.bufreg.c_r _0985_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2103_ _0095_ net4 mod.cpu.bufreg2.i_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2034_ _0018_ net4 mod.cpu.bufreg2.i_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1212__I _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1611__A1 _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _0645_ _0450_ _0480_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1749_ mod.cpu.bufreg2.i_dat\[26\] _0423_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1678__A1 mod.cpu.bufreg2.i_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1678__B2 mod.cpu.bufreg2.dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1669__B2 mod.cpu.bufreg2.dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1669__A1 mod.cpu.bufreg2.i_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1603_ _0777_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1534_ _0726_ _0265_ _0105_ _0778_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1207__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1465_ mod.cpu.bufreg.data\[28\] _0962_ _0966_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1396_ _0910_ _0915_ _0916_ _0918_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2220__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2017_ _0052_ net4 mod.cpu.bufreg2.i_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1787__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2000__A1 mod.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1250_ _0629_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2243__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1181_ mod.u_arbiter.i_wb_cpu_ack _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1814__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1517_ _0249_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1448_ mod.u_scanchain_local.module_data_in\[88\] _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1379_ mod.cpu.bufreg.data\[11\] _0897_ _0901_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2116__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1024__A2 mod.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1302_ mod.u_scanchain_local.module_data_in\[56\] mod.cpu.bufreg2.dat\[25\] _0843_
+ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1233_ mod.cpu.bufreg2.i_dat\[24\] _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1164_ _0745_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1095_ mod.cpu.state.o_cnt_r\[2\] _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2139__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1220__I _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ _0588_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ _0535_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1851_ _0499_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ _0395_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1215__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1216_ mod.cpu.bufreg2.i_dat\[20\] _0789_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2196_ _0187_ net3 mod.cpu.bufreg.data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1147_ _0680_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1078_ mod.cpu.state.o_cnt_r\[0\] _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1035__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ _0036_ net4 mod.u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1903_ mod.cpu.bufreg.data\[2\] _0522_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1834_ _0489_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1765_ mod.cpu.immdec.imm19_12_20\[0\] _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1696_ _0699_ _0379_ _0385_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2248_ _0236_ net3 mod.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2179_ _0170_ net3 mod.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1209__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1696__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1550_ _0253_ _0277_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ _0698_ _0684_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1136__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2102_ _0094_ net4 mod.cpu.bufreg2.i_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2033_ _0017_ net4 mod.cpu.bufreg2.i_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1611__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1817_ mod.cpu.bufreg2.i_dat\[19\] _0421_ _0449_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1748_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1375__A1 mod.cpu.bufreg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1679_ _0852_ _0327_ _0373_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1127__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1678__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1403__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1669__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2022__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2172__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1602_ _0766_ _0288_ _0319_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1533_ _0267_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1464_ mod.cpu.ctrl.o_ibus_adr\[28\] _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1395_ mod.cpu.bufreg.data\[14\] _0913_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2016_ _0041_ net4 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1596__A1 mod.cpu.bufreg2.i_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1899__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2195__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1339__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1180_ _0756_ mod.cpu.state.ibus_cyc _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1511__A1 mod.cpu.bufreg2.i_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1814__A2 mod.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1578__A1 mod.cpu.bufreg2.dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1050__I0 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1516_ _0760_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1218__I mod.cpu.bufreg2.i_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2068__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1447_ _0754_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1378_ mod.cpu.ctrl.o_ibus_adr\[11\] _0891_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1502__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1024__A3 mod.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2210__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1732__A1 mod.cpu.bufreg2.i_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1301_ _0845_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1232_ _0803_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1163_ mod.cpu.bufreg2.i_dat\[13\] mod.cpu.immdec.imm11_7\[0\] _0643_ _0745_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1094_ mod.cpu.state.o_cnt_r\[3\] _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1501__I _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1799__A1 mod.cpu.bufreg2.i_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ _0444_ _0590_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1723__A1 mod.cpu.bufreg2.i_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2233__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1493__A3 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ mod.cpu.bufreg.data\[12\] mod.cpu.bufreg.data\[13\] _0496_ _0499_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1781_ mod.cpu.immdec.imm19_12_20\[1\] _0252_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1477__B _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1705__A1 mod.cpu.bufreg2.i_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1181__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2106__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1215_ _0630_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2195_ _0186_ net3 mod.cpu.bufreg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1146_ _0662_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2256__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1077_ mod.cpu.mem_bytecnt\[0\] mod.cpu.state.o_cnt\[2\] mod.cpu.mem_bytecnt\[1\]
+ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _0579_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2129__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1252__S _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1902_ _0805_ _0529_ _0530_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1833_ mod.cpu.bufreg.data\[5\] mod.cpu.bufreg.data\[6\] _0485_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1764_ _0984_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ mod.cpu.bufreg2.i_dat\[4\] _0380_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0235_ net3 mod.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2178_ _0169_ net3 mod.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1129_ _0708_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1081__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ _0984_ _0729_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1046__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2101_ _0093_ net4 mod.cpu.bufreg2.i_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2032_ _0016_ net4 mod.cpu.bufreg2.i_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1816_ _0397_ _0477_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1747_ _0760_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1678_ mod.cpu.bufreg2.i_dat\[29\] _0777_ _0328_ mod.cpu.bufreg2.dat\[29\] _0373_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1601_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1532_ _0249_ _0266_ _0764_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1463_ _0923_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1394_ _0867_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _0030_ net4 mod.cpu.i_timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1324__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1511__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1515_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1446_ _0943_ _0955_ _0957_ _0958_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1377_ mod.u_scanchain_local.module_data_in\[74\] _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1502__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1018__A1 mod.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2012__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2162__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1144__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1255__S _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1300_ mod.u_scanchain_local.module_data_in\[55\] mod.cpu.bufreg2.dat\[24\] _0843_
+ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1231_ mod.cpu.bufreg2.i_dat\[23\] _0793_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1162_ _0737_ _0738_ _0740_ _0744_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1093_ _0673_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1995_ _0393_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2035__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1271__I1 mod.cpu.bufreg2.dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2185__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1723__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1429_ mod.cpu.ctrl.o_ibus_adr\[21\] _0940_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1239__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1262__I1 mod.cpu.bufreg2.dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1478__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2058__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2433__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1780_ _0448_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1214_ _0655_ _0786_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2194_ _0185_ net3 mod.cpu.bufreg.data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1145_ _0683_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1076_ _0606_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__A1 mod.cpu.bufreg2.dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__B _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1978_ mod.cpu.ctrl.o_ibus_adr\[26\] _0578_ _0575_ mod.cpu.ctrl.o_ibus_adr\[27\]
+ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2200__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1578__B _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1901_ _0806_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1832_ _0488_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1763_ _0697_ _0675_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1694_ _0384_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1507__I mod.cpu.bufreg2.i_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2246_ _0234_ net3 mod.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2223__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ _0168_ net3 mod.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1128_ _0693_ _0700_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1059_ mod.cpu.immdec.imm19_12_20\[8\] _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2006__C _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1081__A2 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2246__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0091_ net4 mod.u_scanchain_local.module_data_in\[95\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2031_ _0015_ net4 mod.cpu.bufreg2.i_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1062__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1815_ _0778_ _0435_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1746_ mod.cpu.immdec.imm30_25\[2\] mod.cpu.immdec.imm30_25\[1\] _0419_ _0423_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1677_ _0372_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2229_ _0217_ net3 mod.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2119__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1600_ _0289_ _0284_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1531_ _0612_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1462_ mod.u_scanchain_local.module_data_in\[91\] _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1393_ mod.cpu.ctrl.o_ibus_adr\[14\] _0907_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1817__A1 mod.cpu.bufreg2.i_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _0019_ net4 mod.cpu.i_rf_ready vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1729_ mod.cpu.immdec.imm24_20\[2\] _0406_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1430__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2091__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1586__B _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1605__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__B1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1514_ _0604_ _0739_ _0249_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1445_ mod.cpu.bufreg.data\[24\] _0946_ _0950_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1515__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1376_ _0894_ _0899_ _0900_ _0902_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1250__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__C1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__B1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1230_ _0722_ _0800_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1161_ mod.cpu.immdec.imm11_7\[4\] _0741_ _0743_ _0728_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1496__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1092_ _0675_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1070__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1994_ mod.cpu.immdec.imm11_7\[0\] mod.cpu.immdec.imm11_7\[1\] _0588_ _0589_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1420__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1428_ mod.u_scanchain_local.module_data_in\[84\] _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1487__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1359_ mod.cpu.bufreg.data\[7\] _0881_ _0885_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1411__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1155__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1104__B _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1213_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ _0184_ net3 mod.cpu.bufreg.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1469__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1144_ _0629_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1075_ _0658_ _0608_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1641__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2152__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0558_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2025__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2175__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ _0522_ _0996_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ mod.cpu.bufreg.data\[4\] mod.cpu.bufreg.data\[5\] _0485_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1762_ mod.cpu.immdec.imm31 _0620_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1693_ _0984_ mod.cpu.bufreg2.i_dat\[3\] _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1139__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2245_ _0233_ net3 mod.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2176_ _0167_ net3 mod.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1127_ _0700_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1058_ _0644_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2048__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1550__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2198__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1589__B _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1081__A3 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1541__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2030_ _0014_ net4 mod.cpu.bufreg2.i_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1814_ _0701_ mod.cpu.immdec.imm24_20\[0\] _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ _0422_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1676_ mod.cpu.bufreg2.i_dat\[28\] _0293_ _0324_ mod.cpu.bufreg2.dat\[28\] _0359_
+ mod.cpu.bufreg2.dat\[29\] _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2228_ _0216_ net3 mod.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2159_ _0150_ net3 mod.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1523__A1 mod.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2213__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _0667_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1461_ _0959_ _0968_ _0969_ _0970_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1392_ mod.u_scanchain_local.module_data_in\[77\] _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1514__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1817__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0008_ net4 mod.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1022__B mod.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1728_ mod.cpu.bufreg2.i_dat\[22\] _0378_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1659_ _0361_ _0362_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1808__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2236__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1044__I0 mod.cpu.i_rf_ready vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1621__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1735__A1 mod.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ net3 _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1444_ mod.cpu.ctrl.o_ibus_adr\[24\] _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1375_ mod.cpu.bufreg.data\[10\] _0897_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1531__I _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2259__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1671__B1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__B1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__C2 mod.cpu.bufreg2.dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1717__B2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1717__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1160_ _0725_ _0703_ _0742_ _0682_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1091_ mod.cpu.decode.co_mem_word _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _0782_ _0743_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1427_ _0754_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2081__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1358_ mod.cpu.ctrl.o_ibus_adr\[7\] _0874_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1289_ mod.u_scanchain_local.module_data_in\[50\] mod.cpu.bufreg2.dat\[19\] _0838_
+ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1261__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1210__B _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1635__C2 mod.cpu.bufreg2.dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1346__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1282__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1212_ _0774_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2192_ _0183_ net3 mod.cpu.bufreg.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1143_ _0658_ _0724_ _0726_ _0655_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1074_ _0610_ _0624_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1976_ _0577_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1157__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1093__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1084__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _0487_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1761_ mod.cpu.bufreg2.i_dat\[30\] _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1692_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1139__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2244_ _0232_ net3 mod.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2175_ _0166_ net3 mod.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1126_ _0709_ _0710_ _0622_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1057_ mod.cpu.bufreg2.i_dat\[2\] mod.cpu.immdec.imm19_12_20\[7\] _0643_ _0644_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1075__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1959_ _0567_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1714__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1624__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1541__A2 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2142__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1813_ _0451_ _0475_ _0476_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1744_ mod.cpu.bufreg2.i_dat\[25\] _0420_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1675_ _0370_ _0371_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _0215_ net3 mod.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2158_ _0149_ net3 mod.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1109_ mod.cpu.alu.cmp_r _0664_ _0671_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2089_ _0079_ net4 mod.u_scanchain_local.module_data_in\[84\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2015__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2165__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1523__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1211__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1460_ mod.cpu.bufreg.data\[27\] _0962_ _0966_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1391_ _0910_ _0911_ _0912_ _0914_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1354__I _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1514__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0004_ net4 mod.cpu.bufreg2.i_rs2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2038__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1727_ mod.cpu.immdec.imm24_20\[3\] _0387_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2188__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1658_ mod.cpu.bufreg2.i_dat\[20\] _0336_ _0351_ mod.cpu.bufreg2.dat\[20\] _0362_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1589_ _0307_ _0309_ _0303_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1441__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1680__A1 mod.cpu.bufreg2.i_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1432__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1349__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1512_ _0248_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1443_ _0923_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1374_ _0867_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1120__B1 mod.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1671__B2 mod.cpu.bufreg2.dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1671__A1 mod.cpu.bufreg2.i_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__B2 mod.cpu.bufreg2.dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__A1 mod.cpu.bufreg2.i_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1169__I _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1632__I _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1090_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1992_ _0585_ _0587_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1426_ _0927_ _0939_ _0941_ _0942_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2226__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1357_ mod.u_scanchain_local.module_data_in\[70\] _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1288_ _0780_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1635__A1 mod.cpu.bufreg2.i_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2249__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1211_ _0673_ _0701_ _0783_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1362__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2191_ _0182_ net3 mod.cpu.bufreg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1142_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1073_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1975_ mod.cpu.ctrl.o_ibus_adr\[25\] _0572_ _0575_ mod.cpu.ctrl.o_ibus_adr\[26\]
+ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1409_ mod.cpu.ctrl.o_ibus_adr\[17\] _0924_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1165__I0 mod.cpu.bufreg2.i_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1617__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1447__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _0377_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2071__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1691_ _0376_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1293__S _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _0231_ net3 mod.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2174_ _0165_ net3 mod.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1125_ mod.cpu.mem_bytecnt\[0\] mod.cpu.state.o_cnt\[2\] _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1056_ _0630_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1958_ mod.cpu.ctrl.o_ibus_adr\[18\] _0566_ _0563_ mod.cpu.ctrl.o_ibus_adr\[19\]
+ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1889_ _0520_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1138__I0 mod.cpu.bufreg2.dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2094__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1126__B _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__I _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2006__A1 mod.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1812_ mod.cpu.immdec.imm19_12_20\[7\] _0457_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1743_ _0758_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1674_ mod.cpu.bufreg2.i_dat\[27\] _0336_ _0331_ mod.cpu.bufreg2.dat\[27\] _0371_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1751__S _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1532__A3 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2226_ _0214_ net3 mod.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2157_ _0148_ net3 mod.cpu.bufreg2.i_op_b_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1108_ mod.cpu.bufreg.lsb\[0\] _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2088_ _0078_ net4 mod.u_scanchain_local.module_data_in\[83\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1039_ mod.cpu.bufreg2.i_rs2 mod.cpu.immdec.imm24_20\[1\] _0631_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1211__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1836__S _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1390_ mod.cpu.bufreg.data\[13\] _0913_ _0901_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0591_ _0599_ _0600_ _0601_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1746__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1726_ _0402_ _0404_ _0405_ _0407_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1657_ mod.cpu.bufreg2.dat\[21\] _0349_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _0814_ _0302_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _0200_ net3 mod.cpu.bufreg.data\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2132__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1455__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1752__I0 mod.cpu.bufreg2.i_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1190__I mod.cpu.bufreg2.dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1680__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1196__A1 mod.cpu.bufreg2.dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1511_ mod.cpu.bufreg2.i_dat\[12\] _0857_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_99_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1442_ mod.u_scanchain_local.module_data_in\[87\] _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1373_ mod.cpu.ctrl.o_ibus_adr\[10\] _0891_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1671__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2155__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1187__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1709_ _0658_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1662__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2028__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2178__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1991_ mod.cpu.ctrl.i_jump _0733_ _0581_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1425_ mod.cpu.bufreg.data\[20\] _0930_ _0934_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1356_ _0878_ _0883_ _0884_ _0886_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1287_ _0837_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1908__I _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1210_ _0779_ _0784_ _0785_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2190_ _0181_ net3 mod.cpu.bufreg.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1141_ _0686_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1072_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1974_ _0576_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1754__S _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1408_ mod.u_scanchain_local.module_data_in\[80\] _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1165__I1 mod.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1314__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1339_ _0855_ _0870_ _0871_ _0872_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1617__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1463__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1305__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2216__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1690_ _0698_ _0379_ _0381_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1544__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2242_ _0230_ net3 mod.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2173_ _0164_ net3 mod.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1124_ mod.cpu.mem_bytecnt\[1\] _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1055_ _0642_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1749__S _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1957_ _0558_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1888_ mod.cpu.bufreg.data\[29\] mod.cpu.bufreg.data\[30\] _0516_ _0520_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1138__I1 mod.cpu.bufreg2.dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2239__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1774__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1526__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ mod.cpu.bufreg2.i_dat\[18\] _0433_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1742_ mod.cpu.immdec.imm30_25\[1\] mod.cpu.immdec.imm30_25\[0\] _0419_ _0420_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1673_ mod.cpu.bufreg2.dat\[28\] _0321_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2225_ _0213_ net3 mod.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2156_ _0147_ net3 mod.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1107_ mod.cpu.state.stage_two_req _0672_ _0678_ _0681_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2087_ _0077_ net4 mod.u_scanchain_local.module_data_in\[82\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1038_ _0632_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1741__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1188__I _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1211__A3 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ mod.cpu.immdec.imm30_25\[0\] _0421_ _0591_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1098__I mod.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1725_ mod.cpu.immdec.imm24_20\[1\] _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1826__I _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1656_ _0360_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1587_ _0300_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2084__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1561__I _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2208_ _0199_ net3 mod.cpu.bufreg.data\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2139_ _0130_ net3 mod.cpu.bufreg2.dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1196__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1510_ _0247_ _0738_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1441_ _0943_ _0952_ _0953_ _0954_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1372_ mod.u_scanchain_local.module_data_in\[73\] _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1757__S _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1187__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1708_ _0759_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1639_ _0348_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1102__A2 mod.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1990_ mod.cpu.ctrl.i_jump _0716_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1424_ mod.cpu.ctrl.o_ibus_adr\[20\] _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1355_ mod.cpu.bufreg.data\[6\] _0881_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1286_ mod.u_scanchain_local.module_data_in\[49\] mod.cpu.bufreg2.dat\[18\] _0833_
+ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2122__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1096__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2145__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1140_ _0718_ _0719_ _0721_ _0724_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1071_ mod.cpu.csr_d_sel _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1087__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1882__I0 mod.cpu.bufreg.data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1973_ mod.cpu.ctrl.o_ibus_adr\[24\] _0572_ _0575_ mod.cpu.ctrl.o_ibus_adr\[25\]
+ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1562__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1407_ _0877_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1338_ mod.cpu.bufreg.data\[3\] _0795_ _0868_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1269_ _0827_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1078__A1 mod.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2168__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1553__A2 mod.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1654__I _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2241_ _0229_ net3 mod.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0163_ net3 mod.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1123_ mod.cpu.ctrl.pc_plus_offset_cy_r _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1054_ mod.cpu.bufreg2.i_dat\[1\] mod.cpu.immdec.imm19_12_20\[6\] _0637_ _0642_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1480__A1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1956_ _0565_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1887_ _0519_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1564__I _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1535__A2 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1138__I2 mod.cpu.bufreg2.dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1846__I0 mod.cpu.bufreg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1223__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1810_ _0645_ _0403_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1741_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1672_ _0847_ _0325_ _0369_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2224_ _0212_ net3 mod.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2155_ _0146_ net3 mod.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1106_ _0682_ _0684_ _0689_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2086_ _0076_ net4 mod.u_scanchain_local.module_data_in\[81\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1037_ net1 mod.cpu.immdec.imm24_20\[0\] _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1939_ _0554_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1508__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2206__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1295__I1 mod.cpu.bufreg2.dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1724_ _0400_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1655_ mod.cpu.bufreg2.i_dat\[19\] _0347_ _0355_ mod.cpu.bufreg2.dat\[19\] _0359_
+ mod.cpu.bufreg2.dat\[20\] _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_1586_ _0810_ mod.cpu.bufreg2.dat\[1\] _0814_ _0285_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2229__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2207_ _0198_ net3 mod.cpu.bufreg.data\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2138_ _0129_ net3 mod.cpu.bufreg2.dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1674__B2 mod.cpu.bufreg2.dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1674__A1 mod.cpu.bufreg2.i_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2069_ _0057_ net4 mod.u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1277__I1 mod.cpu.bufreg2.dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1665__B2 mod.cpu.bufreg2.dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__A1 mod.cpu.bufreg2.i_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1268__I1 mod.cpu.bufreg2.dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1968__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1440_ mod.cpu.bufreg.data\[23\] _0946_ _0950_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1371_ _0894_ _0895_ _0896_ _0898_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1259__I1 mod.cpu.bufreg2.dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2051__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1707_ mod.cpu.bufreg2.i_dat\[14\] _0382_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1638_ mod.cpu.bufreg2.i_dat\[14\] _0347_ _0341_ mod.cpu.bufreg2.dat\[14\] _0344_
+ mod.cpu.bufreg2.dat\[15\] _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1569_ _0776_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__A1 mod.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1747__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1638__A1 mod.cpu.bufreg2.i_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1638__B2 mod.cpu.bufreg2.dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2074__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1810__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1423_ _0923_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1354_ _0867_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1285_ _0836_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_180 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2097__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1161__B _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1070_ _0619_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1087__A2 mod.cpu.bufreg2.dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _0562_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1406_ _0910_ _0922_ _0925_ _0926_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1337_ mod.cpu.ctrl.o_ibus_adr\[3\] _0861_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1268_ mod.u_scanchain_local.module_data_in\[41\] mod.cpu.bufreg2.dat\[10\] _0823_
+ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1199_ _0639_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2112__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1935__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2240_ _0228_ net3 mod.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2171_ _0162_ net3 mod.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1122_ mod.cpu.ctrl.o_ibus_adr\[0\] _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1053_ _0641_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2009__A1 mod.cpu.bufreg2.i_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1480__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1955_ mod.cpu.ctrl.o_ibus_adr\[17\] _0559_ _0563_ mod.cpu.ctrl.o_ibus_adr\[18\]
+ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1886_ mod.cpu.bufreg.data\[28\] mod.cpu.bufreg.data\[29\] _0516_ _0519_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1845__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1138__I3 mod.cpu.bufreg2.dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2135__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1223__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1774__A3 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1704__B _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1740_ _0604_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1671_ mod.cpu.bufreg2.i_dat\[26\] _0291_ _0327_ mod.cpu.bufreg2.dat\[27\] _0369_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ _0211_ net3 mod.cpu.ctrl.o_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2154_ _0145_ net3 mod.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1105_ mod.cpu.state.init_done _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1150__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ _0075_ net4 mod.u_scanchain_local.module_data_in\[80\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1036_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2158__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ mod.cpu.ctrl.o_ibus_adr\[11\] _0552_ _0549_ mod.cpu.ctrl.o_ibus_adr\[12\]
+ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1869_ _0509_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1819__I1 mod.cpu.bufreg2.i_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1755__I0 mod.cpu.bufreg2.i_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1683__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1199__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1723_ mod.cpu.bufreg2.i_dat\[21\] _0397_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1994__I0 mod.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ _0332_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1585_ mod.cpu.bufreg2.dat\[3\] _0771_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _0197_ net3 mod.cpu.bufreg.data\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2137_ _0128_ net3 mod.cpu.bufreg2.dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1674__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2068_ _0056_ net4 mod.u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1019_ _0613_ mod.cpu.immdec.imm11_7\[0\] _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1665__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1370_ mod.cpu.bufreg.data\[9\] _0897_ _0885_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1706_ _0661_ _0380_ _0391_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1637_ _0776_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1568_ _0812_ _0288_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1344__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1499_ _1000_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1895__A2 mod.cpu.bufreg.data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1583__A1 mod.cpu.bufreg2.i_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1335__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1638__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1810__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1422_ mod.u_scanchain_local.module_data_in\[83\] _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1353_ mod.cpu.ctrl.o_ibus_adr\[6\] _0874_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1284_ mod.u_scanchain_local.module_data_in\[48\] mod.cpu.bufreg2.dat\[17\] _0833_
+ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_170 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2156__D _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1565__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1161__C _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ _0574_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2191__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1405_ mod.cpu.bufreg.data\[16\] _0913_ _0917_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1336_ mod.u_scanchain_local.module_data_in\[66\] _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput1 io_in[12] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1267_ _0826_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1198_ _0756_ mod.cpu.state.ibus_cyc _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1786__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2064__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1777__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1951__I _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _0161_ net3 mod.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1701__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1121_ _0614_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1052_ mod.cpu.bufreg2.i_dat\[0\] mod.cpu.immdec.imm19_12_20\[5\] _0637_ _0641_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2009__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0564_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1885_ _0518_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2087__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1319_ _0854_ _0855_ _0856_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1302__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1101__I mod.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1670_ _0368_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _0210_ net3 mod.cpu.ctrl.o_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2153_ _0144_ net3 mod.cpu.bufreg2.dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1104_ _0685_ _0687_ _0688_ _0619_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1150__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2084_ _0073_ net4 mod.u_scanchain_local.module_data_in\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1035_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ _0553_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1610__B1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ mod.cpu.bufreg.data\[20\] mod.cpu.bufreg.data\[21\] _0506_ _0509_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1792__S _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ mod.cpu.bufreg2.i_dat\[15\] _0383_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2102__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2252__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__S _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1199__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1722_ mod.cpu.immdec.imm24_20\[2\] _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1653_ _0357_ _0358_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1994__I1 mod.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1584_ _0306_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2125__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0196_ net3 mod.cpu.bufreg.data\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _0127_ net3 mod.cpu.bufreg2.dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2067_ _0055_ net4 mod.u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1018_ mod.cpu.decode.opcode\[0\] mod.cpu.decode.opcode\[1\] mod.cpu.decode.opcode\[2\]
+ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_81_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2148__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1445__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ mod.cpu.bufreg2.i_dat\[13\] _0382_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1636_ _0346_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1567_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1498_ mod.cpu.bufreg2.i_dat\[4\] _0857_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2119_ _0110_ net3 mod.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1032__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ _0927_ _0936_ _0937_ _0938_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1890__S _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1352_ mod.u_scanchain_local.module_data_in\[69\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1283_ _0835_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_160 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_171 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1565__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1619_ _0737_ _0330_ _0335_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1970_ mod.cpu.ctrl.o_ibus_adr\[23\] _0572_ _0569_ mod.cpu.ctrl.o_ibus_adr\[24\]
+ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1404_ mod.cpu.ctrl.o_ibus_adr\[16\] _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1335_ _0855_ _0865_ _0866_ _0869_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput2 io_in[13] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1266_ mod.u_scanchain_local.module_data_in\[40\] mod.cpu.bufreg2.dat\[9\] _0823_
+ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1197_ _0658_ _0661_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1483__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2209__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1474__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1226__A1 mod.cpu.bufreg2.i_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1009__I _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1162__B1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1120_ _0686_ _0616_ mod.cpu.decode.co_ebreak _0702_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1051_ _0640_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1953_ mod.cpu.ctrl.o_ibus_adr\[16\] _0559_ _0563_ mod.cpu.ctrl.o_ibus_adr\[17\]
+ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1768__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ mod.cpu.bufreg.data\[27\] mod.cpu.bufreg.data\[28\] _0516_ _0518_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1318_ _0652_ mod.u_scanchain_local.module_data_in\[62\] _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1249_ _0815_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1456__A1 mod.cpu.bufreg.data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1208__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2031__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2181__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1695__A1 mod.cpu.bufreg2.i_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1298__I1 mod.cpu.bufreg2.dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _0002_ net3 mod.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ _0143_ net3 mod.cpu.bufreg2.dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1103_ mod.cpu.csr_d_sel mod.cpu.decode.co_mem_word _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1150__A3 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2083_ _0072_ net4 mod.u_scanchain_local.module_data_in\[78\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1034_ net2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1289__I1 mod.cpu.bufreg2.dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1202__I _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1989__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1936_ mod.cpu.ctrl.o_ibus_adr\[10\] _0552_ _0549_ mod.cpu.ctrl.o_ibus_adr\[11\]
+ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1867_ _0508_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1798_ mod.cpu.immdec.imm19_12_20\[5\] _0424_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1872__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1112__I mod.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1721_ _0377_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1652_ mod.cpu.bufreg2.i_dat\[18\] _0323_ _0351_ mod.cpu.bufreg2.dat\[18\] _0358_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ mod.cpu.bufreg2.i_dat\[1\] _0298_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _0195_ net3 mod.cpu.bufreg.data\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ _0126_ net3 mod.cpu.bufreg2.dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2066_ _0054_ net4 mod.u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1017_ mod.cpu.bufreg2.i_op_b_sel _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _0542_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1017__I mod.cpu.bufreg2.i_op_b_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1704_ _0607_ _0379_ _0390_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1635_ mod.cpu.bufreg2.i_dat\[13\] _0339_ _0341_ mod.cpu.bufreg2.dat\[13\] _0344_
+ mod.cpu.bufreg2.dat\[14\] _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1566_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1497_ _0998_ _0999_ _0740_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2242__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2118_ _0109_ net3 mod.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2049_ _0035_ net4 mod.u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2115__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ mod.cpu.bufreg.data\[19\] _0930_ _0934_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1351_ _0878_ _0879_ _0880_ _0882_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1282_ mod.u_scanchain_local.module_data_in\[47\] mod.cpu.bufreg2.dat\[16\] _0833_
+ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_150 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_161 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_172 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1618_ mod.cpu.bufreg2.dat\[7\] _0331_ _0333_ mod.cpu.bufreg2.dat\[8\] _0335_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1549_ _0709_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2138__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1403_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1334_ mod.cpu.bufreg.data\[2\] _0795_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1265_ _0825_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 io_in[15] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1196_ mod.cpu.bufreg2.dat\[6\] _0765_ _0769_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1226__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1162__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1050_ _0639_ mod.cpu.csr_imm _0637_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1465__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1952_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1622__C1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1883_ _0517_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1153__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1317_ _0754_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1248_ mod.cpu.bufreg2.i_dat\[28\] _0814_ _0790_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1456__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1179_ net3 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1208__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1758__I0 mod.cpu.bufreg2.i_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _0003_ net3 mod.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _0142_ net3 mod.cpu.bufreg2.dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1102_ _0686_ mod.cpu.branch_op _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2082_ _0071_ net4 mod.u_scanchain_local.module_data_in\[77\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1033_ _0605_ _0609_ _0628_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1935_ _0539_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1610__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ mod.cpu.bufreg.data\[19\] mod.cpu.bufreg.data\[20\] _0506_ _0508_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1749__I0 mod.cpu.bufreg2.i_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1797_ _0464_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1117__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1720_ _0400_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ mod.cpu.bufreg2.dat\[19\] _0349_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1582_ _0299_ _0302_ _0303_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1108__A1 mod.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2203_ _0194_ net3 mod.cpu.bufreg.data\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2134_ _0125_ net3 mod.cpu.bufreg2.dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2021__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2065_ _0053_ net4 mod.u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1213__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1016_ mod.cpu.bufreg2.i_cnt_done _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2171__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1595__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ mod.cpu.ctrl.o_ibus_adr\[3\] _0540_ _0536_ mod.cpu.ctrl.o_ibus_adr\[4\] _0542_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ _0498_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2044__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2194__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1703_ mod.cpu.bufreg2.i_dat\[12\] _0382_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ _0345_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1565_ _0639_ _0774_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1496_ _0680_ _0730_ _0732_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2117_ _0108_ net3 mod.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2048_ _0034_ net4 mod.u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1804__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1118__I mod.cpu.bufreg2.i_op_b_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2067__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1740__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1054__S _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1350_ mod.cpu.bufreg.data\[5\] _0881_ _0868_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1281_ _0834_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_151 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_140 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_162 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_173 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output5_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1617_ _1001_ _0330_ _0334_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1548_ _0720_ _0274_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1479_ _0616_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1557__B mod.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1713__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2232__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1252__I0 mod.cpu.bufreg2.i_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ _0757_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1704__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1333_ _0867_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1264_ mod.u_scanchain_local.module_data_in\[39\] mod.cpu.bufreg2.dat\[8\] _0823_
+ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_90 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1307__I1 mod.cpu.bufreg2.dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[8] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
X_1195_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1483__A3 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1221__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1171__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2105__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2255__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1162__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1242__S _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0534_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1622__B1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1622__C2 mod.cpu.bufreg2.dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ mod.cpu.bufreg.data\[26\] mod.cpu.bufreg.data\[27\] _0516_ _0517_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2434_ net2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2128__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1316_ mod.cpu.bufreg2.dat\[31\] _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1247_ mod.cpu.bufreg2.dat\[2\] _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1178_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1208__A3 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1216__I0 mod.cpu.bufreg2.i_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1036__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2150_ _0141_ net3 mod.cpu.bufreg2.dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1101_ mod.cpu.decode.opcode\[0\] _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2081_ _0070_ net4 mod.u_scanchain_local.module_data_in\[76\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1032_ _0605_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1934_ _0551_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1865_ _0507_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ mod.cpu.immdec.imm19_12_20\[3\] _0463_ _0449_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1117__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ _0356_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1581_ _0812_ _0287_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1108__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2202_ _0193_ net3 mod.cpu.bufreg.data\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2133_ _0124_ net3 mod.cpu.bufreg2.dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2064_ _0051_ net4 mod.u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1015_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1917_ _0541_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1848_ mod.cpu.bufreg.data\[11\] mod.cpu.bufreg.data\[12\] _0496_ _0498_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1779_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1338__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1510__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__I0 mod.cpu.bufreg.data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1026__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1702_ _1001_ _0762_ _0389_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1633_ mod.cpu.bufreg2.i_dat\[12\] _0339_ _0341_ mod.cpu.bufreg2.dat\[12\] _0344_
+ mod.cpu.bufreg2.dat\[13\] _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1564_ _0285_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1495_ mod.cpu.ctrl.pc_plus_4_cy_r _0859_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1224__I mod.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2116_ _0107_ net3 mod.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2047_ _0033_ net4 mod.u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1245__S _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1280_ mod.u_scanchain_local.module_data_in\[46\] mod.cpu.bufreg2.dat\[15\] _0833_
+ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_141 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2161__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_130 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_152 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_174 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_163 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1798__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1616_ mod.cpu.bufreg2.dat\[6\] _0331_ _0333_ mod.cpu.bufreg2.dat\[7\] _0334_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1970__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1722__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1547_ _0720_ _0274_ _0275_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1478_ _0755_ _0981_ _0982_ _0983_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1486__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2034__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1557__C mod.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2184__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1477__A1 mod.cpu.bufreg.data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1229__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1401_ mod.u_scanchain_local.module_data_in\[79\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1704__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1332_ _0650_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1263_ _0824_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_91 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_80 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1194_ _0739_ _0677_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2057__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1568__B _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1698__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1950_ _0561_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1622__A1 mod.cpu.bufreg2.i_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1622__B2 mod.cpu.bufreg2.dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1881_ _0692_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2433_ net4 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1689__A1 mod.cpu.bufreg2.i_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1315_ _0852_ _0748_ _0853_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1246_ _0813_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1177_ _0650_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1216__I1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1407__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2222__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1907__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1317__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1100_ mod.cpu.decode.co_mem_word mod.cpu.bne_or_bge _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0069_ net4 mod.u_scanchain_local.module_data_in\[75\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1031_ _0611_ _0624_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ mod.cpu.ctrl.o_ibus_adr\[9\] _0546_ _0549_ mod.cpu.ctrl.o_ibus_adr\[10\] _0551_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ mod.cpu.bufreg.data\[18\] mod.cpu.bufreg.data\[19\] _0506_ _0507_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1795_ _0392_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2245__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1229_ _0718_ _0651_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1137__I mod.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2118__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1248__S _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ _0290_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ _0192_ net3 mod.cpu.bufreg.data\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2132_ _0123_ net3 mod.cpu.bufreg2.dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2063_ _0050_ net4 mod.u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1816__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1014_ mod.cpu.alu.i_rs1 mod.cpu.alu.add_cy_r _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1916_ mod.cpu.ctrl.o_ibus_adr\[2\] _0540_ _0536_ mod.cpu.ctrl.o_ibus_adr\[3\] _0541_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1847_ _0497_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1778_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__A1 mod.cpu.bufreg2.i_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1586__A3 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1897__I1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1701_ _0778_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1632_ _0332_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1563_ _0284_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1494_ _0997_ _0714_ _0740_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1505__I mod.cpu.bufreg2.i_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2115_ _0106_ net3 mod.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2046_ _0032_ net4 mod.u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1415__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1879__I1 mod.cpu.bufreg.data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_131 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_142 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_120 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_164 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_175 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_153 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1060__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1615_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1546_ _0720_ _0274_ _0269_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1235__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1477_ mod.cpu.bufreg.data\[31\] _0788_ _0648_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1486__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2029_ _0013_ net4 mod.cpu.bufreg2.i_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1477__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1229__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ _0910_ _0919_ _0920_ _0921_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1331_ mod.cpu.ctrl.o_ibus_adr\[2\] _0861_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1262_ mod.u_scanchain_local.module_data_in\[38\] mod.cpu.bufreg2.dat\[7\] _0823_
+ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_81 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_70 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_92 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1193_ _0766_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1625__C1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1529_ _0258_ _0260_ _0263_ _0259_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1631__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2151__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1603__I _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2434__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1622__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1880_ _0515_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1494__B _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1689__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1314_ _0652_ mod.u_scanchain_local.module_data_in\[61\] _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1245_ mod.cpu.bufreg2.i_dat\[27\] _0812_ _0790_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1513__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1176_ _0753_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2174__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1423__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2047__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1333__I _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1030_ _0625_ mod.cpu.alu.add_cy_r _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2197__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ _0550_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1863_ _0495_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1794_ mod.cpu.csr_imm _0252_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1228_ _0667_ _0797_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1159_ _0686_ _0684_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1770__A1 mod.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1761__A1 mod.cpu.bufreg2.i_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _0191_ net3 mod.cpu.bufreg.data\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2131_ _0122_ net3 mod.cpu.bufreg2.dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1063__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2062_ _0049_ net4 mod.u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1013_ mod.cpu.bufreg2.i_op_b_sel mod.cpu.bufreg.i_sh_signed _0608_ mod.cpu.branch_op
+ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1915_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ mod.cpu.bufreg.data\[10\] mod.cpu.bufreg.data\[11\] _0496_ _0497_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2212__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1777_ _0782_ _0447_ _0758_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1238__I mod.cpu.bufreg2.i_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1052__I0 mod.cpu.bufreg2.i_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1807__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2235__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1259__S _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1700_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1631_ _0247_ _0330_ _0343_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1562_ _0810_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1493_ _0859_ mod.cpu.ctrl.pc_plus_offset_cy_r _0706_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2114_ _0105_ net3 mod.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2045_ _0031_ net4 mod.u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1829_ mod.cpu.bufreg.data\[3\] mod.cpu.bufreg.data\[4\] _0485_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1725__A1 mod.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2108__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2258__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1716__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_132 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_110 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_121 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_154 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_143 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_165 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_176 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1341__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1652__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1497__B _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1255__I0 mod.cpu.bufreg2.i_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1707__A1 mod.cpu.bufreg2.i_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ _0320_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1516__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1545_ _0253_ _0273_ _0274_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1476_ mod.cpu.ctrl.o_ibus_adr\[31\] _0972_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1251__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2028_ _0012_ net4 mod.cpu.bufreg2.i_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1643__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1174__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2080__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1330_ mod.u_scanchain_local.module_data_in\[65\] _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1261_ _0816_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_71 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_60 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_93 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1192_ mod.cpu.bufreg2.dat\[4\] _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xtiny_user_project_82 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1071__I mod.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1625__B1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__C2 mod.cpu.bufreg2.dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1528_ _0627_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1459_ mod.cpu.ctrl.o_ibus_adr\[27\] _0956_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1616__B1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1092__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1147__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1066__I _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1313_ mod.cpu.bufreg2.dat\[30\] _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1244_ mod.cpu.bufreg2.dat\[1\] _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1175_ mod.cpu.bufreg2.i_dat\[17\] mod.cpu.immdec.imm11_7\[4\] _0643_ _0753_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1614__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1931_ mod.cpu.ctrl.o_ibus_adr\[8\] _0546_ _0549_ mod.cpu.ctrl.o_ibus_adr\[9\] _0550_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1862_ _0505_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0461_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2141__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1227_ _0799_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1158_ mod.cpu.immdec.imm11_7\[1\] mod.cpu.immdec.imm11_7\[2\] mod.cpu.immdec.imm11_7\[3\]
+ mod.cpu.immdec.imm11_7\[0\] _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1089_ _0619_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1770__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1522__A2 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2014__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1761__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2164__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2130_ _0121_ net3 mod.cpu.bufreg2.dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1280__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2061_ _0048_ net4 mod.u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1012_ _0606_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ _0250_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1845_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1776_ _0984_ _0682_ _0656_ _0702_ _0436_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1504__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ _0246_ net3 mod.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1203__B _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2037__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2187__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1282__I1 mod.cpu.bufreg2.dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ mod.cpu.bufreg2.dat\[11\] _0296_ _0333_ mod.cpu.bufreg2.dat\[12\] _0343_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1561_ _0770_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ _0987_ _0993_ _0996_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1498__A1 mod.cpu.bufreg2.i_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2113_ _0104_ net3 mod.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2044_ _0029_ net4 mod.u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1273__I1 mod.cpu.bufreg2.dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1828_ _0486_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1973__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1759_ _0432_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1489__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1661__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1264__I1 mod.cpu.bufreg2.dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1823__S _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_111 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_133 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_100 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_122 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_155 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_144 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_166 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_177 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2202__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A1 mod.cpu.bufreg2.i_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1613_ _0324_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1544_ _0679_ mod.cpu.state.o_cnt\[2\] _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1475_ mod.u_scanchain_local.module_data_in\[94\] _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2027_ _0011_ net4 mod.cpu.bufreg2.i_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1643__A1 mod.cpu.bufreg2.i_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2225__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1260_ _0822_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_50 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1191_ mod.cpu.bufreg2.dat\[0\] mod.cpu.bufreg2.dat\[1\] mod.cpu.bufreg2.dat\[2\]
+ mod.cpu.bufreg2.dat\[3\] _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_61 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_72 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_83 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_94 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1625__B2 mod.cpu.bufreg2.dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__A1 mod.cpu.bufreg2.i_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2248__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1527_ _0668_ _0670_ _0261_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1458_ mod.u_scanchain_local.module_data_in\[90\] _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1389_ _0794_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1616__A1 mod.cpu.bufreg2.dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1616__B2 mod.cpu.bufreg2.dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1083__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1312_ _0851_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1243_ _0811_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1174_ _0751_ _0748_ _0752_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1720__I _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2093__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1930_ _0535_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1861_ mod.cpu.bufreg.data\[17\] mod.cpu.bufreg.data\[18\] _0501_ _0505_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1792_ mod.cpu.immdec.imm19_12_20\[2\] _0460_ _0449_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1226_ mod.cpu.bufreg2.i_dat\[22\] _0738_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1157_ _0603_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1088_ mod.cpu.state.init_done _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1842__I1 mod.cpu.bufreg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1770__A3 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1450__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1833__I1 mod.cpu.bufreg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _0047_ net4 mod.u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1011_ mod.cpu.bne_or_bge _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1913_ _0538_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1985__B1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1844_ _0692_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1775_ _0444_ _0445_ _0446_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2258_ _0245_ net3 mod.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1209_ mod.cpu.bufreg2.i_dat\[19\] _0749_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1270__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2189_ _0180_ net3 mod.cpu.bufreg.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1203__C _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2131__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1560_ _0682_ _0676_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ _0994_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1291__S _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1498__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2112_ _0103_ net3 mod.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2043_ _0028_ net4 mod.u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__C1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1827_ mod.cpu.bufreg.data\[2\] mod.cpu.bufreg.data\[3\] _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1186__A1 mod.cpu.bufreg2.i_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1758_ mod.cpu.bufreg2.i_dat\[29\] _0431_ _0425_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1689_ mod.cpu.bufreg2.i_dat\[2\] _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1214__B _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1661__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_123 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_112 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_101 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_134 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_145 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_156 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_178 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_167 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1286__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1612_ _0291_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1543_ _0679_ mod.cpu.state.o_cnt\[2\] _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ _0755_ _0978_ _0979_ _0980_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2027__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ _0010_ net4 mod.cpu.bufreg2.i_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__C1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2177__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1643__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_40 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_73 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_51 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_62 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1190_ mod.cpu.bufreg2.dat\[5\] _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xtiny_user_project_84 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_95 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1744__S _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1526_ _0656_ mod.cpu.bne_or_bge _0676_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1457_ _0959_ _0964_ _0965_ _0967_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1388_ mod.cpu.ctrl.o_ibus_adr\[13\] _0907_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2009_ mod.cpu.bufreg2.i_dat\[11\] _0380_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1543__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1311_ mod.u_scanchain_local.module_data_in\[60\] mod.cpu.bufreg2.dat\[29\] _0781_
+ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1242_ mod.cpu.bufreg2.i_dat\[26\] _0810_ _0790_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1173_ mod.cpu.bufreg2.i_dat\[16\] _0749_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2215__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1782__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1534__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1509_ mod.cpu.bufreg2.i_dat\[11\] _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1183__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2238__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1300__I1 mod.cpu.bufreg2.dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _0504_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _0391_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1764__A1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1225_ _0797_ _0722_ _0728_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1156_ _0690_ _0689_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1087_ _0656_ mod.cpu.bufreg2.dat\[5\] _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ mod.cpu.ctrl.o_ibus_adr\[31\] _0251_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1178__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1842__S _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1010_ mod.cpu.decode.co_mem_word _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__B1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1289__S _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1912_ mod.cpu.ctrl.o_ibus_adr\[1\] _0251_ _0536_ mod.cpu.ctrl.o_ibus_adr\[2\] _0538_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1843_ _0494_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1774_ _0605_ _0435_ _0388_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1752__S _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2257_ _0244_ net3 mod.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1208_ _0673_ _0781_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2188_ _0179_ net3 mod.cpu.bufreg.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1139_ _0718_ _0721_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1728__A1 mod.cpu.bufreg2.i_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2083__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ mod.cpu.state.stage_two_req _0672_ _0678_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1742__I1 mod.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2111_ _0102_ net3 mod.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ _0027_ net4 mod.u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1655__B1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1826_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1757_ mod.cpu.immdec.imm30_25\[5\] mod.cpu.immdec.imm30_25\[4\] _0418_ _0431_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1186__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1688_ _0376_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_113 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_102 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_124 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_157 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_146 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_135 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_179 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_168 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ _0772_ _0327_ _0329_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1366__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1542_ _0272_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ mod.cpu.bufreg.data\[30\] _0788_ _0648_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2025_ _0009_ net4 mod.cpu.bufreg2.i_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__C2 mod.cpu.bufreg2.dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1809_ _0451_ _0472_ _0473_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1225__B _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2121__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1570__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__I _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_41 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_30 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_74 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_63 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_85 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_96 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1525_ _0659_ _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1456_ mod.cpu.bufreg.data\[26\] _0962_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2144__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1387_ mod.u_scanchain_local.module_data_in\[76\] _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2008_ mod.cpu.immdec.imm11_7\[4\] _0761_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1077__A1 mod.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1068__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2017__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2167__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1310_ _0850_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1241_ mod.cpu.bufreg2.dat\[0\] _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1172_ mod.cpu.immdec.imm11_7\[3\] _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1231__A1 mod.cpu.bufreg2.i_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__S _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1508_ _1005_ _1002_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1439_ mod.cpu.ctrl.o_ibus_adr\[23\] _0940_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1470__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1222__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1773__A2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1836__I0 mod.cpu.bufreg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1790_ mod.cpu.immdec.imm19_12_20\[3\] _0252_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1374__I _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1224_ mod.cpu.bufreg.lsb\[0\] _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1155_ _0728_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1086_ _0657_ _0666_ _0669_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1827__I0 mod.cpu.bufreg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1988_ _0584_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1143__B _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1682__A1 mod.cpu.bufreg2.i_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1682__B2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1369__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1911_ _0537_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1842_ mod.cpu.bufreg.data\[9\] mod.cpu.bufreg.data\[10\] _0490_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1773_ mod.cpu.immdec.imm7 _0783_ _0421_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1037__I1 mod.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2256_ _0243_ net3 mod.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1207_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2187_ _0178_ net3 mod.cpu.bufreg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1673__A1 mod.cpu.bufreg2.dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1138_ mod.cpu.bufreg2.dat\[0\] mod.cpu.bufreg2.dat\[8\] mod.cpu.bufreg2.dat\[16\]
+ mod.cpu.bufreg2.dat\[24\] mod.cpu.bufreg.lsb\[0\] _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1069_ mod.cpu.bufreg2.i_dat\[5\] _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1279__I _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2228__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1664__A1 mod.cpu.bufreg2.dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2110_ _0101_ net3 mod.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2041_ _0026_ net4 mod.cpu.bufreg2.i_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1655__B2 mod.cpu.bufreg2.dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1655__A1 mod.cpu.bufreg2.i_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1825_ _0692_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1756_ _0430_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1687_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2239_ _0227_ net3 mod.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__B2 mod.cpu.bufreg2.dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1646__A1 mod.cpu.bufreg2.i_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2050__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_103 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_114 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_136 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_147 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_125 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_158 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_169 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ mod.cpu.bufreg2.i_dat\[5\] _0293_ _0328_ _0766_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1573__B1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1541_ _0673_ _0254_ _0105_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1472_ mod.cpu.ctrl.o_ibus_adr\[30\] _0972_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1382__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2024_ _0007_ net4 mod.cpu.bufreg2.i_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__A1 mod.cpu.bufreg2.i_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1628__B2 mod.cpu.bufreg2.dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1758__S _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2073__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1808_ mod.cpu.immdec.imm19_12_20\[6\] _0457_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1739_ _0725_ _0699_ _0704_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1619__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1890__I1 mod.cpu.bufreg.data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_31 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_20 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_75 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_42 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_64 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_53 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_86 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_97 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2096__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1524_ _0657_ _0718_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1455_ _0647_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1386_ _0877_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ _1005_ _0379_ _0598_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1776__B1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1925__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1240_ _0808_ _0649_ _0801_ _0809_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1171_ _0747_ _0748_ _0750_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_8 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__A1 mod.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1231__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1835__I _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1507_ mod.cpu.bufreg2.i_dat\[10\] _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1438_ mod.u_scanchain_local.module_data_in\[86\] _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1369_ _0794_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1222__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1773__A3 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2134__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1223_ _0792_ _0738_ _0796_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1154_ mod.cpu.bufreg2.i_dat\[7\] _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1085_ _0625_ _0665_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1987_ mod.cpu.ctrl.o_ibus_adr\[30\] _0539_ _0581_ mod.cpu.ctrl.o_ibus_adr\[31\]
+ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1676__C1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1140__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2157__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1131__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1910_ _0859_ _0251_ _0536_ mod.cpu.ctrl.o_ibus_adr\[1\] _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1841_ _0493_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1772_ mod.cpu.bufreg2.i_dat\[7\] _0433_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1334__B _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2255_ _0242_ net3 mod.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2186_ _0177_ net3 mod.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1206_ _0681_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1137_ mod.cpu.bufreg.lsb\[1\] _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1673__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1068_ _0645_ _0649_ _0653_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1425__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1189__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1664__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1416__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0025_ net4 mod.cpu.bufreg2.i_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1655__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ _0483_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1755_ mod.cpu.bufreg2.i_dat\[28\] _0429_ _0425_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1686_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2238_ _0226_ net3 mod.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1646__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ _0160_ net3 mod.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1334__A1 mod.cpu.bufreg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_104 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_115 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_126 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_137 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_148 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_159 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1540_ _0271_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1573__A1 mod.cpu.bufreg2.i_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ mod.u_scanchain_local.module_data_in\[93\] _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2023_ _0006_ net4 mod.cpu.bufreg2.i_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2218__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1807_ mod.cpu.bufreg2.i_dat\[17\] _0433_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1738_ _0402_ _0415_ _0416_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1669_ mod.cpu.bufreg2.i_dat\[25\] _0293_ _0355_ mod.cpu.bufreg2.dat\[25\] _0359_
+ mod.cpu.bufreg2.dat\[26\] _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1619__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_21 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_32 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_10 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_43 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_54 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_65 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_98 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_87 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_76 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1523_ mod.cpu.state.o_cnt_r\[0\] _0730_ mod.cpu.alu.cmp_r _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1454_ mod.cpu.ctrl.o_ibus_adr\[26\] _0956_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1385_ _0894_ _0906_ _0908_ _0909_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2006_ mod.cpu.immdec.imm11_7\[4\] _0592_ _0597_ _0403_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2040__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2190__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1776__A1 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1170_ mod.cpu.bufreg2.i_dat\[15\] _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2063__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_9 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1767__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1519__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1506_ _1004_ _1002_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1437_ _0943_ _0948_ _0949_ _0951_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1368_ mod.cpu.ctrl.o_ibus_adr\[9\] _0891_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1299_ _0844_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1222__A3 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2086__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1222_ _0703_ _0793_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1153_ _0654_ _0649_ _0696_ _0736_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1084_ _0667_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1986_ _0583_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1676__C2 mod.cpu.bufreg2.dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1676__B1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1903__A1 mod.cpu.bufreg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1667__B1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2101__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1440__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ mod.cpu.bufreg.data\[8\] mod.cpu.bufreg.data\[9\] _0490_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2251__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ _0434_ _0442_ _0443_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2254_ _0000_ net3 mod.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1658__B1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2185_ _0176_ net3 mod.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1205_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1136_ _0607_ _0720_ _0709_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1122__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1350__B _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1067_ mod.cpu.bufreg2.i_dat\[3\] _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1189__A2 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1969_ _0573_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1649__B1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2124__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1823_ mod.cpu.alu.cmp_r _0264_ _0605_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1754_ mod.cpu.immdec.imm30_25\[4\] mod.cpu.immdec.imm30_25\[3\] _0418_ _0429_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1718__I1 mod.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1343__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2237_ _0225_ net3 mod.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2168_ _0159_ net3 mod.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1119_ _0683_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2099_ _0090_ net4 mod.u_scanchain_local.module_data_in\[94\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1300__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1334__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_105 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_138 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_116 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_127 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_149 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1022__A1 mod.cpu.bufreg2.i_op_b_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1470_ _0755_ _0975_ _0976_ _0977_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1325__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2022_ _0005_ net4 mod.cpu.bufreg2.i_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1806_ mod.cpu.immdec.imm19_12_20\[7\] _0424_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1013__A1 mod.cpu.bufreg2.i_op_b_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ mod.cpu.immdec.imm24_20\[4\] _0406_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1854__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1668_ _0804_ _0298_ _0367_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1599_ _0288_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_11 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_22 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_44 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_33 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_55 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_66 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_88 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_99 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_77 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1875__S _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1522_ mod.cpu.ctrl.i_jump _0254_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1453_ mod.u_scanchain_local.module_data_in\[89\] _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1384_ mod.cpu.bufreg.data\[12\] _0897_ _0901_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2005_ _0751_ _0592_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1482__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1785__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1767__A2 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1519__A2 _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1505_ mod.cpu.bufreg2.i_dat\[9\] _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1436_ mod.cpu.bufreg.data\[22\] _0946_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1367_ mod.u_scanchain_local.module_data_in\[72\] _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1298_ mod.u_scanchain_local.module_data_in\[54\] mod.cpu.bufreg2.dat\[23\] _0843_
+ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1446__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2030__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2180__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1221_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1152_ _0700_ _0717_ _0101_ _0727_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1083_ _0625_ _0665_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1437__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1985_ mod.cpu.ctrl.o_ibus_adr\[29\] _0578_ _0581_ mod.cpu.ctrl.o_ibus_adr\[30\]
+ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1912__A2 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1419_ mod.cpu.ctrl.o_ibus_adr\[19\] _0924_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1676__A1 mod.cpu.bufreg2.i_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1676__B2 mod.cpu.bufreg2.dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1140__A3 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2053__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1667__A1 mod.cpu.bufreg2.dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__B2 mod.cpu.bufreg2.dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1770_ mod.cpu.immdec.imm30_25\[5\] _0388_ _0419_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2253_ _0241_ net3 mod.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1658__A1 mod.cpu.bufreg2.i_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2184_ _0175_ net3 mod.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1204_ _0629_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1135_ mod.cpu.mem_bytecnt\[0\] _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1066_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2076__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1968_ mod.cpu.ctrl.o_ibus_adr\[22\] _0572_ _0569_ mod.cpu.ctrl.o_ibus_adr\[23\]
+ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1899_ _0602_ _0730_ _0764_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 mod.cpu.bufreg2.i_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A1 mod.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1451__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2099__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1822_ _0434_ _0482_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1753_ _0428_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1684_ _0639_ _0757_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2236_ _0224_ net3 mod.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2167_ _0158_ net3 mod.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1788__S _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1118_ mod.cpu.bufreg2.i_op_b_sel _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2098_ _0089_ net4 mod.u_scanchain_local.module_data_in\[93\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1049_ mod.u_arbiter.i_wb_cpu_ack _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1803__A1 mod.cpu.bufreg2.i_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_106 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_117 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_139 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_128 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2241__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2021_ _0092_ net4 mod.cpu.bufreg2.i_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1805_ _0450_ _0469_ _0470_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2114__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ mod.cpu.bufreg2.i_dat\[24\] _0378_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1013__A2 mod.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1667_ mod.cpu.bufreg2.dat\[24\] _0296_ _0337_ mod.cpu.bufreg2.dat\[25\] _0367_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1598_ _0819_ _0767_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2219_ _0209_ net3 mod.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1311__S _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_23 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1780__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_12 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_56 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_34 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_45 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_89 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_78 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_67 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2137__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1521_ _0251_ _0255_ _0256_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1452_ _0959_ _0960_ _0961_ _0963_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1383_ mod.cpu.ctrl.o_ibus_adr\[12\] _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2004_ _1004_ _0393_ _0596_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1719_ _0401_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1170__A1 mod.cpu.bufreg2.i_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1473__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1225__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1216__S _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1161__A1 mod.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1504_ _1003_ _1002_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1435_ _0647_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1152__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1366_ _0877_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1297_ _0780_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1796__S _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1143__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1757__I0 mod.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1220_ _0774_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1151_ _0728_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1082_ mod.cpu.bne_or_bge _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _0582_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1373__A1 mod.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1418_ mod.u_scanchain_local.module_data_in\[82\] _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1125__A1 mod.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1676__A2 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1349_ _0794_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1600__A2 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1667__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1355__A1 mod.cpu.bufreg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2252_ _0240_ net3 mod.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1203_ _0655_ _0773_ _0777_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2183_ _0174_ net3 mod.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1658__A2 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1134_ mod.cpu.mem_if.signbit _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1065_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1967_ _0558_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1898_ _0527_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1649__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2020__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1821__A2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2170__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1812__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1821_ mod.cpu.bufreg.i_sh_signed _0388_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1752_ mod.cpu.bufreg2.i_dat\[27\] _0427_ _0425_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1576__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1683_ _0854_ _0325_ _0375_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2235_ _0223_ net3 mod.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2166_ _0157_ net3 mod.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2043__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1117_ _0675_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2097_ _0088_ net4 mod.u_scanchain_local.module_data_in\[92\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1048_ _0638_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1817__B _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1309__S _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_107 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_118 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_129 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2066__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2020_ _0085_ net4 mod.cpu.bufreg2.i_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1688__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1804_ mod.cpu.immdec.imm19_12_20\[5\] _0457_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1735_ mod.cpu.immdec.imm30_25\[0\] _0387_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ _0365_ _0366_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1597_ _0317_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2218_ _0208_ net3 mod.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2149_ _0140_ net3 mod.cpu.bufreg2.dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2089__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_13 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_46 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1712__A1 mod.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_24 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_57 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_35 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_68 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_79 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1520_ mod.cpu.state.ibus_cyc _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1451_ mod.cpu.bufreg.data\[25\] _0962_ _0950_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1382_ _0860_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1703__A1 mod.cpu.bufreg2.i_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2003_ mod.cpu.immdec.imm11_7\[2\] _0591_ _0595_ _0761_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2231__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1242__I0 mod.cpu.bufreg2.i_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1718_ _0399_ mod.cpu.immdec.imm24_20\[0\] _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1649_ mod.cpu.bufreg2.i_dat\[17\] _0347_ _0355_ mod.cpu.bufreg2.dat\[17\] _0344_
+ mod.cpu.bufreg2.dat\[18\] _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__I _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1170__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1630__B1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1933__B2 mod.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2104__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2254__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ mod.cpu.bufreg2.i_dat\[8\] _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1434_ mod.cpu.ctrl.o_ibus_adr\[22\] _0940_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1365_ _0878_ _0890_ _0892_ _0893_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1296_ _0842_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2127__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1560__B _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1052__S _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1150_ _0726_ _0729_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1081_ _0661_ _0634_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1897__S _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1693__I0 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1983_ mod.cpu.ctrl.o_ibus_adr\[28\] _0578_ _0581_ mod.cpu.ctrl.o_ibus_adr\[29\]
+ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1417_ _0927_ _0932_ _0933_ _0935_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1348_ mod.cpu.ctrl.o_ibus_adr\[5\] _0874_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1279_ _0816_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1047__S _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2251_ _0239_ net3 mod.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1202_ _0729_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2182_ _0173_ net3 mod.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1133_ _0676_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1064_ _0646_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _0571_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1897_ mod.cpu.bufreg.data\[31\] _0526_ _0484_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1820_ _0481_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1025__A1 mod.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1751_ mod.cpu.immdec.imm30_25\[3\] mod.cpu.immdec.imm30_25\[2\] _0418_ _0427_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1682_ mod.cpu.bufreg2.i_dat\[31\] _0291_ _0327_ _0665_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1328__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2234_ _0222_ net3 mod.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2165_ _0156_ net3 mod.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1116_ _0683_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2096_ _0087_ net4 mod.u_scanchain_local.module_data_in\[91\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1047_ mod.cpu.i_timer_irq mod.cpu.immdec.imm24_20\[4\] _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1949_ mod.cpu.ctrl.o_ibus_adr\[15\] _0559_ _0555_ mod.cpu.ctrl.o_ibus_adr\[16\]
+ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1319__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_108 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_119 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1558__A2 mod.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1034__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1803_ mod.cpu.bufreg2.i_dat\[16\] _0383_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1734_ _0402_ _0412_ _0413_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ mod.cpu.bufreg2.i_dat\[23\] _0336_ _0331_ mod.cpu.bufreg2.dat\[23\] _0366_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1596_ mod.cpu.bufreg2.i_dat\[3\] _0298_ _0316_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2160__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ _0001_ net3 mod.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2148_ _0139_ net3 mod.cpu.bufreg2.dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2079_ _0068_ net4 mod.u_scanchain_local.module_data_in\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_14 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_115_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_36 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_25 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_47 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_58 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_69 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1228__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2033__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ _0787_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2183__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1381_ mod.u_scanchain_local.module_data_in\[75\] _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1473__B _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _0751_ _0592_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1699__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1482__A4 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1717_ _0726_ _0702_ _0386_ _0376_ _0604_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1648_ _0295_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1579_ _0300_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1402__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2056__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__A1 mod.cpu.bufreg2.dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1630__B2 mod.cpu.bufreg2.dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1502_ _1001_ _1002_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1433_ mod.u_scanchain_local.module_data_in\[85\] _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1364_ mod.cpu.bufreg.data\[8\] _0881_ _0885_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1295_ mod.u_scanchain_local.module_data_in\[53\] mod.cpu.bufreg2.dat\[22\] _0838_
+ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2079__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1892__I _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1080_ _0623_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1693__I1 mod.cpu.bufreg2.i_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1982_ _0562_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1416_ mod.cpu.bufreg.data\[18\] _0930_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1347_ mod.u_scanchain_local.module_data_in\[68\] _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1278_ _0832_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2010__A1 mod.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2244__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2250_ _0238_ net3 mod.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1201_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _0172_ net3 mod.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1132_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1063_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1815__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2117__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1965_ mod.cpu.ctrl.o_ibus_adr\[21\] _0566_ _0569_ mod.cpu.ctrl.o_ibus_adr\[22\]
+ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1896_ _0524_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1410__I _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1320__I _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1750_ _0426_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0852_ _0325_ _0321_ _0854_ _0374_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2233_ _0221_ net3 mod.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2164_ _0155_ net3 mod.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1115_ _0698_ _0699_ _0684_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ _0086_ net4 mod.u_scanchain_local.module_data_in\[90\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1046_ _0630_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1948_ _0560_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1879_ mod.cpu.bufreg.data\[25\] mod.cpu.bufreg.data\[26\] _0511_ _0515_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_109 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1191__A1 mod.cpu.bufreg2.dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1802_ mod.cpu.immdec.imm19_12_20\[6\] _0424_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1733_ mod.cpu.immdec.imm24_20\[3\] _0406_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ mod.cpu.bufreg2.dat\[24\] _0321_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1595_ _0303_ _0313_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0207_ net3 mod.cpu.bufreg.data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2147_ _0138_ net3 mod.cpu.bufreg2.dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2078_ _0067_ net4 mod.u_scanchain_local.module_data_in\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1029_ mod.cpu.alu.i_rs1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1173__A1 mod.cpu.bufreg2.i_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_15 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_26 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_37 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1135__I mod.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_48 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_59 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ _0894_ _0903_ _0904_ _0905_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2001_ _1003_ _0762_ _0594_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1716_ _0395_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1647_ _0353_ _0354_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1578_ mod.cpu.bufreg2.dat\[0\] _0812_ _0285_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1630__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1697__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2150__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1501_ _0781_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1432_ _0943_ _0944_ _0945_ _0947_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1363_ mod.cpu.ctrl.o_ibus_adr\[8\] _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1294_ _0841_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1503__I mod.cpu.bufreg2.i_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1128__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2023__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2173__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1323__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1981_ _0580_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1415_ _0647_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2046__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1346_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1530__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1277_ mod.u_scanchain_local.module_data_in\[45\] mod.cpu.bufreg2.dat\[14\] _0828_
+ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1233__I mod.cpu.bufreg2.i_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2196__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2010__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1521__A1 _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2109__CLKN net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1588__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2001__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2069__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2180_ _0171_ net3 mod.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1200_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1131_ _0663_ _0714_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1062_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1964_ _0570_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1895_ mod.cpu.bufreg.i_sh_signed mod.cpu.bufreg.data\[31\] _0522_ _0525_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1329_ _0863_ _0864_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1806__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2211__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1042__I0 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1582__B _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1601__I _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1680_ mod.cpu.bufreg2.i_dat\[30\] _0303_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2232_ _0220_ net3 mod.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2163_ _0154_ net3 mod.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1114_ _0675_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2094_ _0084_ net4 mod.u_scanchain_local.module_data_in\[89\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1045_ _0636_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2234__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1947_ mod.cpu.ctrl.o_ibus_adr\[14\] _0559_ _0555_ mod.cpu.ctrl.o_ibus_adr\[15\]
+ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ _0514_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1660__B1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1715__A1 mod.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2107__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ _0450_ _0466_ _0467_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1732_ mod.cpu.bufreg2.i_dat\[23\] _0378_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _0364_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1706__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ _0819_ _0771_ _0300_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1309__I1 mod.cpu.bufreg2.dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _0206_ net3 mod.cpu.bufreg.data\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0137_ net3 mod.cpu.bufreg2.dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1241__I mod.cpu.bufreg2.dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2077_ _0066_ net4 mod.u_scanchain_local.module_data_in\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1028_ _0609_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1245__I0 mod.cpu.bufreg2.i_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_27 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1173__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_16 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_38 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_49 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1936__A1 mod.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2000_ mod.cpu.immdec.imm11_7\[1\] _0591_ _0593_ _0761_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1715_ mod.cpu.immdec.imm24_20\[1\] _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1646_ mod.cpu.bufreg2.i_dat\[16\] _0323_ _0351_ mod.cpu.bufreg2.dat\[16\] _0354_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1577_ _0284_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2129_ _0120_ net3 mod.cpu.bufreg2.dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1606__B1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1257__S _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ mod.cpu.bufreg2.i_dat\[6\] _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1056__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1431_ mod.cpu.bufreg.data\[21\] _0946_ _0934_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1362_ _0860_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1293_ mod.u_scanchain_local.module_data_in\[52\] mod.cpu.bufreg2.dat\[21\] _0838_
+ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1629_ _0342_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1128__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1119__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ mod.cpu.ctrl.o_ibus_adr\[27\] _0578_ _0575_ mod.cpu.ctrl.o_ibus_adr\[28\]
+ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1414_ mod.cpu.ctrl.o_ibus_adr\[18\] _0924_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1345_ _0650_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1276_ _0831_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2140__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1130_ _0708_ _0713_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1061_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1963_ mod.cpu.ctrl.o_ibus_adr\[20\] _0566_ _0569_ mod.cpu.ctrl.o_ibus_adr\[21\]
+ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0989_ _0992_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1509__I mod.cpu.bufreg2.i_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2013__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2163__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1328_ mod.cpu.ctrl.o_ibus_adr\[1\] _0793_ _0861_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1259_ mod.u_scanchain_local.module_data_in\[37\] mod.cpu.bufreg2.dat\[6\] _0817_
+ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1154__I mod.cpu.bufreg2.i_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2186__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2231_ _0219_ net3 mod.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2100__D _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2162_ _0153_ net3 mod.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1113_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2093_ _0083_ net4 mod.u_scanchain_local.module_data_in\[88\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1044_ mod.cpu.i_rf_ready mod.cpu.immdec.imm24_20\[3\] _0631_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1877_ mod.cpu.bufreg.data\[24\] mod.cpu.bufreg.data\[25\] _0511_ _0514_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2059__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1660__A1 mod.cpu.bufreg2.dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1660__B2 mod.cpu.bufreg2.dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1715__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1612__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1651__A1 mod.cpu.bufreg2.dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ mod.cpu.csr_imm _0451_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1731_ mod.cpu.immdec.imm24_20\[4\] _0387_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ mod.cpu.bufreg2.i_dat\[22\] _0347_ _0355_ mod.cpu.bufreg2.dat\[22\] _0359_
+ mod.cpu.bufreg2.dat\[23\] _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__1706__A2 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1593_ _0771_ _0767_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2214_ _0205_ net3 mod.cpu.bufreg.data\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2145_ _0136_ net3 mod.cpu.bufreg2.dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2201__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2076_ _0065_ net4 mod.u_scanchain_local.module_data_in\[71\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1027_ mod.cpu.bufreg2.i_rs2 _0622_ _0613_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1929_ _0548_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_17 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_28 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_39 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__A1 mod.cpu.bufreg2.i_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1633__B2 mod.cpu.bufreg2.dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2224__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1714_ _0760_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1718__S _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1645_ mod.cpu.bufreg2.dat\[17\] _0349_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1576_ _0814_ _0288_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1163__I0 mod.cpu.bufreg2.i_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2128_ _0119_ net3 mod.cpu.bufreg2.dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2059_ _0046_ net4 mod.u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1427__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2247__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__B1 mod.cpu.i_rf_ready vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1606__A1 mod.cpu.bufreg2.i_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1430_ _0787_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1361_ mod.u_scanchain_local.module_data_in\[71\] _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1292_ _0840_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1072__I _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1628_ mod.cpu.bufreg2.i_dat\[10\] _0339_ _0341_ mod.cpu.bufreg2.dat\[10\] _0337_
+ mod.cpu.bufreg2.dat\[11\] _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1559_ _0603_ _0281_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2004__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1413_ mod.u_scanchain_local.module_data_in\[81\] _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1344_ _0855_ _0873_ _0875_ _0876_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1275_ mod.u_scanchain_local.module_data_in\[44\] mod.cpu.bufreg2.dat\[13\] _0828_
+ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1818__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2092__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1615__I _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1060_ net2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1962_ _0562_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1893_ _0989_ _0992_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1327_ _0857_ mod.u_scanchain_local.module_data_in\[64\] _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1258_ _0821_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1189_ _0612_ _0764_ _0677_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1019__A2 mod.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1435__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1194__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2230_ _0218_ net3 mod.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2161_ _0152_ net3 mod.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1112_ mod.cpu.decode.opcode\[0\] _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2092_ _0082_ net4 mod.u_scanchain_local.module_data_in\[87\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1043_ _0635_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1013__C mod.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1945_ _0250_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1876_ _0513_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2130__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1660__A2 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1651__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2153__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1730_ _0402_ _0409_ _0410_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1661_ _0792_ _0330_ _0363_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1592_ mod.cpu.bufreg2.dat\[3\] _0309_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2213_ _0204_ net3 mod.cpu.bufreg.data\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2144_ _0135_ net3 mod.cpu.bufreg2.dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2075_ _0064_ net4 mod.u_scanchain_local.module_data_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1026_ _0612_ _0615_ _0618_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1928_ mod.cpu.ctrl.o_ibus_adr\[7\] _0546_ _0543_ mod.cpu.ctrl.o_ibus_adr\[8\] _0548_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1859_ mod.cpu.bufreg.data\[16\] mod.cpu.bufreg.data\[17\] _0501_ _0504_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1158__A1 mod.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_18 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_29 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2026__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2176__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1321__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1713_ _0395_ _0396_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1644_ _0350_ _0352_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ _0290_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2049__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1163__I1 mod.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2199__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2127_ _0118_ net3 mod.cpu.bufreg2.dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2058_ _0045_ net4 mod.u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1009_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1708__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__B2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1443__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1606__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1819__S _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1360_ _0878_ _0887_ _0888_ _0889_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1291_ mod.u_scanchain_local.module_data_in\[51\] mod.cpu.bufreg2.dat\[20\] _0838_
+ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1627_ _0295_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1558_ mod.cpu.mem_bytecnt\[1\] mod.cpu.bufreg.lsb\[1\] _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1489_ _0782_ _0691_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1772__A1 mod.cpu.bufreg2.i_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1284__S _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ _0927_ _0928_ _0929_ _0931_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1343_ mod.cpu.bufreg.data\[4\] _0795_ _0868_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1274_ _0830_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2237__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1054__I0 mod.cpu.bufreg2.i_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1506__A1 _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1993__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1168__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1681__B1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _0568_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0764_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1736__A1 mod.cpu.bufreg2.i_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1742__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1326_ _0858_ _0862_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1257_ mod.cpu.bufreg2.i_dat\[31\] _0766_ _0817_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1188_ _0739_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2082__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _0151_ net3 mod.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1111_ _0655_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2091_ _0081_ net4 mod.u_scanchain_local.module_data_in\[86\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1042_ _0634_ mod.cpu.immdec.imm24_20\[2\] _0631_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2109__D mod.u_scanchain_local.module_data_in\[95\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1257__I0 mod.cpu.bufreg2.i_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1944_ _0557_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ mod.cpu.bufreg.data\[23\] mod.cpu.bufreg.data\[24\] _0511_ _0513_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1709__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1309_ mod.u_scanchain_local.module_data_in\[59\] mod.cpu.bufreg2.dat\[28\] _0781_
+ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1248__I0 mod.cpu.bufreg2.i_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1660_ mod.cpu.bufreg2.dat\[21\] _0296_ _0333_ mod.cpu.bufreg2.dat\[22\] _0363_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1591_ _0312_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2212_ _0203_ net3 mod.cpu.bufreg.data\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2143_ _0134_ net3 mod.cpu.bufreg2.dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ _0062_ net4 mod.u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1025_ mod.cpu.bufreg2.i_cnt_done mod.cpu.immdec.imm31 _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1927_ _0547_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1858_ _0503_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1789_ _0458_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_19 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1618__B1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1109__C _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1840__S _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2120__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1712_ mod.cpu.decode.co_ebreak _0393_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1643_ mod.cpu.bufreg2.i_dat\[15\] _0323_ _0351_ mod.cpu.bufreg2.dat\[15\] _0352_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1574_ _0287_ _0292_ _0297_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2126_ _0117_ net3 mod.cpu.bufreg2.dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2057_ _0044_ net4 mod.u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1008_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1724__I _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1551__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2143__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1067__A1 mod.cpu.bufreg2.i_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1290_ _0839_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2016__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1230__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1781__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1626_ _0340_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2166__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1557_ mod.cpu.mem_bytecnt\[1\] mod.cpu.bufreg.lsb\[1\] mod.cpu.bufreg.lsb\[0\] mod.cpu.mem_bytecnt\[0\]
+ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1488_ _0989_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ mod.u_scanchain_local.module_data_in\[95\] net4 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1772__A2 _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1524__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2039__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2189__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1763__A2 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1411_ mod.cpu.bufreg.data\[17\] _0930_ _0917_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1342_ mod.cpu.ctrl.o_ibus_adr\[4\] _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1273_ mod.u_scanchain_local.module_data_in\[43\] mod.cpu.bufreg2.dat\[12\] _0828_
+ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1506__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1609_ _0295_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1690__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1293__I1 mod.cpu.bufreg2.dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1184__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1960_ mod.cpu.ctrl.o_ibus_adr\[19\] _0566_ _0563_ mod.cpu.ctrl.o_ibus_adr\[20\]
+ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1891_ _0521_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1295__S _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1325_ _0859_ _0793_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2204__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1256_ _0820_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1187_ _0755_ _0762_ _0763_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_91_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1027__I1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1266__I1 mod.cpu.bufreg2.dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1179__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2227__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1642__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1110_ _0660_ _0694_ _0687_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2090_ _0080_ net4 mod.u_scanchain_local.module_data_in\[85\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1041_ _0625_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1089__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1943_ mod.cpu.ctrl.o_ibus_adr\[13\] _0552_ _0555_ mod.cpu.ctrl.o_ibus_adr\[14\]
+ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1874_ _0512_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1308_ _0849_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1239_ _0667_ _0797_ _0806_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1248__I1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1838__S _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1590_ mod.cpu.bufreg2.i_dat\[2\] _0298_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1175__I0 mod.cpu.bufreg2.i_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _0202_ net3 mod.cpu.bufreg.data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2142_ _0133_ net3 mod.cpu.bufreg2.dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2073_ _0061_ net4 mod.u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1024_ _0619_ mod.cpu.branch_op mod.cpu.csr_d_sel _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1926_ mod.cpu.ctrl.o_ibus_adr\[6\] _0546_ _0543_ mod.cpu.ctrl.o_ibus_adr\[7\] _0547_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1857_ mod.cpu.bufreg.data\[15\] mod.cpu.bufreg.data\[16\] _0501_ _0503_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1788_ mod.cpu.immdec.imm19_12_20\[1\] _0456_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__B _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1618__A1 mod.cpu.bufreg2.dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1618__B2 mod.cpu.bufreg2.dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2072__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1085__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1711_ mod.cpu.bufreg2.i_dat\[20\] _0377_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1642_ _0324_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1573_ mod.cpu.bufreg2.i_dat\[0\] _0293_ _0296_ _0810_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2125_ _0116_ net3 mod.cpu.bufreg2.dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2056_ _0043_ net4 mod.u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1007_ mod.cpu.state.o_cnt_r\[3\] mod.cpu.state.o_cnt_r\[2\] _0602_ _0603_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2095__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1909_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1226__B _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1067__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1915__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1298__S _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1625_ mod.cpu.bufreg2.i_dat\[9\] _0339_ _0328_ mod.cpu.bufreg2.dat\[9\] _0337_ mod.cpu.bufreg2.dat\[10\]
+ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__1825__I _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1556_ _0280_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1487_ _0699_ _0622_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2108_ _0100_ net3 mod.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2039_ _0024_ net4 mod.cpu.bufreg2.i_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2110__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1460__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ _0787_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1341_ _0860_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1272_ _0829_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1451__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1987__B1 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2133__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1608_ _0290_ _0300_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1539_ _0709_ _0710_ _0112_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_59_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1690__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1681__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2156__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1890_ mod.cpu.bufreg.data\[30\] mod.cpu.bufreg.data\[31\] _0484_ _0521_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1197__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1744__I0 mod.cpu.bufreg2.i_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1324_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1255_ mod.cpu.bufreg2.i_dat\[30\] _0819_ _0817_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1186_ mod.cpu.bufreg2.i_dat\[18\] _0749_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1672__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2029__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2179__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1195__I _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1040_ _0633_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1103__A1 mod.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1942_ _0556_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1873_ mod.cpu.bufreg.data\[22\] mod.cpu.bufreg.data\[23\] _0511_ _0512_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1590__A1 mod.cpu.bufreg2.i_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1307_ mod.u_scanchain_local.module_data_in\[58\] mod.cpu.bufreg2.dat\[27\] _0843_
+ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1238_ mod.cpu.bufreg2.i_dat\[25\] _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1645__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1169_ _0651_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1899__B _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0201_ net3 mod.cpu.bufreg.data\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1175__I1 mod.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2141_ _0132_ net3 mod.cpu.bufreg2.dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2072_ _0060_ net4 mod.u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1023_ mod.cpu.decode.opcode\[2\] _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1925_ _0539_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1856_ _0502_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1787_ _0448_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1158__A4 mod.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1563__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2217__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1710_ _0392_ _0394_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1641_ mod.cpu.bufreg2.dat\[16\] _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1572_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1545__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2124_ _0115_ net3 mod.cpu.bufreg2.dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2055_ _0042_ net4 mod.u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1006_ mod.cpu.state.o_cnt_r\[0\] mod.cpu.state.o_cnt_r\[1\] _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1908_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1784__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1839_ _0492_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1311__I1 mod.cpu.bufreg2.dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput5 net5 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1138__S0 mod.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1302__I1 mod.cpu.bufreg2.dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2007__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1766__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1624_ _0777_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1518__A1 _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1555_ _0269_ mod.cpu.state.o_cnt_r\[1\] _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1486_ _0701_ _0663_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2062__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2107_ _0099_ net4 mod.cpu.bufreg2.i_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2038_ _0023_ net4 mod.cpu.bufreg2.i_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1057__I0 mod.cpu.bufreg2.i_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2085__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1340_ mod.u_scanchain_local.module_data_in\[67\] _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1271_ mod.u_scanchain_local.module_data_in\[42\] mod.cpu.bufreg2.dat\[11\] _0828_
+ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1607_ _0322_ _0326_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1538_ _0270_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1469_ mod.cpu.bufreg.data\[29\] _0788_ _0966_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1197__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1323_ _0757_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1254_ mod.cpu.bufreg2.dat\[4\] _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1185_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2100__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2250__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1941_ mod.cpu.ctrl.o_ibus_adr\[12\] _0552_ _0555_ mod.cpu.ctrl.o_ibus_adr\[13\]
+ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1872_ _0495_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1386__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1306_ _0847_ _0748_ _0848_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1237_ _0804_ _0649_ _0807_ _0801_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1168_ _0648_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1099_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2146__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1021__A1 mod.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2140_ _0131_ net3 mod.cpu.bufreg2.dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _0059_ net4 mod.u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1022_ mod.cpu.bufreg2.i_op_b_sel _0617_ mod.cpu.immdec.imm24_20\[0\] _0618_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1602__C _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2019__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ _0545_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1855_ mod.cpu.bufreg.data\[14\] mod.cpu.bufreg.data\[15\] _0501_ _0502_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1786_ _0390_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__I _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1315__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1306__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1640_ _0332_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1571_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2123_ _0114_ net3 mod.cpu.bufreg2.dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2054_ _0040_ net4 mod.u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1481__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1907_ _0249_ _0740_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1838_ mod.cpu.bufreg.data\[7\] mod.cpu.bufreg.data\[8\] _0490_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1769_ _0403_ _0419_ _0440_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput6 net6 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1138__S1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1623_ _0338_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1518__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1394__I _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1554_ _0279_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1485_ _0725_ _0616_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2207__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

