* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12902__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09671_ _03868_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08622_ _02053_ _02928_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14966__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08553_ _01949_ _02859_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09287__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12130__I1 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07504_ _01787_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08484_ _02041_ mod.u_cpu.rf_ram.memory\[356\]\[1\] _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12830__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07435_ _01560_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07366_ mod.u_cpu.rf_ram.memory\[388\]\[0\] mod.u_cpu.rf_ram.memory\[389\]\[0\] mod.u_cpu.rf_ram.memory\[390\]\[0\]
+ mod.u_cpu.rf_ram.memory\[391\]\[0\] _01673_ _01666_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_176_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09105_ net2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _01604_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14346__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09036_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _03259_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08014__A2 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14496__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13146__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09938_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13846__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11029__B _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09869_ _04001_ mod.u_cpu.rf_ram.memory\[538\]\[0\] _04020_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11900_ _05415_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14120__S _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12880_ _06076_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11831_ _05365_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14550_ _00404_ net3 mod.u_cpu.rf_ram.memory\[412\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10132__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _05318_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13501_ _06559_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15121__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10713_ _04172_ _04570_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14023__A1 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14481_ _00335_ net3 mod.u_cpu.rf_ram.memory\[447\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12575__S _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11693_ _05271_ mod.u_cpu.rf_ram.memory\[251\]\[1\] _05269_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13432_ _03508_ _06511_ _06514_ _03507_ _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10644_ _04556_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13363_ _06458_ _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10575_ _04498_ mod.u_cpu.rf_ram.memory\[430\]\[1\] _04508_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15271__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15102_ _00956_ net3 mod.u_cpu.rf_ram.memory\[489\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12314_ _03696_ _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13294_ _06281_ _06284_ _06391_ _06392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14839__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15033_ _00887_ net3 mod.u_cpu.rf_ram.memory\[201\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__S _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12245_ _05635_ mod.u_cpu.rf_ram.memory\[196\]\[1\] _05646_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12176_ _05600_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10899__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13137__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11127_ _04847_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13837__A1 _06340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14989__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _03984_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10009_ _04115_ mod.u_cpu.rf_ram.memory\[516\]\[1\] _04113_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10371__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14817_ _00671_ net3 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11453__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14748_ _00602_ net3 mod.u_cpu.rf_ram.memory\[313\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11871__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14679_ _00533_ net3 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14369__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _01527_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15614__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07151_ _01439_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09441__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12328__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09744__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13128__I0 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11628__I _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13828__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ _02124_ _02282_ _02290_ _02291_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09723_ _03711_ _03788_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07507__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09654_ _03854_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07841__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08605_ _01738_ _02874_ _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_76_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15144__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09585_ _03763_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _02730_ _02842_ _02207_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07366__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08467_ _02303_ mod.u_cpu.rf_ram.memory\[374\]\[1\] _02773_ _01867_ _02774_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15294__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07418_ _01605_ _01725_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08398_ _02500_ mod.u_cpu.rf_ram.memory\[436\]\[1\] _02704_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13603__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _01532_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11614__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10707__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _04364_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09019_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _03324_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10291_ _04313_ mod.u_cpu.rf_ram.memory\[476\]\[1\] _04316_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10643__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12030_ _05498_ mod.u_cpu.rf_ram.memory\[19\]\[0\] _05503_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13819__A1 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13981_ _06946_ _06948_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09499__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11474__S _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12932_ _06110_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12863_ _05786_ _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13047__A2 _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08068__B _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14602_ _00456_ net3 mod.u_cpu.rf_ram.memory\[386\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11814_ _05354_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14511__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15582_ _01353_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _06019_ mod.u_cpu.rf_ram.memory\[130\]\[1\] _06015_ _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15637__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14533_ _00387_ net3 mod.u_cpu.rf_ram.memory\[421\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _05265_ _05306_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__S _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__I1 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14464_ _00318_ net3 mod.u_cpu.rf_ram.memory\[455\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11676_ _05243_ mod.u_cpu.rf_ram.memory\[256\]\[0\] _05259_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12558__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10408__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13415_ _06354_ mod.u_cpu.rf_ram.memory\[139\]\[1\] _06503_ _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14661__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08515__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10627_ _04546_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14395_ _00249_ net3 mod.u_cpu.rf_ram.memory\[490\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09423__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11230__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13346_ _06424_ _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10558_ _04498_ mod.u_cpu.rf_ram.memory\[433\]\[1\] _04494_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11649__S _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13277_ _06321_ _06373_ _06374_ _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10489_ _04452_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15017__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15016_ _00870_ net3 mod.u_cpu.rf_ram.memory\[207\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09726__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12030__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12228_ _05636_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07737__A1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12159_ _03727_ _04379_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10592__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15167__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13286__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__I0 mod.u_cpu.rf_ram.memory\[288\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13530__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08162__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09370_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _02592_ _02620_ _02627_ _01658_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11844__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11911__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08252_ _02559_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07203_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08425__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08183_ _02321_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _01438_ _01441_ _01442_ _01443_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10024__A2 _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11772__A2 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07728__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12721__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07967_ _02272_ mod.u_cpu.rf_ram.memory\[254\]\[0\] _02274_ _02252_ _02275_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13277__A2 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__11288__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14534__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07898_ _02202_ _02203_ _02205_ _02049_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07571__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09637_ _03779_ _03820_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__A1 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ _03704_ _03747_ _03748_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__B1 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12788__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ mod.u_cpu.rf_ram.memory\[341\]\[1\] _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14684__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11835__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ mod.u_cpu.cpu.immdec.imm11_7\[3\] mod.u_cpu.cpu.immdec.imm11_7\[4\] _03724_
+ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10263__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11530_ _05161_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08335__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__A2 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09405__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ _05113_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08839__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13200_ _06283_ _06285_ _06296_ _06306_ _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10412_ _04347_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14180_ _07081_ mod.u_cpu.rf_ram.memory\[8\]\[1\] _07083_ _07085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11392_ _05046_ mod.u_cpu.rf_ram.memory\[300\]\[0\] _05067_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07967__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13131_ _06255_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12960__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10343_ _04302_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07746__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12012__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10274_ _04305_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13062_ mod.u_cpu.rf_ram.memory\[69\]\[1\] _06005_ _06209_ _06211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__C _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11268__I _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _05492_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11279__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10326__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13964_ _06920_ _06934_ _06935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09192__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09341__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12915_ _04955_ _04644_ _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13895_ _06581_ mod.u_cpu.rf_ram.memory\[112\]\[1\] _06882_ _06884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14217__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15634_ _01405_ net3 mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12846_ _03743_ _06052_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13976__B1 _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15565_ _01336_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12777_ _05992_ mod.u_cpu.rf_ram.memory\[132\]\[0\] _06007_ _06008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14516_ _00370_ net3 mod.u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11728_ _05295_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15496_ _01267_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14447_ _00301_ net3 mod.u_cpu.rf_ram.memory\[464\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11659_ _04973_ _05120_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14378_ _00232_ net3 mod.u_cpu.rf_ram.memory\[498\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14407__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12951__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13329_ _06425_ _06402_ _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10801__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08870_ mod.u_cpu.rf_ram.memory\[552\]\[1\] mod.u_cpu.rf_ram.memory\[553\]\[1\] mod.u_cpu.rf_ram.memory\[554\]\[1\]
+ mod.u_cpu.rf_ram.memory\[555\]\[1\] _02472_ _02473_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14557__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08383__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07821_ _02047_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15525__D _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10810__I _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ mod.u_cpu.rf_ram.memory\[148\]\[0\] mod.u_cpu.rf_ram.memory\[149\]\[0\] mod.u_cpu.rf_ram.memory\[150\]\[0\]
+ mod.u_cpu.rf_ram.memory\[151\]\[0\] _02059_ _01723_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07605__B _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09183__I0 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07683_ _01850_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14208__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _03650_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _03415_ mod.u_scanchain_local.module_data_in\[56\] _03408_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\]
+ _03596_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11817__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10458__S _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08304_ _02350_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11442__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _03521_
+ _03532_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__07110__A2 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ _01855_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13195__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08950__I _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08166_ mod.u_cpu.rf_ram.memory\[552\]\[0\] mod.u_cpu.rf_ram.memory\[553\]\[0\] mod.u_cpu.rf_ram.memory\[554\]\[0\]
+ mod.u_cpu.rf_ram.memory\[555\]\[0\] _02472_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12942__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15332__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11745__A2 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07117_ mod.u_cpu.cpu.decode.op26 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08097_ _02154_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08374__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15482__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10181__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08999_ _03301_ _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10961_ _04746_ _04770_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__A2 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12700_ _05938_ mod.u_cpu.rf_ram.memory\[140\]\[1\] _05956_ _05958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10484__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13680_ _06689_ _06690_ _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10892_ _04724_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12631_ _05870_ _03886_ _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11808__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12647__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08429__A2 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13422__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15350_ _01125_ net3 mod.u_cpu.rf_ram.memory\[369\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12562_ _05865_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14301_ _00155_ net3 mod.u_cpu.rf_ram.memory\[537\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11513_ _05144_ mod.u_cpu.rf_ram.memory\[281\]\[0\] _05150_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15281_ _00039_ net4 mod.u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12493_ _05821_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14232_ _00086_ net3 mod.u_cpu.rf_ram.memory\[571\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11444_ _05101_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11036__I1 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__S1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13478__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14163_ _06062_ _06568_ _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _01968_ _05055_ _05056_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09892__S _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13114_ _06244_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ _04330_ mod.u_cpu.rf_ram.memory\[470\]\[1\] _04339_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14094_ _07029_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13045_ _06199_ mod.u_cpu.rf_ram.memory\[107\]\[1\] _06197_ _06200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10257_ _04292_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A2 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10188_ _04217_ mod.u_cpu.rf_ram.memory\[490\]\[0\] _04243_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14996_ _00850_ net3 mod.u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13110__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13947_ _03430_ _03433_ _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08668__A2 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13661__A2 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15205__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13878_ _06422_ _06864_ _06866_ _06811_ _06870_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_15617_ _01388_ net3 mod.u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12829_ _06042_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12472__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15548_ _01319_ net3 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15355__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10077__I _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15479_ _01251_ net3 mod.u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08020_ _02297_ mod.u_cpu.rf_ram.memory\[116\]\[0\] _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09971_ _03762_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07319__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08922_ _02527_ mod.u_cpu.rf_ram.memory\[540\]\[1\] _03228_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10538__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08853_ _01608_ mod.u_cpu.rf_ram.memory\[38\]\[1\] _03159_ _02212_ _03160_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10163__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10540__I _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07804_ mod.u_cpu.rf_ram.memory\[173\]\[0\] _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08784_ mod.u_cpu.rf_ram.memory\[84\]\[1\] mod.u_cpu.rf_ram.memory\[85\]\[1\] mod.u_cpu.rf_ram.memory\[86\]\[1\]
+ mod.u_cpu.rf_ram.memory\[87\]\[1\] _01857_ _02054_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09305__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07735_ _02042_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07666_ _01956_ _01959_ _01973_ _01812_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09405_ _03439_ mod.u_scanchain_local.module_data_in\[64\] _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13404__A2 _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07597_ _01875_ mod.u_cpu.rf_ram.memory\[356\]\[0\] _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09336_ _03578_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13800__B _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09267_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08831__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14722__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _02084_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09198_ _03471_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12915__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08149_ _01634_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07296__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12391__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11160_ _04896_ mod.u_cpu.rf_ram.memory\[337\]\[1\] _04907_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14872__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11747__S _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _04178_ mod.u_cpu.rf_ram.memory\[501\]\[1\] _04185_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11091_ _04796_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10042_ _01612_ _04138_ _04139_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09217__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13891__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14850_ _00704_ net3 mod.u_cpu.rf_ram.memory\[262\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15228__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09147__I0 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13801_ _06789_ _06774_ _06800_ _06801_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14140__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14781_ _00635_ net3 mod.u_cpu.rf_ram.memory\[297\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11993_ _05470_ mod.u_cpu.rf_ram.memory\[569\]\[0\] _05478_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13732_ _06722_ _06657_ _06737_ _06738_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_17_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10944_ _04758_ _04759_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11654__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14252__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15378__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10098__S _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13663_ _06661_ _06369_ _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _04703_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15402_ _01177_ net3 mod.u_cpu.rf_ram.memory\[359\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12614_ _05283_ _05900_ _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08791__S _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13594_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] mod.u_arbiter.i_wb_cpu_dbus_adr\[30\]
+ _06614_ _06618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15333_ _01108_ net3 mod.u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12545_ _05854_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15264_ _00021_ net4 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12476_ _02535_ _05809_ _05810_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14215_ _03735_ mod.u_cpu.rf_ram.memory\[259\]\[1\] _07103_ _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11427_ _05071_ mod.u_cpu.rf_ram.memory\[294\]\[0\] _05090_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15195_ _01048_ net3 mod.u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08586__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14146_ _07062_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11358_ _05044_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13936__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10309_ _04266_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14077_ _03910_ _04996_ _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11289_ _01921_ _04997_ _04998_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07934__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13331__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12134__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13331__B2 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13028_ _06184_ mod.u_cpu.rf_ram.memory\[84\]\[1\] _06187_ _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11456__I _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10940__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11392__S _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14979_ _00833_ net3 mod.u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07520_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A1 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07451_ _01758_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07602__C _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14745__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07382_ mod.u_cpu.rf_ram.memory\[396\]\[0\] mod.u_cpu.rf_ram.memory\[397\]\[0\] mod.u_cpu.rf_ram.memory\[398\]\[0\]
+ mod.u_cpu.rf_ram.memory\[399\]\[0\] _01689_ _01683_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09121_ _03419_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11948__A2 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09596__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09052_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08433__C _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08003_ _02105_ _02292_ _02310_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14895__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10384__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ _02547_ _04078_ _04079_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08329__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13322__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07844__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _02500_ _03211_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13322__B2 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09885_ _04018_ mod.u_cpu.rf_ram.memory\[536\]\[1\] _04030_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10136__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13873__A2 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10270__I _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ mod.u_cpu.rf_ram.memory\[48\]\[1\] mod.u_cpu.rf_ram.memory\[49\]\[1\] mod.u_cpu.rf_ram.memory\[50\]\[1\]
+ mod.u_cpu.rf_ram.memory\[51\]\[1\] _02421_ _02393_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14275__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08767_ _02303_ _03073_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15520__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08188__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ _01757_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11636__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08698_ mod.u_cpu.rf_ram.memory\[199\]\[1\] _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13514__C _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07935__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _01919_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10660_ _04560_ mod.u_cpu.rf_ram.memory\[416\]\[1\] _04565_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11239__I1 mod.u_cpu.rf_ram.memory\[324\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__A2 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _03497_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _04520_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14118__S _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08804__A2 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13022__S _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08360__S0 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12330_ _05705_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__C _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12261_ _05645_ mod.u_cpu.rf_ram.memory\[193\]\[0\] _05658_ _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14000_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _06954_ _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08112__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11212_ _04943_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput7 net7 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_12192_ _05334_ _05611_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07240__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11143_ _04897_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15050__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13313__A1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12116__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11074_ _04841_ mod.u_cpu.rf_ram.memory\[351\]\[1\] _04849_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14618__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10180__I _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10025_ mod.u_cpu.rf_ram.memory\[513\]\[0\] _03925_ _04126_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12911__I1 mod.u_cpu.rf_ram.memory\[399\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14902_ _00756_ net3 mod.u_cpu.rf_ram.memory\[233\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08740__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14833_ _00687_ net3 mod.u_cpu.rf_ram.memory\[271\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15623__D _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13616__A2 _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14764_ _00618_ net3 mod.u_cpu.rf_ram.memory\[305\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12675__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14768__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11976_ _02458_ _05466_ _05467_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13715_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10927_ _04739_ mod.u_cpu.rf_ram.memory\[373\]\[1\] _04745_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14695_ _00549_ net3 mod.u_cpu.rf_ram.memory\[340\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13646_ _06655_ _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10858_ _03990_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_158_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12835__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13577_ _06608_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10789_ _04641_ mod.u_cpu.rf_ram.memory\[395\]\[1\] _04652_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15316_ mod.u_cpu.cpu.o_wdata1 net3 mod.u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12528_ _01574_ _05842_ _05844_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10602__A2 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15247_ _00052_ net4 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12459_ _03338_ _03668_ _03359_ _03394_ _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12771__S _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08559__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15178_ _01031_ net3 mod.u_cpu.rf_ram.memory\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09220__A2 mod.u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13666__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14129_ _07051_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07664__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12107__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14298__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11186__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15543__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10090__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _03847_ mod.u_cpu.rf_ram.memory\[561\]\[0\] _03867_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08731__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08621_ mod.u_cpu.rf_ram.memory\[140\]\[1\] mod.u_cpu.rf_ram.memory\[141\]\[1\] mod.u_cpu.rf_ram.memory\[142\]\[1\]
+ mod.u_cpu.rf_ram.memory\[143\]\[1\] _02070_ _02071_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08709__B _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08552_ mod.u_cpu.rf_ram.memory\[319\]\[1\] _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07503_ _01773_ _01805_ _01810_ _01785_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ _01520_ _02789_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ _01741_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14032__A2 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09104_ _03403_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13791__A1 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07296_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09035_ _03338_ mod.u_cpu.cpu.genblk3.csr.mcause31 _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15073__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09598__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12480__I _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07574__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A1 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04066_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13846__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09868_ _03797_ _04003_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09770__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14910__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08819_ mod.u_cpu.rf_ram.memory\[31\]\[1\] _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11830_ _05364_ mod.u_cpu.rf_ram.memory\[39\]\[1\] _05362_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _05304_ mod.u_cpu.rf_ram.memory\[239\]\[1\] _05316_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13500_ _03642_ _06557_ _06558_ _03648_ _06559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10712_ _04602_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14480_ _00334_ net3 mod.u_cpu.rf_ram.memory\[447\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _05249_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13431_ _06516_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10643_ mod.u_cpu.rf_ram.memory\[41\]\[1\] _04532_ _04554_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12034__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08789__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07749__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15416__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13362_ _06391_ _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _04509_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10596__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15101_ _00955_ net3 mod.u_cpu.rf_ram.memory\[175\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08073__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12313_ _05693_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07461__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13293_ mod.u_arbiter.i_wb_cpu_rdt\[9\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _03499_ _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15032_ _00886_ net3 mod.u_cpu.rf_ram.memory\[201\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12244_ _05647_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14440__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15566__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12175_ _05583_ mod.u_cpu.rf_ram.memory\[76\]\[1\] _05598_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10899__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11126_ _04886_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11057_ _04837_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11848__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12896__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14590__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10008_ _04090_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14816_ _00670_ net3 mod.u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08248__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11959_ _05442_ mod.u_cpu.rf_ram.memory\[529\]\[0\] _05456_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14747_ _00601_ net3 mod.u_cpu.rf_ram.memory\[314\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14678_ _00532_ net3 mod.u_cpu.rf_ram.memory\[348\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13629_ _06332_ _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13073__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15096__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07150_ _01458_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12820__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09441__A2 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12328__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07394__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13128__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14933__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ _01533_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09722_ _03908_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08004__I0 mod.u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08704__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ _03832_ mod.u_cpu.rf_ram.memory\[563\]\[1\] _03852_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08604_ _01977_ _02893_ _02910_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09584_ _03799_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12639__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09114__I _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08158__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08535_ mod.u_cpu.rf_ram.memory\[296\]\[1\] mod.u_cpu.rf_ram.memory\[297\]\[1\] mod.u_cpu.rf_ram.memory\[298\]\[1\]
+ mod.u_cpu.rf_ram.memory\[299\]\[1\] _01753_ _01916_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11311__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14313__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15439__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _01864_ _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07417_ mod.u_cpu.rf_ram.memory\[405\]\[0\] _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08397_ _02111_ _02703_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07348_ _01483_ _01590_ _01655_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10578__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14463__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15589__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13516__A1 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ _03259_ _03322_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ _04317_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10750__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13819__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13980_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06938_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _06948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A2 mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12931_ _06105_ mod.u_cpu.rf_ram.memory\[369\]\[1\] _06108_ _06110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11554__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12862_ _06062_ _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11813_ _05350_ mod.u_cpu.rf_ram.memory\[49\]\[1\] _05352_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14601_ _00455_ net3 mod.u_cpu.rf_ram.memory\[387\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08068__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15581_ _01352_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12793_ _06018_ _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14532_ _00386_ net3 mod.u_cpu.rf_ram.memory\[421\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11744_ _04983_ _03823_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12007__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14463_ _00317_ net3 mod.u_cpu.rf_ram.memory\[456\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13055__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07682__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14806__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11675_ _04838_ _05120_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07700__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07479__I mod.u_cpu.raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12558__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13414_ _06504_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _04523_ mod.u_cpu.rf_ram.memory\[422\]\[0\] _04545_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14394_ _00248_ net3 mod.u_cpu.rf_ram.memory\[490\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12802__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13345_ _06441_ _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10557_ _04497_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11230__A2 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09694__I _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14956__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13276_ _06300_ _06374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10488_ _04247_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11369__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15015_ _00869_ net3 mod.u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12227_ _05635_ mod.u_cpu.rf_ram.memory\[119\]\[1\] _05632_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12030__I1 mod.u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A2 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12158_ _03712_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08103__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11109_ _04864_ mod.u_cpu.rf_ram.memory\[345\]\[0\] _04874_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12869__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12089_ _05533_ mod.u_cpu.rf_ram.memory\[65\]\[1\] _05540_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__I1 mod.u_cpu.rf_ram.memory\[289\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08162__A2 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14336__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09111__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08320_ _02611_ _02623_ _02626_ _01742_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14486__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _01757_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07389__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _01509_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13746__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _02476_ _02482_ _02488_ _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _01427_ _01432_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07425__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11221__A2 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08722__B _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14171__A1 _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10032__I0 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__I _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09973__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12721__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08013__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15111__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11780__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08948__I _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07966_ _02180_ _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09705_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07897_ _02204_ mod.u_cpu.rf_ram.memory\[216\]\[0\] _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11532__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _03840_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08784__S0 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15261__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09567_ _03785_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12237__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14829__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09102__A1 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__B2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12788__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ mod.u_cpu.rf_ram.memory\[336\]\[1\] mod.u_cpu.rf_ram.memory\[337\]\[1\] mod.u_cpu.rf_ram.memory\[338\]\[1\]
+ mod.u_cpu.rf_ram.memory\[339\]\[1\] _01841_ _01844_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09498_ _01441_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08616__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _02337_ _02755_ _01591_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13037__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13588__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14979__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11460_ _05108_ mod.u_cpu.rf_ram.memory\[28\]\[1\] _05111_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08839__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _04399_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11391_ _04784_ _05058_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13130_ mod.u_arbiter.i_wb_cpu_rdt\[17\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _06253_ _06255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07967__A2 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12960__A2 _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10342_ _03850_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14162__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13061_ _02353_ _06209_ _06210_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10273_ _04298_ mod.u_cpu.rf_ram.memory\[478\]\[0\] _04304_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12012_ _05470_ mod.u_cpu.rf_ram.memory\[57\]\[0\] _05491_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14359__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15604__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13963_ _03444_ _05794_ _06934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10326__I1 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11284__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11523__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09341__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12914_ _06098_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13894_ _06883_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14217__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12845_ _01478_ _06052_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15633_ _01404_ net3 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13205__S _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13976__A1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07711__B _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15564_ _01335_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13976__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12776_ _03960_ _05978_ _06007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14515_ _00369_ net3 mod.u_cpu.rf_ram.memory\[430\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13028__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11727_ _05289_ mod.u_cpu.rf_ram.memory\[242\]\[0\] _05294_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15495_ _01266_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14446_ _00300_ net3 mod.u_cpu.rf_ram.memory\[464\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _05246_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10609_ _04533_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07407__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14377_ _00231_ net3 mod.u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11589_ _05199_ mod.u_cpu.rf_ram.memory\[268\]\[0\] _05200_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13328_ _06298_ _06304_ _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12951__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15134__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13259_ _05787_ _06356_ _06357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10014__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13900__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10714__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11395__S _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08383__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ mod.u_cpu.rf_ram.memory\[160\]\[0\] mod.u_cpu.rf_ram.memory\[161\]\[0\] mod.u_cpu.rf_ram.memory\[162\]\[0\]
+ mod.u_cpu.rf_ram.memory\[163\]\[0\] _02125_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15284__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07751_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12467__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07605__C _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08135__A2 _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07682_ _01979_ _01980_ _01988_ _01989_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09421_ _03496_ mod.u_scanchain_local.module_data_in\[67\] _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _03593_ _03595_ _03488_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08303_ mod.u_cpu.rf_ram.memory\[472\]\[1\] mod.u_cpu.rf_ram.memory\[473\]\[1\] mod.u_cpu.rf_ram.memory\[474\]\[1\]
+ mod.u_cpu.rf_ram.memory\[475\]\[1\] _02593_ _02454_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07646__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13019__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _03528_ _03534_ _03537_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08234_ _01688_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08165_ _02388_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12753__I _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07847__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ mod.u_cpu.cpu.decode.op21 _01420_ _01424_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08071__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08096_ mod.u_cpu.rf_ram.memory\[16\]\[0\] mod.u_cpu.rf_ram.memory\[17\]\[0\] mod.u_cpu.rf_ram.memory\[18\]\[0\]
+ mod.u_cpu.rf_ram.memory\[19\]\[0\] _02403_ _02367_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14144__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14501__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15627__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08998_ _03276_ _03302_ _03261_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10181__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07582__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12458__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07949_ mod.u_cpu.rf_ram.memory\[240\]\[0\] mod.u_cpu.rf_ram.memory\[241\]\[0\] mod.u_cpu.rf_ram.memory\[242\]\[0\]
+ mod.u_cpu.rf_ram.memory\[243\]\[0\] _02242_ _02172_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_47_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14651__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A2 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10960_ _04369_ _04713_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07885__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _03745_ _03820_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10891_ mod.u_cpu.rf_ram.memory\[37\]\[1\] _04661_ _04722_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11832__I _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15007__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12630_ _05911_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12561_ _05858_ mod.u_cpu.rf_ram.memory\[161\]\[1\] _05863_ _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11433__A2 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14300_ _00154_ net3 mod.u_cpu.rf_ram.memory\[537\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11512_ _04873_ _05149_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15280_ _00038_ net4 mod.u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12492_ _05813_ mod.u_cpu.rf_ram.memory\[170\]\[0\] _05820_ _05821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15157__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14231_ _00085_ net3 mod.u_cpu.rf_ram.memory\[572\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11443_ _05096_ mod.u_cpu.rf_ram.memory\[291\]\[0\] _05100_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14162_ _03363_ _06631_ _07072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12933__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _05022_ _05055_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13113_ _06237_ mod.u_cpu.rf_ram.memory\[100\]\[1\] _06242_ _06244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10325_ _04340_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14093_ _07028_ mod.u_cpu.rf_ram.memory\[245\]\[1\] _07025_ _07029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13044_ _06104_ _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10256_ _04276_ mod.u_cpu.rf_ram.memory\[480\]\[0\] _04291_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12697__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10187_ _04242_ _04234_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07425__C _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14995_ _00849_ net3 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13110__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13946_ _06912_ _06920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07876__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13249__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12838__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13877_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _06867_ _06869_ _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15616_ _01387_ net3 mod.u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12828_ _06038_ mod.u_cpu.rf_ram.memory\[125\]\[1\] _06040_ _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09212__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07628__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10358__I _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15547_ _01318_ net3 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12774__S _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12759_ _04668_ _05978_ _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15478_ _01250_ net3 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14429_ _00283_ net3 mod.u_cpu.rf_ram.memory\[473\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12573__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14524__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11983__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ _04089_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08921_ _02528_ _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09928__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14674__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10538__I1 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _02190_ _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07803_ _02047_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08783_ _02051_ _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08108__A2 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07734_ _01499_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07665_ _01961_ _01966_ _01971_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09404_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] _03615_ _03639_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _01759_ _01903_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07619__A1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ _03546_ _03580_ _03581_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09266_ _03506_ _03522_ _03523_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _02454_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09197_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] _03469_
+ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12215__I1 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08148_ _02129_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14117__A1 _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ mod.u_cpu.rf_ram.memory\[0\]\[0\] mod.u_cpu.rf_ram.memory\[1\]\[0\] mod.u_cpu.rf_ram.memory\[2\]\[0\]
+ mod.u_cpu.rf_ram.memory\[3\]\[0\] _02385_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10110_ _01594_ _04185_ _04187_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11090_ _04861_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12679__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10041_ _04044_ _04138_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08201__I _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__C _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13800_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _06772_ _06416_ _06801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14140__I1 mod.u_cpu.rf_ram.memory\[289\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11992_ _03767_ _04026_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14780_ _00634_ net3 mod.u_cpu.rf_ram.memory\[297\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12151__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13731_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _06483_ _06709_ _06738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10943_ _04708_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12851__A1 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13662_ _06434_ _06644_ _06673_ _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10874_ _04712_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15401_ _01176_ net3 mod.u_cpu.rf_ram.memory\[359\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12613_ _05373_ _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13593_ _06617_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09967__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14547__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15332_ _00007_ net3 mod.u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12544_ _05837_ mod.u_cpu.rf_ram.memory\[164\]\[1\] _05852_ _05854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08283__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13489__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08804__C _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15263_ _00020_ net4 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12475_ _05759_ _05809_ _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10217__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11426_ _04812_ _05089_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08035__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14214_ _07104_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15194_ _01047_ net3 mod.u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14697__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14145_ _07057_ mod.u_cpu.rf_ram.memory\[90\]\[0\] _07061_ _07062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08586__A2 _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11357_ _05032_ mod.u_cpu.rf_ram.memory\[306\]\[1\] _05042_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10308_ _04329_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14076_ _07017_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11288_ _04746_ _04997_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11717__I0 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09535__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13027_ _06188_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10239_ _04267_ mod.u_cpu.rf_ram.memory\[483\]\[1\] _04278_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13331__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11342__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09299__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14978_ _00832_ net3 mod.u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12142__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13929_ _06904_ mod.u_cpu.rf_ram.memory\[111\]\[1\] _06901_ _06905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12568__I _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12693__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15322__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07450_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13901__B _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07381_ _01633_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09120_ _03412_ _03415_ _03418_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15472__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13399__I _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09051_ _03307_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08002_ _02293_ _02296_ _02309_ _02122_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08026__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11956__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10384__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09953_ _03899_ _04078_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11647__I _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08904_ mod.u_cpu.rf_ram.memory\[519\]\[1\] _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13322__A2 _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09884_ _04031_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10136__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11184__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09117__I _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08835_ mod.u_cpu.rf_ram.memory\[52\]\[1\] mod.u_cpu.rf_ram.memory\[53\]\[1\] mod.u_cpu.rf_ram.memory\[54\]\[1\]
+ mod.u_cpu.rf_ram.memory\[55\]\[1\] _02151_ _02152_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11583__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ mod.u_cpu.rf_ram.memory\[127\]\[1\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07860__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08188__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07717_ _02022_ mod.u_cpu.rf_ram.memory\[268\]\[0\] _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08697_ _02204_ mod.u_cpu.rf_ram.memory\[196\]\[1\] _03003_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07648_ _01914_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07935__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13389__A2 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13633__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07579_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _03567_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10590_ _04506_ mod.u_cpu.rf_ram.memory\[427\]\[0\] _04519_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08360__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09249_ _03502_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13102__I _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _05657_ _05650_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11211_ _04938_ mod.u_cpu.rf_ram.memory\[328\]\[0\] _04942_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08112__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12191_ _05432_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11142_ _04896_ mod.u_cpu.rf_ram.memory\[340\]\[1\] _04894_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13313__A2 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11073_ _04850_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12372__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09027__I _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _04125_ _04002_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_14901_ _00755_ net3 mod.u_cpu.rf_ram.memory\[234\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15345__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14832_ _00686_ net3 mod.u_cpu.rf_ram.memory\[271\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12388__I _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14763_ _00617_ net3 mod.u_cpu.rf_ram.memory\[306\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11975_ _05322_ _05466_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13714_ _03364_ _06657_ _06720_ _06721_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10686__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10926_ _01876_ _04745_ _04747_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15495__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14694_ _00548_ net3 mod.u_cpu.rf_ram.memory\[340\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13721__B _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13645_ _06656_ _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _04699_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10438__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13576_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] mod.u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _06604_ _06608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10788_ _04653_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15315_ mod.u_cpu.rf_ram_if.wdata1_r\[1\] net3 mod.u_cpu.rf_ram_if.wdata1_r\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08534__C _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12527_ _05843_ _05842_ _05844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_185_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15246_ _00041_ net4 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12458_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _05795_ _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08559__A2 _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ _05078_ _05062_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15177_ _01030_ net3 mod.u_cpu.rf_ram.memory\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12389_ _05745_ mod.u_cpu.rf_ram.memory\[177\]\[1\] _05743_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14128_ _07043_ mod.u_cpu.rf_ram.memory\[118\]\[0\] _07050_ _07051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14059_ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] _07000_ _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07881__S _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08620_ _02046_ _02926_ _02051_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08731__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14712__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08551_ _01962_ mod.u_cpu.rf_ram.memory\[316\]\[1\] _02857_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08709__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07502_ _01807_ mod.u_cpu.rf_ram.memory\[446\]\[0\] _01809_ _01783_ _01810_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10677__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08495__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ mod.u_cpu.rf_ram.memory\[357\]\[1\] _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _01630_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14862__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07364_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09103_ _03261_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14018__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ _01495_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15218__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09034_ mod.u_cpu.cpu.bufreg2.i_cnt_done _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11929__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09598__I1 mod.u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14242__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15368__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10281__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08970__A2 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _03818_ _03883_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09867_ _04019_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14392__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13059__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _02302_ mod.u_cpu.rf_ram.memory\[28\]\[1\] _03124_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09798_ _03967_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12806__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _02611_ _03052_ _03055_ _01680_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10668__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12001__I _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11760_ _02250_ _05316_ _05317_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08030__S0 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08486__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10293__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10711_ _04593_ mod.u_cpu.rf_ram.memory\[408\]\[1\] _04600_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09511__S _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11691_ _05270_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10642_ _04555_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13430_ _03492_ _06511_ _06514_ _03508_ _06516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12034__A2 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08354__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10456__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13361_ _06437_ _06447_ _06453_ _06456_ _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__A2 _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13782__A2 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10573_ _04506_ mod.u_cpu.rf_ram.memory\[430\]\[0\] _04508_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15100_ _00954_ net3 mod.u_cpu.rf_ram.memory\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09450__A3 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12312_ _05692_ mod.u_cpu.rf_ram.memory\[185\]\[1\] _05690_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13292_ _06389_ _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07461__A2 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15031_ _00885_ net3 mod.u_cpu.rf_ram.memory\[202\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12243_ _05645_ mod.u_cpu.rf_ram.memory\[196\]\[0\] _05646_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08410__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12174_ _05599_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11125_ _04880_ mod.u_cpu.rf_ram.memory\[343\]\[1\] _04884_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13298__B2 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09980__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14735__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12345__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11056_ _04825_ mod.u_cpu.rf_ram.memory\[353\]\[1\] _04835_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09210__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10007_ _04114_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14098__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14815_ _00669_ net3 mod.u_cpu.rf_ram.memory\[280\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14885__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14746_ _00600_ net3 mod.u_cpu.rf_ram.memory\[314\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08477__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11958_ _05047_ _04118_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10909_ _04720_ mod.u_cpu.rf_ram.memory\[376\]\[1\] _04734_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14677_ _00531_ net3 mod.u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11889_ _05407_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11750__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13628_ _06640_ _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13773__A2 _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13559_ _06598_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14265__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15510__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15229_ _01082_ net3 mod.u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__A1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07982_ _02283_ _02286_ _02289_ _02141_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _03890_ mod.u_cpu.rf_ram.memory\[556\]\[1\] _03906_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09201__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11839__A2 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11925__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _03853_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08603_ _02898_ _02900_ _02046_ _02909_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09583_ _03740_ mod.u_cpu.rf_ram.memory\[570\]\[0\] _03798_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09504__I1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ _02188_ _02837_ _02840_ _01833_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08468__A1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08465_ mod.u_cpu.rf_ram.memory\[375\]\[1\] _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07416_ mod.u_cpu.rf_ram.memory\[400\]\[0\] mod.u_cpu.rf_ram.memory\[401\]\[0\] mod.u_cpu.rf_ram.memory\[402\]\[0\]
+ mod.u_cpu.rf_ram.memory\[403\]\[0\] _01722_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15040__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ mod.u_cpu.rf_ram.memory\[437\]\[1\] _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14608__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ _01591_ _01620_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10578__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08640__A1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07278_ _01532_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13587__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15190__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09017_ _03320_ mod.u_cpu.cpu.ctrl.i_iscomp _03321_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07585__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14758__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12575__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13819__A3 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ _04055_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09499__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _06109_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12861_ _03338_ _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14600_ _00454_ net3 mod.u_cpu.rf_ram.memory\[387\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11812_ _05353_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15580_ _01351_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12792_ _06017_ _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14531_ _00385_ net3 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10387__S _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _05305_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14462_ _00316_ net3 mod.u_cpu.rf_ram.memory\[456\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _05258_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07682__A2 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14288__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13413_ _06351_ mod.u_cpu.rf_ram.memory\[139\]\[0\] _06503_ _06504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10186__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15533__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10625_ _04262_ _04534_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13755__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14393_ _00247_ net3 mod.u_cpu.rf_ram.memory\[491\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10813__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13344_ _06121_ _06441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10556_ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08631__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10914__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13275_ _06359_ _06360_ _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10487_ _04451_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15014_ _00868_ net3 mod.u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12226_ _05634_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12157_ _05587_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12318__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11108_ _04873_ _04869_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12088_ _05541_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12869__I1 mod.u_cpu.rf_ram.memory\[409\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08537__I2 mod.u_cpu.rf_ram.memory\[290\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11039_ _04825_ mod.u_cpu.rf_ram.memory\[356\]\[1\] _04823_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__I1 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15063__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09151__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09111__A2 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14729_ _00583_ net3 mod.u_cpu.rf_ram.memory\[323\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08250_ _02541_ _02557_ _01447_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07201_ _01506_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10096__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _01717_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _01439_ _01440_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07425__A2 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14900__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14171__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08481__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12309__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07965_ mod.u_cpu.rf_ram.memory\[255\]\[0\] _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09704_ _03702_ _03883_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15406__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ _01993_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11532__I1 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10496__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _03832_ mod.u_cpu.rf_ram.memory\[565\]\[1\] _03838_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08784__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07900__A3 _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ _03764_ mod.u_cpu.rf_ram.memory\[572\]\[1\] _03783_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13434__B2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10248__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14430__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11296__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _02778_ _02823_ _01788_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13985__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15556__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ _03722_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08185__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08448_ _02747_ _02754_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _02561_ _02682_ _02685_ _02080_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ mod.u_cpu.rf_ram.memory\[457\]\[1\] _04383_ _04397_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14580__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11390_ _05066_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10341_ _04351_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10420__A1 _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13060_ _05948_ _06209_ _06210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10272_ _04299_ _04303_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12011_ _04294_ _04026_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15086__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13962_ _06932_ _06933_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13673__A1 _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12913_ _06086_ mod.u_cpu.rf_ram.memory\[399\]\[1\] _06096_ _06098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13893_ _06578_ mod.u_cpu.rf_ram.memory\[112\]\[0\] _06882_ _06883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15632_ _01403_ net3 mod.u_cpu.rf_ram.memory\[244\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12844_ _05788_ _05803_ _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13425__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08807__C _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13976__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15563_ _01334_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12775_ _06006_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11987__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14514_ _00368_ net3 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11726_ _05293_ _05284_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15494_ _01265_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14923__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08852__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14445_ _00299_ net3 mod.u_cpu.rf_ram.memory\[465\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11657_ _05234_ mod.u_cpu.rf_ram.memory\[258\]\[1\] _05244_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12936__B1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10608_ mod.u_cpu.rf_ram.memory\[425\]\[1\] _04532_ _04529_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08604__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14376_ _00230_ net3 mod.u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11588_ _04784_ _05191_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13327_ _06385_ _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10539_ _04485_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13258_ _03390_ _03672_ _06356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13955__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11211__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12209_ _04195_ _04125_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09955__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14303__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _06282_ _06289_ _06295_ _06285_ _06296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15429__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07591__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07750_ _01603_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13664__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12467__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14453__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ _01886_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15579__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09420_ _03623_ _03652_ _03653_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12219__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09351_ _03590_ _03594_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09096__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08302_ _02040_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09282_ _03535_ mod.u_scanchain_local.module_data_in\[45\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08843__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _02523_ _02524_ _02540_ _02469_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_166_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08164_ _02329_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_147_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07115_ _01423_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14026__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08095_ _01856_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14144__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11202__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ mod.u_cpu.rf_ram_if.rdata1 _03248_ mod.u_cpu.rf_ram_if.rtrig1 _03302_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07948_ _01740_ _02241_ _02255_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13655__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07334__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ _02149_ _02169_ _02186_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09618_ _03826_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13407__A1 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12210__S _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07885__A2 mod.u_cpu.rf_ram.memory\[220\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14946__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10890_ _02427_ _04722_ _04723_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09549_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11969__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12560_ _05864_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08834__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11511_ _05124_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12491_ _05334_ _05767_ _05820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14230_ _00084_ net3 mod.u_cpu.rf_ram.memory\[572\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11442_ _04965_ _05089_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14161_ _07067_ mod.u_cpu.cpu.ctrl.i_jump _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11373_ _04369_ _05020_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14326__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08693__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10944__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _04326_ mod.u_cpu.rf_ram.memory\[470\]\[0\] _04339_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13112_ _06243_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14092_ _06903_ _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12146__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _04290_ _04137_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13043_ _06198_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__A1 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08445__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13708__C _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A4 _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14476__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10186_ _03918_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07573__A1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14994_ _00848_ net3 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13945_ _06918_ _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__B _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13876_ _06868_ _06837_ _06869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15615_ _01386_ net3 mod.u_cpu.rf_ram.memory\[289\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12827_ _02313_ _06040_ _06041_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15546_ _01317_ net3 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12758_ _05995_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15101__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10632__A1 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11709_ _05271_ mod.u_cpu.rf_ram.memory\[253\]\[1\] _05280_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15477_ _01249_ net3 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12689_ mod.u_cpu.rf_ram.memory\[77\]\[1\] _05950_ _05947_ _05951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14428_ _00282_ net3 mod.u_cpu.rf_ram.memory\[473\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12385__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08272__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14359_ _00213_ net3 mod.u_cpu.rf_ram.memory\[508\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15251__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13185__I0 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14819__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ mod.u_cpu.rf_ram.memory\[541\]\[1\] _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08436__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07683__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ mod.u_cpu.rf_ram.memory\[39\]\[1\] _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13637__A1 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08782_ mod.u_cpu.rf_ram.memory\[80\]\[1\] mod.u_cpu.rf_ram.memory\[81\]\[1\] mod.u_cpu.rf_ram.memory\[82\]\[1\]
+ mod.u_cpu.rf_ram.memory\[83\]\[1\] _02249_ _02107_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14969__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07733_ _01743_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11499__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07316__A1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12030__S _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07664_ _01686_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ _03614_ _03636_ _03638_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_168_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07595_ mod.u_cpu.rf_ram.memory\[357\]\[0\] _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14062__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__I0 mod.u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ _03554_ mod.u_scanchain_local.module_data_in\[53\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_21_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _03516_ mod.u_scanchain_local.module_data_in\[42\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14349__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08216_ mod.u_cpu.rf_ram.memory\[512\]\[0\] mod.u_cpu.rf_ram.memory\[513\]\[0\] mod.u_cpu.rf_ram.memory\[514\]\[0\]
+ mod.u_cpu.rf_ram.memory\[515\]\[0\] _02494_ _02495_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09196_ _03470_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08182__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10226__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11423__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _02454_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14117__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08078_ _01581_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14499__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10040_ _03991_ _04137_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11991_ _05477_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13730_ _06456_ _06725_ _06728_ _06736_ _06640_ _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_84_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ _03857_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09313__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15124__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13661_ _06309_ _06404_ _06402_ _06673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14053__A1 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10873_ _04698_ mod.u_cpu.rf_ram.memory\[382\]\[1\] _04710_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15400_ _01175_ net3 mod.u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12612_ _05899_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08807__A1 _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09855__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13592_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] mod.u_arbiter.i_wb_cpu_dbus_adr\[29\]
+ _06614_ _06617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15331_ _01107_ net3 mod.u_cpu.rf_ram.memory\[246\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12543_ _05853_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08283__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09480__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15274__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15262_ _00018_ net4 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12474_ _05395_ _04033_ _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14213_ _03699_ mod.u_cpu.rf_ram.memory\[259\]\[0\] _07103_ _07104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10194__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11425_ _04995_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15193_ _01046_ net3 mod.u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08035__A2 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__A1 _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14144_ _03796_ _05397_ _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11356_ _05043_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _04326_ mod.u_cpu.rf_ram.memory\[473\]\[0\] _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14075_ _06904_ mod.u_cpu.rf_ram.memory\[114\]\[1\] _07015_ _07017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07717__B _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11287_ _04994_ _04996_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11717__I1 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09535__A2 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13026_ _06186_ mod.u_cpu.rf_ram.memory\[84\]\[0\] _06187_ _06188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10238_ _04279_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10169_ _04230_ _04229_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14977_ _00831_ net3 mod.u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13928_ _06903_ _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09223__I _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13859_ _06664_ _06851_ _06852_ _06464_ _06853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07380_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15617__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15529_ _01300_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _03250_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _02283_ _02301_ _02307_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14641__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08026__A2 _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11956__I1 mod.u_cpu.rf_ram.memory\[218\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08730__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _03896_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14791__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08903_ _02527_ mod.u_cpu.rf_ram.memory\[516\]\[1\] _03209_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09526__A2 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08302__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09883_ _04023_ mod.u_cpu.rf_ram.memory\[536\]\[0\] _04030_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ _01693_ _03121_ _03140_ _02380_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15147__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ _02297_ mod.u_cpu.rf_ram.memory\[124\]\[1\] _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11663__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07716_ _01729_ _02023_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _03001_ _03002_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10279__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12695__S _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07647_ _01915_ _01945_ _01954_ _01768_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11892__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15297__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ _01532_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13633__I1 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09317_ _03415_ mod.u_scanchain_local.module_data_in\[50\] _03562_ _03566_ _03567_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12494__I _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__A1 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09179_ mod.u_arbiter.i_wb_cpu_rdt\[16\] mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] _03459_
+ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11210_ _04804_ _04926_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11021__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12190_ _05610_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11141_ _04879_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08212__I _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09517__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11072_ _04843_ mod.u_cpu.rf_ram.memory\[351\]\[0\] _04849_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12372__I1 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14900_ _00754_ net3 mod.u_cpu.rf_ram.memory\[234\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10023_ _03979_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14831_ _00685_ net3 mod.u_cpu.rf_ram.memory\[272\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12669__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11088__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14514__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14762_ _00616_ net3 mod.u_cpu.rf_ram.memory\[306\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11974_ _03893_ _04108_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13713_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _06704_ _06471_ _06693_ _06656_ _06721_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10925_ _04746_ _04745_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11883__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14693_ _00547_ net3 mod.u_cpu.rf_ram.memory\[341\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07700__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13644_ _06655_ _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ _04698_ mod.u_cpu.rf_ram.memory\[384\]\[1\] _04696_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12588__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10438__I1 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14664__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10917__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13575_ _06607_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10787_ _04637_ mod.u_cpu.rf_ram.memory\[395\]\[0\] _04652_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07498__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15314_ mod.u_cpu.cpu.o_wen0 net3 mod.u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12526_ _05487_ _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15245_ _00030_ net4 mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12457_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _05794_ _05795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13001__A2 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _03712_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15176_ _01029_ net3 mod.u_cpu.rf_ram.memory\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12388_ _05710_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14127_ _03828_ _05631_ _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11339_ _05031_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14058_ _07003_ _07005_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13009_ _06176_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09154__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08550_ _01934_ _02856_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12815__A2 _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07501_ _01779_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08481_ mod.u_cpu.rf_ram.memory\[352\]\[1\] mod.u_cpu.rf_ram.memory\[353\]\[1\] mod.u_cpu.rf_ram.memory\[354\]\[1\]
+ mod.u_cpu.rf_ram.memory\[355\]\[1\] _01920_ _02666_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_78_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08495__A2 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07432_ _01488_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11626__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07363_ _01537_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09444__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09102_ _03383_ _03387_ _03397_ _03402_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07294_ _01492_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09033_ _03258_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10763__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12051__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09935_ _04065_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12503__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11594__S _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _04018_ mod.u_cpu.rf_ram.memory\[53\]\[1\] _04015_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14537__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10365__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07871__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _02369_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09797_ _03788_ _03966_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07930__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10003__S _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10117__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _02585_ _03053_ _03054_ _01751_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__12806__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14687__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ mod.u_cpu.rf_ram.memory\[210\]\[1\] mod.u_cpu.rf_ram.memory\[211\]\[1\] _01807_
+ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08030__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10710_ _04601_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11690_ _05268_ mod.u_cpu.rf_ram.memory\[251\]\[0\] _05269_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10641_ mod.u_cpu.rf_ram.memory\[41\]\[0\] _04396_ _04554_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13360_ _06455_ _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09986__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _04218_ _04507_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08207__I _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07997__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11769__S _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _05634_ _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12990__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13291_ _06384_ _06385_ _06387_ _06388_ _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_154_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15030_ _00884_ net3 mod.u_cpu.rf_ram.memory\[202\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12042__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12242_ _05367_ _05611_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15312__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12173_ _05575_ mod.u_cpu.rf_ram.memory\[76\]\[0\] _05598_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08410__A2 _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _04885_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13298__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11055_ _04836_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10356__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15462__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10006_ _04096_ mod.u_cpu.rf_ram.memory\[516\]\[0\] _04113_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14098__I1 mod.u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__A1 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14814_ _00668_ net3 mod.u_cpu.rf_ram.memory\[280\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14745_ _00599_ net3 mod.u_cpu.rf_ram.memory\[315\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11957_ _05455_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__B _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ _04735_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14676_ _00530_ net3 mod.u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11888_ _05406_ mod.u_cpu.rf_ram.memory\[227\]\[1\] _05402_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13627_ _06415_ _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11608__I0 mod.u_cpu.rf_ram.memory\[265\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ _04569_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13558_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] mod.u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _06594_ _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12281__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07532__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12509_ _05343_ _05831_ _05832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13489_ _06539_ _06552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15228_ _01081_ net3 mod.u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15159_ _01012_ net3 mod.u_cpu.rf_ram.memory\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08401__A2 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07981_ _02135_ mod.u_cpu.rf_ram.memory\[102\]\[0\] _02288_ _02139_ _02289_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13289__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09720_ _03907_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10347__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__B _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08004__I2 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__B1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _03847_ mod.u_cpu.rf_ram.memory\[563\]\[0\] _03852_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08602_ _01852_ _02901_ _02908_ _01887_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09582_ _03758_ _03797_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08533_ _02225_ _02838_ _02839_ _01683_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07640__B _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11472__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13361__C _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _02059_ mod.u_cpu.rf_ram.memory\[372\]\[1\] _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _01500_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10557__I _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09417__A1 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ mod.u_cpu.rf_ram.memory\[432\]\[1\] mod.u_cpu.rf_ram.memory\[433\]\[1\] mod.u_cpu.rf_ram.memory\[434\]\[1\]
+ mod.u_cpu.rf_ram.memory\[435\]\[1\] _02688_ _02475_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_195_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09968__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07346_ _01489_ _01629_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13868__I _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07523__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15335__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12972__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ _01572_ _01576_ _01583_ _01584_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07866__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ mod.u_cpu.cpu.state.o_cnt_r\[2\] mod.u_cpu.cpu.ctrl.i_iscomp _03321_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12024__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08079__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13921__B1 _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15485__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09918_ _04054_ mod.u_cpu.rf_ram.memory\[531\]\[1\] _04052_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10338__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08156__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09353__B1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _03771_ _03996_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12860_ _06060_ mod.u_cpu.rf_ram_if.rtrig1 _06061_ mod.u_cpu.rf_ram.regzero _01102_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11811_ _05342_ mod.u_cpu.rf_ram.memory\[49\]\[0\] _05352_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12791_ _05105_ _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14530_ _00384_ net3 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11742_ _05304_ mod.u_cpu.rf_ram.memory\[240\]\[1\] _05302_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11463__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14461_ _00315_ net3 mod.u_cpu.rf_ram.memory\[457\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _05250_ mod.u_cpu.rf_ram.memory\[250\]\[1\] _05256_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09408__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10018__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13412_ _03910_ _06011_ _06503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10624_ _04544_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14392_ _00246_ net3 mod.u_cpu.rf_ram.memory\[491\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__S0 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11499__S _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13343_ _06437_ _06418_ _06403_ _06439_ _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _03761_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07285__I3 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14702__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _06371_ _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10486_ _04450_ mod.u_cpu.rf_ram.memory\[445\]\[1\] _04448_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07709__C _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12715__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15013_ _00867_ net3 mod.u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12225_ _05404_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13727__B _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _05583_ mod.u_cpu.rf_ram.memory\[206\]\[1\] _05585_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14852__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12318__I1 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _04024_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10329__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12087_ _05539_ mod.u_cpu.rf_ram.memory\[65\]\[0\] _05540_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09195__I0 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11038_ _04796_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08537__I3 mod.u_cpu.rf_ram.memory\[291\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09895__A1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13691__A2 _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15208__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12989_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _06161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14728_ _00582_ net3 mod.u_cpu.rf_ram.memory\[323\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14232__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15358__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14659_ _00513_ net3 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_159_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08180_ _02483_ mod.u_cpu.rf_ram.memory\[558\]\[0\] _02486_ _02487_ _02488_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07131_ _01437_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08622__A2 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14382__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07686__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10568__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08511__S _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08481__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07964_ _01537_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08138__A1 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09186__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _03724_ _03892_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07895_ mod.u_cpu.rf_ram.memory\[217\]\[0\] _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09634_ _02510_ _03838_ _03839_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09565_ _03784_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08516_ mod.u_cpu.rf_ram.memory\[344\]\[1\] mod.u_cpu.rf_ram.memory\[345\]\[1\] mod.u_cpu.rf_ram.memory\[346\]\[1\]
+ mod.u_cpu.rf_ram.memory\[347\]\[1\] _02751_ _02748_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11296__I1 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09496_ _03718_ _03721_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08310__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10287__I _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08447_ _02230_ _02750_ _02753_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14725__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12245__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _02560_ _02683_ _02684_ _02594_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _01568_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08613__A2 _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10340_ _04345_ mod.u_cpu.rf_ram.memory\[468\]\[1\] _04349_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14875__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _04302_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12010_ _05490_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08129__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__I0 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13122__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08220__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13961_ mod.u_arbiter.i_wb_cpu_rdt\[3\] _06906_ _06928_ _03441_ _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09877__A1 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13673__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12912_ _06097_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11684__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13892_ _03872_ _06223_ _06882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10731__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14255__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12843_ _06051_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15631_ _01402_ net3 mod.u_cpu.rf_ram.memory\[244\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09629__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15500__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13425__A2 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15562_ _01333_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12484__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12774_ mod.u_cpu.rf_ram.memory\[133\]\[1\] _06005_ _06003_ _06006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14513_ _00367_ net3 mod.u_cpu.rf_ram.memory\[431\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11987__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10197__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11725_ _03857_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15493_ _01264_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14444_ _00298_ net3 mod.u_cpu.rf_ram.memory\[465\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11039__I1 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11656_ _05245_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12936__B2 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10607_ _04531_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14375_ _00229_ net3 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08604__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ _05143_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13326_ _06130_ _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10538_ _04481_ mod.u_cpu.rf_ram.memory\[436\]\[1\] _04483_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12539__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13257_ _06355_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10469_ _04043_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08368__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13361__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12208_ _03698_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13188_ _06291_ _06293_ _06281_ _06294_ _06295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10175__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12139_ _05520_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15030__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__I0 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09226__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07591__A2 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11675__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07680_ _01981_ _01984_ _01987_ _01972_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10722__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__A1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07974__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15180__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12587__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09350_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _03594_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14748__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09096__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08301_ _02590_ _02596_ _02102_ _02607_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09281_ _03517_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08232_ _02525_ _02531_ _02538_ _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_166_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12227__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14898__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08163_ _01688_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13211__I _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09643__I1 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10789__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _01421_ _01422_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _02348_ _02394_ _02401_ _02185_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10166__A1 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10570__I _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08996_ _03261_ mod.u_cpu.cpu.bufreg.i_sh_signed _03300_ _01422_ _03301_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__09159__I0 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14152__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14278__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08040__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _02170_ _02243_ _02254_ _02207_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12698__S _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13655__A2 _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15523__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08975__I mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11666__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07878_ _02170_ _02173_ _02184_ _02185_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08908__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _03800_ mod.u_cpu.rf_ram.memory\[567\]\[1\] _03824_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09548_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11969__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ mod.u_cpu.cpu.decode.op21 _01426_ _01440_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A2 _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ _05148_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12490_ _05819_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _05099_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09244__C1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13121__I _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14160_ _07070_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11372_ _05054_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08215__I _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08693__S1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13111_ _06230_ mod.u_cpu.rf_ram.memory\[100\]\[0\] _06242_ _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10323_ _04180_ _04327_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14091_ _02258_ _07025_ _07027_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15053__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13343__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13042_ _06186_ mod.u_cpu.rf_ram.memory\[107\]\[0\] _06197_ _06198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10254_ _03985_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09011__A2 _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08445__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10185_ _04241_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14993_ _00847_ net3 mod.u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13944_ _06913_ _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10704__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13875_ mod.u_cpu.cpu.immdec.imm24_20\[4\] _06868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15614_ _01385_ net3 mod.u_cpu.rf_ram.memory\[289\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11409__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12826_ _06032_ _06040_ _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15545_ _01316_ net3 mod.u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12757_ _05984_ mod.u_cpu.rf_ram.memory\[80\]\[1\] _05993_ _05995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11708_ _02269_ _05280_ _05281_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15476_ _00006_ net3 mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ _03734_ _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14427_ _00281_ net3 mod.u_cpu.rf_ram.memory\[474\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11639_ _05177_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08589__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12385__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14358_ _00212_ net3 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10396__A1 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13966__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13309_ _06405_ _06406_ _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14289_ _00143_ net3 mod.u_cpu.rf_ram.memory\[543\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07651__I3 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08436__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13885__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14420__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15546__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11486__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _02356_ mod.u_cpu.rf_ram.memory\[36\]\[1\] _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07801_ _01701_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08781_ _02104_ _03068_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ _01444_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11648__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14570__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07663_ _01697_ mod.u_cpu.rf_ram.memory\[302\]\[0\] _01969_ _01970_ _01971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10171__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13206__I _06312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09402_ _03637_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07594_ mod.u_cpu.rf_ram.memory\[352\]\[0\] mod.u_cpu.rf_ram.memory\[353\]\[0\] mod.u_cpu.rf_ram.memory\[354\]\[0\]
+ mod.u_cpu.rf_ram.memory\[355\]\[0\] _01841_ _01844_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09333_ _03578_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12073__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _03520_ _03521_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_21_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11671__I1 mod.u_cpu.rf_ram.memory\[250\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _02097_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09195_ mod.u_arbiter.i_wb_cpu_rdt\[23\] mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] _03469_
+ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15076__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08146_ _02453_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ _01924_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14913__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14125__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08979_ mod.u_cpu.cpu.state.init_done _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11990_ _05464_ mod.u_cpu.rf_ram.memory\[559\]\[1\] _05475_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08504__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ _04757_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13660_ _06671_ _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _04711_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14053__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12611_ _05891_ mod.u_cpu.rf_ram.memory\[153\]\[1\] _05897_ _05899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12064__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13591_ _06616_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11111__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09855__I1 mod.u_cpu.rf_ram.memory\[540\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13800__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15330_ _01106_ net3 mod.u_cpu.rf_ram.memory\[246\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12542_ _05827_ mod.u_cpu.rf_ram.memory\[164\]\[0\] _05852_ _05853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15419__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15261_ _00017_ net4 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10475__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07491__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12473_ _05808_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08115__S0 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14212_ _03968_ _05120_ _07103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11424_ _05088_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15192_ _01045_ net3 mod.u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09232__A2 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14443__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15569__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14143_ _07060_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11355_ _05028_ mod.u_cpu.rf_ram.memory\[306\]\[0\] _05042_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13316__A1 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10306_ _04163_ _04327_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08991__A1 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14074_ _07016_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11286_ _04995_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11178__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13025_ _05535_ _06080_ _06187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10237_ _04276_ mod.u_cpu.rf_ram.memory\[483\]\[0\] _04278_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14593__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09791__I0 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10168_ _03898_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _04179_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14976_ _00830_ net3 mod.u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13927_ _06017_ _06903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11350__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13858_ _06435_ _06370_ _06436_ _06852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12809_ mod.u_cpu.rf_ram.memory\[229\]\[1\] _06005_ _06027_ _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13789_ mod.u_arbiter.i_wb_cpu_rdt\[26\] _03449_ _03502_ _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07959__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15099__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15528_ _01299_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08283__C _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07482__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15459_ _01233_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08000_ _01716_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08982__A1 mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14936__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ _01463_ _03722_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_144_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11169__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13858__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08902_ _02507_ _03208_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09882_ _03805_ _04003_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08734__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09782__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08833_ _01592_ _03130_ _03139_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13137__S _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08764_ _02298_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07715_ mod.u_cpu.rf_ram.memory\[269\]\[0\] _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08695_ mod.u_cpu.rf_ram.memory\[197\]\[1\] _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14316__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07646_ _01918_ _01948_ _01953_ _01929_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13094__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07577_ _01874_ _01878_ _01883_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09316_ _03563_ _03565_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13794__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A2 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14466__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07473__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _03460_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08129_ _02157_ _02436_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11140_ _04895_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13849__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11071_ _04845_ _04848_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08725__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10022_ _04124_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11580__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14830_ _00684_ net3 mod.u_cpu.rf_ram.memory\[272\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08368__C _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11973_ _05465_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12285__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11088__A2 _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14761_ _00615_ net3 mod.u_cpu.rf_ram.memory\[307\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11332__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13712_ _06363_ _06712_ _06719_ _06135_ _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10924_ _04541_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14692_ _00546_ net3 mod.u_cpu.rf_ram.memory\[341\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15241__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__A2 _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13643_ _03390_ _06654_ _06137_ _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13085__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14809__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10855_ _04640_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12685__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12588__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13574_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] mod.u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _06604_ _06607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _04238_ _04648_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09453__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15391__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12525_ _05164_ _04302_ _05842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15313_ mod.u_scanchain_local.module_data_in\[69\] net4 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14959__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12456_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _05793_ _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15244_ _00019_ net4 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11399__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _05077_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15175_ _01028_ net3 mod.u_cpu.rf_ram.memory\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12387_ _05744_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14126_ _07049_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11338_ _04795_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14057_ mod.u_arbiter.i_wb_cpu_rdt\[27\] _06998_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _07005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11269_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08716__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13008_ _06107_ mod.u_cpu.rf_ram.memory\[86\]\[0\] _06175_ _06176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08811__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14339__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09234__I _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14959_ _00813_ net3 mod.u_cpu.rf_ram.memory\[549\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07500_ mod.u_cpu.rf_ram.memory\[447\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08480_ _02778_ _02779_ _02786_ _02007_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14489__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07431_ _01458_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__S0 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07689__I _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13776__A1 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07362_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12823__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__I1 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07293_ _01536_ _01593_ _01600_ _01587_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09032_ _03334_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11939__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15114__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04054_ mod.u_cpu.rf_ram.memory\[528\]\[1\] _04063_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08707__A1 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09755__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12503__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10514__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11562__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ mod.u_cpu.rf_ram.memory\[29\]\[1\] _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15264__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _03704_ _03938_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12267__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ _02156_ mod.u_cpu.rf_ram.memory\[108\]\[1\] _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10117__I1 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11314__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _02543_ _02981_ _02984_ _01632_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13822__C _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08916__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ _01643_ mod.u_cpu.rf_ram.memory\[308\]\[0\] _01936_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13067__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _04527_ _04389_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09435__A2 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10571_ _04436_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13519__A1 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12310_ _05691_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13290_ mod.u_arbiter.i_wb_cpu_rdt\[4\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _06122_ _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12241_ _05604_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12172_ _05325_ _05576_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _04883_ mod.u_cpu.rf_ram.memory\[343\]\[0\] _04884_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15607__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11054_ _04827_ mod.u_cpu.rf_ram.memory\[353\]\[0\] _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10005_ _03961_ _04087_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14813_ _00667_ net3 mod.u_cpu.rf_ram.memory\[281\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11305__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14631__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09123__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08557__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14744_ _00598_ net3 mod.u_cpu.rf_ram.memory\[315\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11956_ _05450_ mod.u_cpu.rf_ram.memory\[218\]\[1\] _05453_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _04728_ mod.u_cpu.rf_ram.memory\[376\]\[0\] _04734_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14675_ _00529_ net3 mod.u_cpu.rf_ram.memory\[350\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11887_ _05405_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14781__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _04686_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13626_ _06111_ _06112_ _06639_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13557_ _06597_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10769_ _04496_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__S1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12508_ _05725_ _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13488_ _06537_ _06551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15137__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14183__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12439_ _05778_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10663__I _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15227_ _01080_ net3 mod.u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10044__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15158_ _01011_ net3 mod.u_cpu.rf_ram.memory\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10744__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13974__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14109_ _07038_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15089_ _00943_ net3 mod.u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07980_ _02136_ _02287_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15287__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12497__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08289__B _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09362__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09650_ _03814_ _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09362__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08601_ _02323_ _02904_ _02907_ _01631_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09581_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12249__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13415__S _06503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08548__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ _02059_ mod.u_cpu.rf_ram.memory\[300\]\[1\] _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08463_ _01858_ _02769_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07676__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11472__A2 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13214__I _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07414_ _01633_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08394_ _02686_ _02690_ _02105_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _01632_ _01639_ _01652_ _01618_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07428__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__S1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07276_ _01528_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09015_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14504__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13921__A1 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13921__B2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10735__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07600__A1 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07882__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _04017_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10338__I1 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__C _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14654__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09848_ _04006_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _03936_ mod.u_cpu.rf_ram.memory\[550\]\[1\] _03952_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _04808_ _03866_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12790_ _06016_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09602__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08646__C _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11741_ _05249_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07667__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11463__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12660__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14460_ _00314_ net3 mod.u_cpu.rf_ram.memory\[457\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11672_ _05257_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08218__I _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10623_ _04537_ mod.u_cpu.rf_ram.memory\[423\]\[1\] _04540_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07419__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13411_ _06502_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12963__I _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14391_ _00245_ net3 mod.u_cpu.rf_ram.memory\[492\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13342_ _06438_ _06390_ _06439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07514__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08711__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10554_ _04495_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08092__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A1 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14165__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13273_ _06322_ _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _04429_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09049__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13912__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12224_ _02330_ _05632_ _05633_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15012_ _00866_ net3 mod.u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10726__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09592__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12155_ _05586_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13727__C _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09719__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11106_ _04872_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12086_ _04973_ _05388_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10329__I1 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11037_ _04824_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09647__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12988_ _06160_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14727_ _00581_ net3 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07658__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11939_ _03780_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14658_ _00512_ net3 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13609_ _03365_ _06625_ _06627_ _06628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14589_ _00443_ net3 mod.u_cpu.rf_ram.memory\[393\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14527__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07130_ mod.u_cpu.rf_ram_if.rtrig0 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07830__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09958__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14677__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07963_ _02244_ mod.u_cpu.rf_ram.memory\[252\]\[0\] _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07635__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08138__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09186__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _03807_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07894_ _01779_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09633_ _03775_ _03838_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07897__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11952__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09564_ _03740_ mod.u_cpu.rf_ram.memory\[572\]\[0\] _03783_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _02759_ _02818_ _02821_ _02764_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09495_ _03374_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15302__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A2 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _02730_ _02752_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13198__A2 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08377_ _02656_ mod.u_cpu.rf_ram.memory\[428\]\[1\] _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12245__I1 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07877__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07328_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__15452__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08074__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07259_ _01495_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09949__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10708__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11756__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08377__A2 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13960_ _03444_ _06917_ _06918_ _06931_ _06932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11133__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09877__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12911_ _06088_ mod.u_cpu.rf_ram.memory\[399\]\[0\] _06096_ _06097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12958__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13891_ _01426_ _06881_ _06800_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12881__A1 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10731__I1 mod.u_cpu.rf_ram.memory\[404\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11862__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15630_ _01401_ net3 mod.u_cpu.rf_ram.memory\[279\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _06038_ mod.u_cpu.rf_ram.memory\[123\]\[1\] _06049_ _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09629__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15561_ _01332_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12773_ _03734_ _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13830__B1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13830__C2 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14512_ _00366_ net3 mod.u_cpu.rf_ram.memory\[431\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11724_ _05292_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15492_ _01263_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14443_ _00297_ net3 mod.u_cpu.rf_ram.memory\[466\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ _05243_ mod.u_cpu.rf_ram.memory\[258\]\[0\] _05244_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10606_ _03733_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14374_ _00228_ net3 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11586_ _05198_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11995__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10537_ _04484_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13325_ _06421_ _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _03991_ _04437_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13256_ _06354_ mod.u_cpu.rf_ram.memory\[95\]\[1\] _06352_ _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11747__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08368__A2 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12207_ _05621_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13187_ _06284_ _06294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10399_ mod.u_cpu.rf_ram.memory\[45\]\[1\] _04383_ _04390_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10175__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _05574_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12069_ _05521_ mod.u_cpu.rf_ram.memory\[63\]\[0\] _05528_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07879__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15325__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11675__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08540__A2 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07974__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08679__I0 mod.u_cpu.rf_ram.memory\[210\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08300_ _02083_ _02598_ _02605_ _02606_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10486__I0 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09280_ _03495_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15475__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08231_ _02120_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07697__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ _02449_ _02452_ _02468_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08056__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__B1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ mod.u_cpu.cpu.branch_op _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08093_ _02352_ _02397_ _02400_ _02361_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13888__B1 _06877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10851__I _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10166__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08995_ _03280_ _03299_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07946_ _02174_ _02248_ _02253_ _01766_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07877_ _01551_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09616_ _02513_ _03824_ _03825_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08196__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10298__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09547_ _03768_ _03749_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10477__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09478_ _01660_ _03703_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08429_ _02534_ mod.u_cpu.rf_ram.memory\[404\]\[1\] _02735_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14842__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13415__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11440_ _05087_ mod.u_cpu.rf_ram.memory\[292\]\[1\] _05097_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08047__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09244__B1 _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09244__C2 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11371_ _05050_ mod.u_cpu.rf_ram.memory\[304\]\[1\] _05052_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08940__B _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10322_ _04338_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13110_ _03960_ _06223_ _06242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14090_ _07026_ _07025_ _07027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14992__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11729__I0 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13041_ _05606_ _06092_ _06197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10253_ _04289_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13343__A2 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11354__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__I _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10184_ _04215_ mod.u_cpu.rf_ram.memory\[491\]\[1\] _04239_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14222__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15348__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__I1 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08770__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14992_ _00846_ net3 mod.u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12154__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13943_ _06912_ _06917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12854__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14372__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13874_ _06412_ _06834_ _06867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15498__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15613_ _01384_ net3 mod.u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11409__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12825_ _03770_ _06030_ _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09997__I _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15544_ _01315_ net3 mod.u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12756_ _05994_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10093__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11707_ _05265_ _05280_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15475_ _00005_ net3 mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12687_ _02370_ _05947_ _05949_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14426_ _00280_ net3 mod.u_cpu.rf_ram.memory\[474\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08038__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _05233_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07310__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08589__A2 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14357_ _00211_ net3 mod.u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11569_ _04066_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10396__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11593__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13308_ _06374_ _06362_ _06406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14288_ _00142_ net3 mod.u_cpu.rf_ram.memory\[543\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10671__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13239_ _06343_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08141__I _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12799__S _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ mod.u_cpu.rf_ram.memory\[168\]\[0\] mod.u_cpu.rf_ram.memory\[169\]\[0\] mod.u_cpu.rf_ram.memory\[170\]\[0\]
+ mod.u_cpu.rf_ram.memory\[171\]\[0\] _02106_ _02107_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08780_ _01446_ _03077_ _03086_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13098__A1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14715__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07731_ _01485_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12845__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13893__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09710__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11208__S _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08513__A2 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07662_ _01701_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10320__A2 _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09401_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _03627_
+ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14865__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07593_ _01852_ _01892_ _01900_ _01677_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_92_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11007__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _03574_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03560_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12073__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09263_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _03498_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_08214_ _02039_ _02493_ _02521_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09194_ _03451_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11959__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07220__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _01782_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ mod.u_cpu.rf_ram.memory\[4\]\[0\] mod.u_cpu.rf_ram.memory\[5\]\[0\] mod.u_cpu.rf_ram.memory\[6\]\[0\]
+ mod.u_cpu.rf_ram.memory\[7\]\[0\] _02366_ _02383_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14245__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10581__I _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14125__I1 mod.u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14395__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13089__A1 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08978_ _01430_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] mod.u_cpu.cpu.state.init_done
+ _03282_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07890__I _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15640__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ mod.u_cpu.rf_ram.memory\[231\]\[0\] _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08504__A2 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ _04756_ mod.u_cpu.rf_ram.memory\[371\]\[1\] _04754_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08060__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10871_ _04695_ mod.u_cpu.rf_ram.memory\[382\]\[0\] _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12610_ _05898_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13261__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13590_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] mod.u_arbiter.i_wb_cpu_dbus_adr\[28\]
+ _06614_ _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08654__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12541_ _05367_ _05831_ _05852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15020__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15260_ _00016_ net4 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08226__I _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12472_ _05807_ mod.u_cpu.rf_ram.memory\[419\]\[1\] _05804_ _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09768__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08115__S1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14211_ _07102_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11423_ _05087_ mod.u_cpu.rf_ram.memory\[295\]\[1\] _05085_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15191_ _01044_ net3 mod.u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14142_ _07055_ mod.u_cpu.rf_ram.memory\[289\]\[1\] _07058_ _07060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11354_ _04758_ _05038_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08440__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15170__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11587__I _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10305_ _04302_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13316__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08991__A2 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14073_ _06578_ mod.u_cpu.rf_ram.memory\[114\]\[0\] _07015_ _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11285_ _04988_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12375__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11178__I1 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14738__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10236_ _04277_ _04263_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13024_ _06072_ _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09940__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09791__I1 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _03896_ _04228_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08594__I2 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ _04178_ mod.u_cpu.rf_ram.memory\[503\]\[1\] _04174_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14975_ _00829_ net3 mod.u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14888__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13926_ _02304_ _06901_ _06902_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _06487_ _06850_ _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12808_ _02234_ _06027_ _06028_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13252__A1 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13788_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15527_ _01298_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12739_ _02215_ _05982_ _05983_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13004__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15458_ _01232_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14268__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14409_ _00263_ net3 mod.u_cpu.rf_ram.memory\[483\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15513__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15389_ _01164_ net3 mod.u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10369__A2 _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07975__I _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13307__A2 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09950_ _04076_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08982__A2 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08901_ mod.u_cpu.rf_ram.memory\[517\]\[1\] _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09881_ _04029_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09931__A1 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08832_ _02150_ _03131_ _03138_ _02363_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08739__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08763_ mod.u_cpu.rf_ram.memory\[125\]\[1\] _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12121__I _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07714_ _01704_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08498__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08694_ _01560_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07215__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13618__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07645_ _01938_ mod.u_cpu.rf_ram.memory\[294\]\[0\] _01951_ _01952_ _01953_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15043__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12046__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07576_ _01630_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09315_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13794__A2 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14048__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09246_ _03493_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07473__A2 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08670__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15193__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ _03458_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] _03459_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12791__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__I0 mod.u_cpu.rf_ram.memory\[425\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08128_ mod.u_cpu.rf_ram.memory\[45\]\[0\] _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08422__A1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _01524_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12357__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11070_ _04847_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10021_ _04115_ mod.u_cpu.rf_ram.memory\[514\]\[1\] _04122_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13127__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14760_ _00614_ net3 mod.u_cpu.rf_ram.memory\[307\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08489__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11972_ _05464_ mod.u_cpu.rf_ram.memory\[217\]\[1\] _05462_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12285__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07125__I mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11332__I1 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13711_ _06716_ _06718_ _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10923_ _04184_ _04713_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14691_ _00545_ net3 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07161__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07161__B2 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13642_ _03274_ _06653_ _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10854_ _04697_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10048__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14410__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13785__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15536__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13573_ _06606_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10785_ _04651_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15312_ _00073_ net4 mod.u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12524_ _05841_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08661__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15243_ _00008_ net4 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12455_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _03430_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14560__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11399__I1 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _05069_ mod.u_cpu.rf_ram.memory\[298\]\[1\] _05075_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08413__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15174_ _01027_ net3 mod.u_cpu.rf_ram.memory\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12386_ _05731_ mod.u_cpu.rf_ram.memory\[177\]\[0\] _05743_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14125_ _07041_ mod.u_cpu.rf_ram.memory\[116\]\[1\] _07047_ _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11337_ _05030_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12348__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14056_ _06970_ _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09213__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11268_ _04194_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13238__S _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13007_ _03828_ _06080_ _06175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08716__A2 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _04176_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12142__S _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11199_ _04918_ mod.u_cpu.rf_ram.memory\[330\]\[0\] _04934_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09515__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11720__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15066__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14958_ _00812_ net3 mod.u_cpu.rf_ram.memory\[549\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13909_ _06311_ _06861_ _06443_ _06647_ _06890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14889_ _00743_ net3 mod.u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08575__B _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ _01474_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13076__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07361_ _01491_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12823__I1 mod.u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09100_ _03385_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_176_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07292_ _01505_ _01596_ _01599_ _01584_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08652__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14903__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09031_ _01435_ mod.u_cpu.cpu.decode.co_ebreak _01452_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08955__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12339__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11020__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09933_ _04064_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09204__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__S _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08707__A2 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09864_ _03762_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15409__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08469__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ mod.u_cpu.rf_ram.memory\[24\]\[1\] mod.u_cpu.rf_ram.memory\[25\]\[1\] mod.u_cpu.rf_ram.memory\[26\]\[1\]
+ mod.u_cpu.rf_ram.memory\[27\]\[1\] _02366_ _02367_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09795_ _03965_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08746_ mod.u_cpu.rf_ram.memory\[109\]\[1\] _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12267__A2 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14433__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ _02462_ mod.u_cpu.rf_ram.memory\[214\]\[1\] _02983_ _02597_ _02984_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15559__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10300__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07628_ _01934_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08891__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11078__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13767__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07559_ _01503_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__A3 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14583__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10570_ _04452_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08643__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08705__S _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _03410_ mod.u_scanchain_local.module_data_in\[38\] _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12227__S _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12578__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12240_ _05644_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12026__I _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12171_ _05597_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11122_ _03879_ _04869_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _04285_ _04822_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15089__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08254__S0 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10004_ _04112_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__C _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14812_ _00666_ net3 mod.u_cpu.rf_ram.memory\[281\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11305__I1 mod.u_cpu.rf_ram.memory\[314\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09123__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14743_ _00597_ net3 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08557__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11955_ _05454_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07134__A1 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ _04732_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08882__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14674_ _00528_ net3 mod.u_cpu.rf_ram.memory\[350\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11886_ _05404_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14926__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13625_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _06111_ _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _04682_ mod.u_cpu.rf_ram.memory\[387\]\[1\] _04684_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13556_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] mod.u_arbiter.i_wb_cpu_dbus_adr\[13\]
+ _06594_ _06597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10768_ _04639_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12507_ _05830_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13487_ _06550_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _04593_ mod.u_cpu.rf_ram.memory\[410\]\[1\] _04591_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15226_ _01079_ net3 mod.u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12438_ _05753_ mod.u_cpu.rf_ram.memory\[172\]\[0\] _05777_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11241__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15157_ _01010_ net3 mod.u_cpu.rf_ram.memory\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12369_ _05732_ _04137_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14306__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14108_ _07028_ mod.u_cpu.rf_ram.memory\[117\]\[1\] _07036_ _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11792__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15088_ _00942_ net3 mod.u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11775__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14039_ _06990_ _06991_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12497__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12741__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14456__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08600_ _02136_ mod.u_cpu.rf_ram.memory\[262\]\[1\] _02906_ _01504_ _02907_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12249__A2 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ mod.u_cpu.rf_ram.memory\[301\]\[1\] _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08462_ mod.u_cpu.rf_ram.memory\[373\]\[1\] _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07676__A2 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10680__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _01696_ _01699_ _01718_ _01720_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13749__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08393_ _02083_ _02691_ _02699_ _02606_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07344_ _01572_ _01642_ _01650_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07275_ _01577_ mod.u_cpu.rf_ram.memory\[470\]\[0\] _01580_ _01582_ _01583_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12047__S _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09014_ _03297_ _03298_ _03255_ _03318_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08324__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12185__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09976__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13921__A2 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11932__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15231__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07600__A2 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09916_ _04053_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08236__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13685__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _03999_ mod.u_cpu.rf_ram.memory\[542\]\[1\] _04004_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15381__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08994__I mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ _03953_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14949__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08927__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08729_ _02632_ mod.u_cpu.rf_ram.memory\[246\]\[1\] _03035_ _01702_ _03036_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _05303_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07667__A2 _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07403__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11671_ _05243_ mod.u_cpu.rf_ram.memory\[250\]\[0\] _05256_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13410_ _06354_ mod.u_cpu.rf_ram.memory\[91\]\[1\] _06500_ _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12799__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10622_ _01760_ _04540_ _04543_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14390_ _00244_ net3 mod.u_cpu.rf_ram.memory\[492\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07419__A2 mod.u_cpu.rf_ram.memory\[404\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09664__I0 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13341_ _06374_ _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10553_ _04486_ mod.u_cpu.rf_ram.memory\[433\]\[0\] _04494_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08711__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__A2 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14329__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10974__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13272_ _06369_ _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08234__I _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _01803_ _04448_ _04449_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15011_ _00865_ net3 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12223_ _05581_ _05632_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09041__B2 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13296__B _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12154_ _05575_ mod.u_cpu.rf_ram.memory\[206\]\[0\] _05585_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14479__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _04862_ mod.u_cpu.rf_ram.memory\[346\]\[1\] _04870_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13676__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12085_ _05520_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13676__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11036_ _04803_ mod.u_cpu.rf_ram.memory\[356\]\[0\] _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13428__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13428__B2 _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10939__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12987_ _06158_ mod.u_cpu.cpu.genblk3.csr.mcause31 _06159_ _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13315__I _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14726_ _00580_ net3 mod.u_cpu.rf_ram.memory\[324\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11938_ _05412_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07658__A2 mod.u_cpu.rf_ram.memory\[300\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15104__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14657_ _00511_ net3 mod.u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11869_ _05385_ mod.u_cpu.rf_ram.memory\[72\]\[0\] _05392_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13608_ _03381_ _06626_ _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08607__A1 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13600__A1 _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14588_ _00442_ net3 mod.u_cpu.rf_ram.memory\[393\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13539_ _06587_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15254__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12167__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15209_ _01062_ net3 mod.u_cpu.rf_ram.memory\[219\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09958__I1 mod.u_cpu.rf_ram.memory\[524\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13903__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09032__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _02245_ _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09701_ _03891_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07346__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07893_ _02198_ _02199_ _02200_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09632_ _03834_ _03837_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09563_ _03758_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08514_ _02526_ _02819_ _02820_ _01501_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08846__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09494_ _01448_ _01454_ _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07223__I mod.u_cpu.raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08445_ mod.u_cpu.rf_ram.memory\[396\]\[1\] mod.u_cpu.rf_ram.memory\[397\]\[1\] mod.u_cpu.rf_ram.memory\[398\]\[1\]
+ mod.u_cpu.rf_ram.memory\[399\]\[1\] _02751_ _02748_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13161__S _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08376_ mod.u_cpu.rf_ram.memory\[429\]\[1\] _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14056__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07327_ _01634_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09271__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ _01536_ _01555_ _01565_ _01552_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_136_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14621__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09949__I1 mod.u_cpu.rf_ram.memory\[526\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09023__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07189_ mod.u_cpu.raddr\[1\] _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09574__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10025__S _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14771__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12910_ _04913_ _04570_ _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13890_ _06704_ _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12881__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__I _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15127__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ _06050_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07561__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14083__A1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13130__I0 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15560_ _01331_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08229__I _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12772_ _06004_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09885__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14511_ _00365_ net3 mod.u_cpu.rf_ram.memory\[432\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _05287_ mod.u_cpu.rf_ram.memory\[243\]\[1\] _05290_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15491_ _01262_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15277__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14442_ _00296_ net3 mod.u_cpu.rf_ram.memory\[466\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11654_ _04831_ _05214_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12397__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08392__C _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10605_ _04530_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14373_ _00227_ net3 mod.u_cpu.rf_ram.memory\[501\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11585_ _05194_ mod.u_cpu.rf_ram.memory\[26\]\[1\] _05196_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11995__I1 mod.u_cpu.rf_ram.memory\[569\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13324_ _06064_ _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10536_ _04469_ mod.u_cpu.rf_ram.memory\[436\]\[0\] _04483_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09014__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13255_ _06236_ _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10467_ _04436_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12206_ _05609_ mod.u_cpu.rf_ram.memory\[200\]\[1\] _05619_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13186_ _06292_ _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10398_ _02436_ _04390_ _04391_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12137_ _05566_ mod.u_cpu.rf_ram.memory\[74\]\[1\] _05572_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12068_ _04294_ _04845_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11019_ _04811_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10635__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14709_ _00563_ net3 mod.u_cpu.rf_ram.memory\[333\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ _02533_ mod.u_cpu.rf_ram.memory\[518\]\[0\] _02536_ _02537_ _02538_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14644__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _02143_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09253__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08056__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07112_ mod.u_cpu.cpu.decode.opcode\[2\] _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08092_ _02356_ mod.u_cpu.rf_ram.memory\[30\]\[0\] _02399_ _02359_ _02400_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13888__B2 _06879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14794__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10410__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ mod.u_cpu.cpu.bne_or_bge _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07945_ _02249_ mod.u_cpu.rf_ram.memory\[238\]\[0\] _02251_ _02252_ _02253_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07319__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12163__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07876_ _02174_ _02178_ _02183_ _02166_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09433__I mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09615_ _03775_ _03824_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _03701_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10477__I1 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09477_ _01439_ _01494_ mod.u_cpu.raddr\[1\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_169_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08428_ _02526_ _02734_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13415__I1 mod.u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12379__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08359_ _01762_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09244__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08047__A2 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11370_ _05053_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _04330_ mod.u_cpu.rf_ram.memory\[471\]\[1\] _04336_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13040_ _06196_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09547__A2 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ _04288_ mod.u_cpu.rf_ram.memory\[481\]\[1\] _04286_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13343__A3 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07558__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10183_ _04240_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14991_ _00845_ net3 mod.u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12303__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13942_ _06123_ _06906_ _06911_ _03431_ _06916_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14517__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10489__I _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13873_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06865_ _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_46_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07730__A1 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13103__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15612_ _01383_ net3 mod.u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12824_ _06039_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15543_ _01314_ net3 mod.u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14667__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12755_ _05992_ mod.u_cpu.rf_ram.memory\[80\]\[0\] _05993_ _05994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10093__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _04994_ _05279_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15474_ _01248_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12686_ _05948_ _05947_ _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14425_ _00279_ net3 mod.u_cpu.rf_ram.memory\[475\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11417__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11637_ _05222_ mod.u_cpu.rf_ram.memory\[260\]\[0\] _05232_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11042__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14356_ _00210_ net3 mod.u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11568_ _05186_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13307_ _06368_ _06404_ _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10519_ _04251_ _03911_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14287_ _00141_ net3 mod.u_cpu.rf_ram.memory\[544\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11499_ _05114_ mod.u_cpu.rf_ram.memory\[283\]\[0\] _05140_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13238_ _06276_ mod.u_cpu.rf_ram.memory\[94\]\[1\] _06341_ _06343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13590__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13169_ _06277_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13098__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07730_ _01481_ _01817_ _02037_ _01469_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12845__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15442__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08297__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07661_ _01967_ _01968_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07721__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ _03635_ _03632_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07592_ _01874_ _01896_ _01899_ _01884_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09331_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15592__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09262_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08213_ _02506_ _02519_ _02520_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ _03468_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11959__I1 mod.u_cpu.rf_ram.memory\[529\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08144_ mod.u_cpu.rf_ram.memory\[544\]\[0\] mod.u_cpu.rf_ram.memory\[545\]\[0\] mod.u_cpu.rf_ram.memory\[546\]\[0\]
+ mod.u_cpu.rf_ram.memory\[547\]\[0\] _02450_ _02451_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12081__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08760__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10862__I _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _01524_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12908__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12533__A1 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ mod.u_cpu.cpu.state.stage_two_req _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07928_ _02175_ mod.u_cpu.rf_ram.memory\[228\]\[0\] _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14038__A1 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ _02155_ _02160_ _02165_ _02166_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08060__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ _04299_ _04709_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08935__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13797__B1 _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _03715_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11134__S _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12540_ _05851_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11272__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07411__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12471_ _05806_ _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14210_ mod.u_cpu.rf_ram.memory\[269\]\[1\] _06221_ _07100_ _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11422_ _05031_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15190_ _01043_ net3 mod.u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08670__C _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15315__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14141_ _07059_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11353_ _05041_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10304_ _04248_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08242__I _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14072_ _03858_ _07014_ _07015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11284_ _03769_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13023_ _06185_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14180__S _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10235_ _03968_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15465__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09940__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10166_ _04225_ _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14974_ _00828_ net3 mod.u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13925_ _06249_ _06901_ _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10012__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13856_ _06397_ _06292_ _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12807_ _05948_ _06027_ _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13787_ _06774_ _06787_ _06788_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10999_ _04797_ mod.u_cpu.rf_ram.memory\[362\]\[1\] _04793_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15526_ _01297_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12738_ _05843_ _05982_ _05983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10310__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12460__B1 _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15457_ _01231_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12669_ _05709_ _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14408_ _00262_ net3 mod.u_cpu.rf_ram.memory\[483\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11015__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15388_ _01163_ net3 mod.u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__I2 mod.u_cpu.rf_ram.memory\[314\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14339_ _00193_ net3 mod.u_cpu.rf_ram.memory\[518\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14154__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12515__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ mod.u_cpu.rf_ram.memory\[512\]\[1\] mod.u_cpu.rf_ram.memory\[513\]\[1\] mod.u_cpu.rf_ram.memory\[514\]\[1\]
+ mod.u_cpu.rf_ram.memory\[515\]\[1\] _02494_ _02495_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09880_ _04018_ mod.u_cpu.rf_ram.memory\[537\]\[1\] _04027_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10377__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08814__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08195__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08831_ _02405_ _03134_ _03137_ _02415_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09931__A2 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14832__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ mod.u_cpu.rf_ram.memory\[120\]\[1\] mod.u_cpu.rf_ram.memory\[121\]\[1\] mod.u_cpu.rf_ram.memory\[122\]\[1\]
+ mod.u_cpu.rf_ram.memory\[123\]\[1\] _02294_ _02295_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ mod.u_cpu.rf_ram.memory\[264\]\[0\] mod.u_cpu.rf_ram.memory\[265\]\[0\] mod.u_cpu.rf_ram.memory\[266\]\[0\]
+ mod.u_cpu.rf_ram.memory\[267\]\[0\] _02020_ _01995_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09695__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08498__A2 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ mod.u_cpu.rf_ram.memory\[192\]\[1\] mod.u_cpu.rf_ram.memory\[193\]\[1\] mod.u_cpu.rf_ram.memory\[194\]\[1\]
+ mod.u_cpu.rf_ram.memory\[195\]\[1\] _01578_ _01714_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_39_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _01782_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14982__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ _01879_ mod.u_cpu.rf_ram.memory\[374\]\[0\] _01881_ _01882_ _01883_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09314_ _03486_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07231__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15338__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09245_ _03505_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12054__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09176_ _03451_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11688__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12754__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ mod.u_cpu.rf_ram.memory\[40\]\[0\] mod.u_cpu.rf_ram.memory\[41\]\[0\] mod.u_cpu.rf_ram.memory\[42\]\[0\]
+ mod.u_cpu.rf_ram.memory\[43\]\[0\] _02151_ _02383_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10604__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14362__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15488__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ _02058_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12357__I1 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10020_ _04123_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07834__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13852__B _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11971_ _05405_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09686__A1 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08489__A2 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13710_ _06694_ _06363_ _06717_ _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10922_ _04744_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14690_ _00544_ net3 mod.u_cpu.rf_ram.memory\[342\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__I _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08665__C _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13641_ _03297_ mod.u_cpu.cpu.decode.opcode\[1\] _06652_ _06653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _04695_ mod.u_cpu.rf_ram.memory\[384\]\[0\] _04696_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13234__A2 _06340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__I _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13572_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] mod.u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _06604_ _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12293__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10784_ _04641_ mod.u_cpu.rf_ram.memory\[396\]\[1\] _04649_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08110__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15311_ _00072_ net4 mod.u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12523_ _05837_ mod.u_cpu.rf_ram.memory\[166\]\[1\] _05839_ _05841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14705__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15242_ _01095_ net3 mod.u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12454_ _03281_ _05791_ _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11405_ _05076_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13942__B1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15173_ _01026_ net3 mod.u_cpu.rf_ram.memory\[148\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12385_ _05742_ _05726_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14124_ _07048_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11336_ _05028_ mod.u_cpu.rf_ram.memory\[30\]\[0\] _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14855__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14055_ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] _07000_ _07003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10359__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11267_ _04981_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13170__A1 _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13006_ _06174_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10218_ _04265_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11198_ _04792_ _04926_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10149_ _01648_ _04213_ _04214_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13762__B _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14957_ _00811_ net3 mod.u_cpu.rf_ram.memory\[217\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__B _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13908_ _03681_ _06641_ _06887_ _06889_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08348__S _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14888_ _00742_ net3 mod.u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14235__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13839_ _06138_ _06834_ _06835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09429__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13053__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08147__I _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _01662_ _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08101__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15509_ _01280_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07291_ _01545_ mod.u_cpu.rf_ram.memory\[502\]\[0\] _01598_ _01582_ _01599_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14385__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07986__I _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09030_ _03290_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15630__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04051_ mod.u_cpu.rf_ram.memory\[528\]\[0\] _04063_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09863_ _04016_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09904__A2 _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07915__A1 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _03117_ _03118_ _03119_ _03120_ _02391_ _01720_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09794_ _03964_ mod.u_cpu.rf_ram.memory\[548\]\[1\] _03962_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15010__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08745_ mod.u_cpu.rf_ram.memory\[110\]\[1\] mod.u_cpu.rf_ram.memory\[111\]\[1\] _01508_
+ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11971__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ _01705_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08340__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ mod.u_cpu.rf_ram.memory\[309\]\[0\] _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15160__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14728__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07558_ _01864_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08057__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__S0 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12975__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09435__A4 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ _01779_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07896__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11412__S _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12027__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _03485_ _03490_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14878__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09159_ mod.u_arbiter.i_wb_cpu_rdt\[9\] mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _03442_
+ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12170_ mod.u_cpu.rf_ram.memory\[205\]\[1\] _05468_ _05595_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13527__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11121_ _04882_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11002__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ _04834_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08254__S1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ mod.u_cpu.rf_ram.memory\[517\]\[1\] _04111_ _04109_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07136__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14258__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14811_ _00665_ net3 mod.u_cpu.rf_ram.memory\[282\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11881__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15503__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11954_ _05442_ mod.u_cpu.rf_ram.memory\[218\]\[0\] _05453_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14742_ _00596_ net3 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10905_ _04708_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14673_ _00527_ net3 mod.u_cpu.rf_ram.memory\[351\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11885_ _05105_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13624_ _06638_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10836_ _04685_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13555_ _06596_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10767_ _04637_ mod.u_cpu.rf_ram.memory\[398\]\[0\] _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12018__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12506_ _05822_ mod.u_cpu.rf_ram.memory\[16\]\[1\] _05828_ _05830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13486_ _03610_ _06545_ _06546_ _03616_ _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10698_ _04578_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15225_ _01078_ net3 mod.u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12437_ _05325_ _05767_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11121__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08398__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15156_ _01009_ net3 mod.u_cpu.rf_ram.memory\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11241__I1 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12368_ _03849_ _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14107_ _02326_ _07036_ _07037_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11319_ _05014_ mod.u_cpu.rf_ram.memory\[312\]\[1\] _05016_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15087_ _00941_ net3 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15033__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12299_ _05684_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__B1 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14038_ mod.u_arbiter.i_wb_cpu_rdt\[22\] _06987_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _06991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15183__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08530_ mod.u_cpu.rf_ram.memory\[302\]\[1\] mod.u_cpu.rf_ram.memory\[303\]\[1\] _02272_
+ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11457__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10504__I0 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08322__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__S0 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08461_ mod.u_cpu.rf_ram.memory\[368\]\[1\] mod.u_cpu.rf_ram.memory\[369\]\[1\] mod.u_cpu.rf_ram.memory\[370\]\[1\]
+ mod.u_cpu.rf_ram.memory\[371\]\[1\] _01837_ _01838_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08873__A2 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07412_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12257__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08392_ _02188_ _02695_ _02698_ _02196_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07343_ _01528_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12009__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09013_ _01431_ _03305_ _03311_ _03317_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12709__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12185__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13159__S _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11932__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09915_ _04051_ mod.u_cpu.rf_ram.memory\[531\]\[0\] _04052_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08236__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09889__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14400__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13685__A2 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15526__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _04005_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09777_ _03916_ mod.u_cpu.rf_ram.memory\[550\]\[0\] _03952_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _02084_ _03034_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14550__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11299__I1 mod.u_cpu.rf_ram.memory\[315\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__I _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07116__A2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07747__S0 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11999__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ mod.u_cpu.rf_ram.memory\[221\]\[1\] _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A1 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08864__A2 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11670_ _04868_ _05255_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12948__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ _04542_ _04540_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13340_ _06436_ _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10552_ _04360_ _04487_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13271_ _06367_ _06368_ _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10483_ _04439_ _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15056__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15010_ _00864_ net3 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13373__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12222_ _05019_ _05631_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13912__A3 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12153_ _05312_ _05568_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10780__I _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10982__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11104_ _04871_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09329__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12084_ _05538_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13676__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11035_ _04821_ _04822_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14201__B _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12487__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12986_ _06063_ _03335_ _03375_ _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14725_ _00579_ net3 mod.u_cpu.rf_ram.memory\[325\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11937_ _05441_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11116__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14656_ _00510_ net3 mod.u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11868_ _05343_ _05388_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08853__C _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13607_ _03309_ _06625_ _06626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10819_ _04674_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11799_ _05342_ mod.u_cpu.rf_ram.memory\[232\]\[0\] _05344_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14587_ _00441_ net3 mod.u_cpu.rf_ram.memory\[394\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13600__A2 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11611__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13538_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] mod.u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _06584_ _06587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07291__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13469_ _06539_ _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10891__S _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13364__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12167__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15208_ _01061_ net3 mod.u_cpu.rf_ram.memory\[219\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09032__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14423__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15549__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15139_ _00992_ net3 mod.u_cpu.rf_ram.memory\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ mod.u_cpu.rf_ram.memory\[253\]\[0\] _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13667__A2 _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09700_ _03890_ mod.u_cpu.rf_ram.memory\[558\]\[1\] _03887_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07892_ _01517_ mod.u_cpu.rf_ram.memory\[218\]\[0\] _01714_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14573__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13934__C _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08543__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09631_ _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07932__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _03781_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07504__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08513_ _01605_ mod.u_cpu.rf_ram.memory\[348\]\[1\] _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09493_ _01448_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08846__A2 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _01919_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08375_ mod.u_cpu.rf_ram.memory\[430\]\[1\] mod.u_cpu.rf_ram.memory\[431\]\[1\] _02585_
+ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15079__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07326_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ _01505_ _01559_ _01564_ _01529_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10169__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07188_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10964__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14916__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12705__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09829_ _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12840_ _06035_ mod.u_cpu.rf_ram.memory\[123\]\[0\] _06049_ _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14083__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07414__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13130__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12771_ mod.u_cpu.rf_ram.memory\[133\]\[0\] _05971_ _06003_ _06004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14510_ _00364_ net3 mod.u_cpu.rf_ram.memory\[432\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11722_ _05291_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15490_ _01261_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _00295_ net3 mod.u_cpu.rf_ram.memory\[467\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11653_ _05221_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10604_ mod.u_cpu.rf_ram.memory\[425\]\[0\] _04396_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14372_ _00226_ net3 mod.u_cpu.rf_ram.memory\[501\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11584_ _05197_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14446__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13323_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _06358_ _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _04189_ _04464_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13254_ _06353_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _04435_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09014__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13897__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12205_ _05620_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13185_ mod.u_arbiter.i_wb_cpu_rdt\[6\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _06126_ _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10397_ _04230_ _04390_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14596__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09076__I _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08773__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12136_ _05573_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12067_ _05527_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13754__C _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _04797_ mod.u_cpu.rf_ram.memory\[35\]\[1\] _04809_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11380__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13326__I _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09025__B _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07324__I _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13770__B _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12969_ _03344_ _06144_ _06145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08384__S0 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14708_ _00562_ net3 mod.u_cpu.rf_ram.memory\[333\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15221__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08583__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14639_ _00493_ net3 mod.u_cpu.rf_ram.memory\[368\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08160_ _02455_ _02460_ _02466_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12632__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07111_ mod.u_cpu.cpu.decode.co_mem_word mod.u_cpu.cpu.bne_or_bge mod.u_cpu.cpu.csr_d_sel
+ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15371__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ _01823_ _02398_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14939__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11199__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13888__A2 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ _03253_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _01827_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13664__C _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09564__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08758__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ _02179_ mod.u_cpu.rf_ram.memory\[206\]\[0\] _02182_ _02164_ _02183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10323__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11371__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14319__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ _03767_ _03823_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12140__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14065__A2 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _03766_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13812__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09476_ _03701_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09492__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14469__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08427_ mod.u_cpu.rf_ram.memory\[405\]\[1\] _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10595__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08127__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12379__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08358_ _01991_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _01572_ _01611_ _01616_ _01584_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08289_ _02592_ _02595_ _02077_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13328__A1 _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _01579_ _04336_ _04337_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10251_ _04266_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12315__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10937__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14128__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10182_ _04217_ mod.u_cpu.rf_ram.memory\[491\]\[0\] _04239_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14990_ _00844_ net3 mod.u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08507__A1 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12303__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13500__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13941_ _03431_ _06912_ _06915_ _06916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13872_ _03503_ mod.u_arbiter.i_wb_cpu_rdt\[23\] _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10865__A2 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15244__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15611_ _01382_ net3 mod.u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13103__I1 mod.u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12823_ _06038_ mod.u_cpu.rf_ram.memory\[126\]\[1\] _06036_ _06039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14178__S _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15542_ _01313_ net3 mod.u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12754_ _03872_ _05576_ _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _05262_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15394__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15473_ _01247_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12685_ _03944_ _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08118__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14424_ _00278_ net3 mod.u_cpu.rf_ram.memory\[475\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11636_ _04821_ _05214_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07246__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14355_ _00209_ net3 mod.u_cpu.rf_ram.memory\[510\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11567_ _05178_ mod.u_cpu.rf_ram.memory\[272\]\[1\] _05184_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10518_ _04472_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13306_ _06387_ _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14286_ _00140_ net3 mod.u_cpu.rf_ram.memory\[544\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11498_ _05139_ _05125_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13237_ _06342_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10449_ _04423_ mod.u_cpu.rf_ram.memory\[450\]\[0\] _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12225__I _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09794__I0 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13590__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13168_ _06276_ mod.u_cpu.rf_ram.memory\[349\]\[1\] _06274_ _06277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _05550_ mod.u_cpu.rf_ram.memory\[210\]\[1\] _05560_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12161__S _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13099_ _06230_ mod.u_cpu.rf_ram.memory\[102\]\[0\] _06234_ _06235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07660_ mod.u_cpu.rf_ram.memory\[303\]\[0\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12058__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07591_ _01879_ mod.u_cpu.rf_ram.memory\[366\]\[0\] _01898_ _01867_ _01899_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11105__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14611__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09330_ _03546_ _03576_ _03577_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07989__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11805__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09474__A2 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _03506_ _03515_ _03519_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08212_ _01489_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] _03464_
+ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14761__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _02152_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12230__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12081__I1 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09709__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ _01483_ _02336_ _02381_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_174_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15117__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07229__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__A1 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13730__A1 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13730__B2 _06736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15267__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _03251_ _03280_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08488__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07927_ _02157_ _02234_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12297__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _01765_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14038__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14291__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07789_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07899__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13797__B2 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09528_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07476__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _03395_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11272__A2 _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12470_ _05709_ _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11421_ _01950_ _05085_ _05086_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14140_ _07057_ mod.u_cpu.rf_ram.memory\[289\]\[0\] _07058_ _07059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11352_ _05032_ mod.u_cpu.rf_ram.memory\[307\]\[1\] _05039_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__A3 _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10303_ _04325_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14071_ _05630_ _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11283_ _04993_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07139__I _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13022_ _06184_ mod.u_cpu.rf_ram.memory\[10\]\[1\] _06182_ _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08728__A1 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10234_ _04248_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10535__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11583__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07400__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10165_ _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A2 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14973_ _00827_ net3 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14634__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13924_ _04067_ _06030_ _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14029__A2 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13855_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_arbiter.i_wb_cpu_rdt\[6\] _06335_
+ _06849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12806_ _05226_ _05320_ _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14784__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13786_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06774_ _06788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10998_ _04796_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09700__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15525_ _01296_ net3 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12460__A1 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12737_ _03865_ _05552_ _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11263__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12460__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15456_ _01230_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12668_ _05936_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14201__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14407_ _00261_ net3 mod.u_cpu.rf_ram.memory\[484\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10963__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11015__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11619_ _05208_ mod.u_cpu.rf_ram.memory\[263\]\[1\] _05218_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15387_ _01162_ net3 mod.u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__I3 mod.u_cpu.rf_ram.memory\[315\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11060__S _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12599_ _05873_ _05891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14338_ _00192_ net3 mod.u_cpu.rf_ram.memory\[518\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14269_ _00123_ net3 mod.u_cpu.rf_ram.memory\[553\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A1 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13712__A1 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__I3 mod.u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08814__S1 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09392__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _02410_ mod.u_cpu.rf_ram.memory\[22\]\[1\] _03136_ _01830_ _03137_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08761_ _03056_ _03058_ _02149_ _03067_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07712_ _01993_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_66_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10203__I _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08692_ _02348_ _02998_ _02377_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09695__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07643_ _01949_ _01950_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13079__I0 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07574_ _01749_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09313_ _03413_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12451__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11034__I _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08750__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09244_ _03496_ mod.u_scanchain_local.module_data_in\[39\] _03497_ _03504_ _03408_
+ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_90_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09175_ mod.u_arbiter.i_wb_cpu_rdt\[15\] _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12203__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14507__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _02365_ _02426_ _02433_ _02168_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12754__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08057_ _02347_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09758__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13554__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14657__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11565__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07233__I1 mod.u_cpu.rf_ram.memory\[457\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07933__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ _03254_ mod.u_cpu.cpu.decode.opcode\[1\] _03263_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11317__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10113__I _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11970_ _02203_ _05462_ _05463_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09686__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09902__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10921_ _04739_ mod.u_cpu.rf_ram.memory\[374\]\[1\] _04742_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11145__S _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13424__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13640_ _03297_ _03681_ _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10852_ _04290_ _04687_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13571_ _06605_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _04650_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15310_ _00071_ net4 mod.u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12522_ _05840_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14195__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15241_ _01094_ net3 mod.u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12453_ _03289_ _03667_ _05791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13242__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15432__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12745__A2 _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13942__A1 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__I _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11404_ _05071_ mod.u_cpu.rf_ram.memory\[298\]\[0\] _05075_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15172_ _01025_ net3 mod.u_cpu.rf_ram.memory\[148\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12384_ _03864_ _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _04196_ _03752_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14123_ _07043_ mod.u_cpu.rf_ram.memory\[116\]\[0\] _07047_ _07048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14054_ _07001_ _07002_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11266_ _04976_ mod.u_cpu.rf_ram.memory\[320\]\[1\] _04979_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11556__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15582__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _04249_ mod.u_cpu.rf_ram.memory\[486\]\[0\] _04264_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13170__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _06173_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _06163_ _06174_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11197_ _04933_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11181__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10148_ _04186_ _04213_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10079_ _04163_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14956_ _00810_ net3 mod.u_cpu.rf_ram.memory\[217\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09921__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08856__C _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13907_ _06647_ _06661_ _06682_ _06861_ _06888_ _06889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_78_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14887_ _00741_ net3 mod.u_cpu.rf_ram.memory\[240\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13334__I _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13838_ _03331_ _03404_ _01424_ _03334_ _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12433__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__S _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13769_ _03670_ _03396_ _06771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15508_ _01279_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08732__S0 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07290_ _01561_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08591__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15439_ _01214_ net3 mod.u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__I _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08163__I _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09195__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _03873_ _04062_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13697__B1 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11547__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09862_ _04001_ mod.u_cpu.rf_ram.memory\[53\]\[0\] _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07915__A2 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08813_ mod.u_cpu.rf_ram.memory\[8\]\[1\] mod.u_cpu.rf_ram.memory\[9\]\[1\] mod.u_cpu.rf_ram.memory\[10\]\[1\]
+ mod.u_cpu.rf_ram.memory\[11\]\[1\] _02171_ _02267_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _03889_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14110__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08744_ _02933_ _02965_ _01481_ _03050_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08675_ mod.u_cpu.rf_ram.memory\[215\]\[1\] _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10868__I _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15305__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10522__I1 mod.u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A2 mod.u_cpu.rf_ram.memory\[508\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _01710_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07242__I mod.u_cpu.raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07557_ mod.u_cpu.rf_ram.memory\[383\]\[0\] _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08723__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__S1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15455__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07488_ mod.u_cpu.rf_ram.memory\[439\]\[0\] _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14177__A1 _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ _03371_ _03489_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07851__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09158_ _03446_ _03435_ _03447_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13924__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ _02150_ _02404_ _02416_ _02363_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07603__A1 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10108__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03388_ _03389_ mod.u_cpu.cpu.state.o_cnt_r\[2\]
+ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_163_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _04620_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11538__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _04825_ mod.u_cpu.rf_ram.memory\[354\]\[1\] _04832_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10002_ _03928_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__I1 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14810_ _00664_ net3 mod.u_cpu.rf_ram.memory\[282\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14741_ _00595_ net3 mod.u_cpu.rf_ram.memory\[317\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11953_ _05452_ _05423_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07580__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13154__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10904_ _03803_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14672_ _00526_ net3 mod.u_cpu.rf_ram.memory\[351\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11884_ _05403_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13623_ _06581_ mod.u_cpu.rf_ram.memory\[309\]\[1\] _06636_ _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12415__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10835_ _04679_ mod.u_cpu.rf_ram.memory\[387\]\[0\] _04684_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08692__B _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13554_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] mod.u_arbiter.i_wb_cpu_dbus_adr\[12\]
+ _06594_ _06596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10766_ _04218_ _04623_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09292__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09831__A2 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10977__A1 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14168__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12505_ _05829_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12018__I1 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14822__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10697_ _04592_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13485_ _06549_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13915__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15224_ _01077_ net3 mod.u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13915__B2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12436_ _05776_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08398__A2 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15155_ _01008_ net3 mod.u_cpu.rf_ram.memory\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12367_ _05695_ _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13757__C _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__I _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14972__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14106_ _07026_ _07036_ _07037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11318_ _05017_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15086_ _00940_ net3 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12298_ _05679_ mod.u_cpu.rf_ram.memory\[187\]\[0\] _05683_ _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11529__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__A1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14037_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] _06989_ _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11249_ _04905_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09347__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07327__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10201__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15328__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14939_ _00793_ net3 mod.u_cpu.rf_ram.memory\[223\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07490__C _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11457__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11701__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14352__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__S1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08460_ _01956_ _02766_ _01788_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15478__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07411_ _01550_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08391_ _02191_ mod.u_cpu.rf_ram.memory\[422\]\[1\] _02697_ _02323_ _02698_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14096__S _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11513__S _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07342_ _01643_ mod.u_cpu.rf_ram.memory\[494\]\[0\] _01649_ _01615_ _01650_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12957__A2 _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07273_ _01523_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09012_ _03312_ _03287_ _03314_ _03315_ _03316_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__13906__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12709__A2 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__B _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09914_ _03851_ _04038_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09889__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07237__I _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08010__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _04001_ mod.u_cpu.rf_ram.memory\[542\]\[0\] _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _03948_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ mod.u_cpu.rf_ram.memory\[247\]\[1\] _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07747__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08658_ _02944_ _02964_ _01738_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ mod.u_cpu.rf_ram.memory\[312\]\[0\] mod.u_cpu.rf_ram.memory\[313\]\[0\] mod.u_cpu.rf_ram.memory\[314\]\[0\]
+ mod.u_cpu.rf_ram.memory\[315\]\[0\] _01774_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14845__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ _01496_ mod.u_cpu.rf_ram.memory\[268\]\[1\] _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11423__S _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12948__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _04541_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10551_ _04493_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07824__A1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14995__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13270_ _06120_ _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10482_ _04307_ _04447_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13373__A2 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ _05630_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13912__A4 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10187__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11384__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12152_ _05584_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14225__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__C _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10982__I1 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11103_ _04864_ mod.u_cpu.rf_ram.memory\[346\]\[0\] _04870_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09329__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12053__I _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12083_ _05533_ mod.u_cpu.rf_ram.memory\[212\]\[1\] _05536_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _04703_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08001__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14375__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15620__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12636__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12985_ _06113_ _03370_ _06158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14724_ _00578_ net3 mod.u_cpu.rf_ram.memory\[325\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11936_ mod.u_cpu.rf_ram.memory\[169\]\[1\] _05230_ _05439_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12239__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14655_ _00509_ net3 mod.u_cpu.rf_ram.memory\[360\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _05391_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13606_ _01429_ _03307_ _03315_ _06625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08068__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _04663_ mod.u_cpu.rf_ram.memory\[390\]\[0\] _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14586_ _00440_ net3 mod.u_cpu.rf_ram.memory\[394\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07610__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11798_ _05343_ _05335_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07815__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13537_ _06586_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10749_ _04627_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15000__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07291__A2 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13468_ _06512_ _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15207_ _01060_ net3 mod.u_cpu.rf_ram.memory\[209\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13364__A2 _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12419_ mod.u_cpu.rf_ram.memory\[489\]\[1\] _05765_ _05763_ _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13399_ _06310_ _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08240__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15138_ _00991_ net3 mod.u_cpu.rf_ram.memory\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15150__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ mod.u_cpu.rf_ram.memory\[248\]\[0\] mod.u_cpu.rf_ram.memory\[249\]\[0\] mod.u_cpu.rf_ram.memory\[250\]\[0\]
+ mod.u_cpu.rf_ram.memory\[251\]\[0\] _02266_ _02267_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15069_ _00923_ net3 mod.u_cpu.rf_ram.memory\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12175__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14718__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07891_ mod.u_cpu.rf_ram.memory\[219\]\[0\] _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11922__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A2 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _03835_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09561_ _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14868__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08512_ mod.u_cpu.rf_ram.memory\[349\]\[1\] _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09492_ _03716_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08443_ _01680_ _02749_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12339__S _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _02148_ _02680_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ _01494_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07256_ _01545_ mod.u_cpu.rf_ram.memory\[478\]\[0\] _01563_ _01525_ _01564_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14248__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07187_ _01494_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14398__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15643__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11913__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09828_ _03749_ _03818_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09759_ _03937_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13633__S _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08298__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__I _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12770_ _04955_ _05952_ _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _05289_ mod.u_cpu.rf_ram.memory\[243\]\[0\] _05290_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13418__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11153__S _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14440_ _00294_ net3 mod.u_cpu.rf_ram.memory\[467\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15023__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11652_ _05242_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07430__I _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10603_ _04527_ _04528_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14371_ _00225_ net3 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11583_ _05180_ mod.u_cpu.rf_ram.memory\[26\]\[0\] _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13322_ _03664_ _06416_ _06339_ _06418_ _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10534_ _04482_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__A1 _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15173__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11887__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ _03755_ _04132_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13253_ _06351_ mod.u_cpu.rf_ram.memory\[95\]\[0\] _06352_ _06353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10404__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12204_ _05605_ mod.u_cpu.rf_ram.memory\[200\]\[0\] _05619_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08222__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13184_ _05783_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _06290_ _06291_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10396_ _04389_ _03896_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A2 _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12135_ _05559_ mod.u_cpu.rf_ram.memory\[74\]\[0\] _05572_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12066_ _05518_ mod.u_cpu.rf_ram.memory\[29\]\[1\] _05525_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12857__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08525__A2 _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _04810_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08081__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11380__I1 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11127__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13543__S _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08289__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12968_ _06142_ _06143_ _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14707_ _00561_ net3 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08384__S1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11919_ _05428_ _05423_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10966__I _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11063__S _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12899_ _03985_ _06048_ _06089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14638_ _00492_ net3 mod.u_cpu.rf_ram.memory\[368\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15516__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14569_ _00423_ net3 mod.u_cpu.rf_ram.memory\[403\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _01418_ mod.u_cpu.cpu.csr_imm _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ mod.u_cpu.rf_ram.memory\[31\]\[0\] _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11797__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14540__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__I _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08992_ _03251_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07943_ _02180_ _02250_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12848__A1 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14690__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12421__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07874_ _02180_ _02181_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09613_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09544_ _03756_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15046__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12320__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09475_ _01500_ _03700_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08426_ mod.u_cpu.rf_ram.memory\[400\]\[1\] mod.u_cpu.rf_ram.memory\[401\]\[1\] mod.u_cpu.rf_ram.memory\[402\]\[1\]
+ mod.u_cpu.rf_ram.memory\[403\]\[1\] _02688_ _02475_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10882__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13025__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14073__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15196__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08127__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08357_ _01890_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _01577_ mod.u_cpu.rf_ram.memory\[510\]\[0\] _01613_ _01615_ _01616_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ mod.u_cpu.rf_ram.memory\[456\]\[1\] mod.u_cpu.rf_ram.memory\[457\]\[1\] mod.u_cpu.rf_ram.memory\[458\]\[1\]
+ mod.u_cpu.rf_ram.memory\[459\]\[1\] _02593_ _02594_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13328__A2 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07239_ _01520_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10250_ _04287_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09952__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14128__I1 mod.u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08014__C _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08755__A2 mod.u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10181_ _04238_ _04234_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12839__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13427__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__A2 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09704__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13940_ _03434_ _06912_ _06914_ _06915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13871_ _06840_ _06859_ _06860_ _06863_ _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15610_ _01381_ net3 mod.u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12822_ _06018_ _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14413__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15541_ _01312_ net3 mod.u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15539__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12753_ _05962_ _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ _05278_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10873__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15472_ _01246_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12684_ _03895_ _05589_ _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07160__I _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14423_ _00277_ net3 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08118__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11635_ _05231_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14563__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14354_ _00208_ net3 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08443__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11566_ _05185_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13305_ _06402_ _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _04467_ mod.u_cpu.rf_ram.memory\[440\]\[1\] _04470_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14285_ _00139_ net3 mod.u_cpu.rf_ram.memory\[545\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11497_ _03789_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_171_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13236_ _06273_ mod.u_cpu.rf_ram.memory\[94\]\[0\] _06341_ _06342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10448_ _04281_ _04407_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__I1 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13167_ _06236_ _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10379_ _03894_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_151_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12118_ _05561_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13098_ _03950_ _06223_ _06234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12241__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12049_ _03770_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15069__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07335__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07590_ _01663_ _01897_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12058__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13007__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09260_ _03516_ mod.u_scanchain_local.module_data_in\[41\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08682__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14906__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08211_ _02471_ _02508_ _02517_ _02518_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09191_ _03467_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _02209_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_147_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__I3 mod.u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ _02337_ _02346_ _02379_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10919__I1 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13730__A2 _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09725__I _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ mod.u_cpu.cpu.decode.co_mem_word _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07926_ mod.u_cpu.rf_ram.memory\[229\]\[0\] _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13494__B2 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14436__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _02161_ mod.u_cpu.rf_ram.memory\[198\]\[0\] _02163_ _02164_ _02165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07173__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__B _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13246__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07788_ _01686_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09527_ _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14586__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07476__A2 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08673__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09458_ mod.u_cpu.cpu.bufreg.c_r _03684_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08409_ mod.u_cpu.rf_ram.memory\[447\]\[1\] _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09389_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_178_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11420_ _05022_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08425__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__I3 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _05040_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10302_ _04313_ mod.u_cpu.rf_ram.memory\[474\]\[1\] _04323_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14070_ _03483_ _06911_ _06919_ _07012_ _07013_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _04976_ mod.u_cpu.rf_ram.memory\[318\]\[1\] _04991_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09925__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13021_ _06104_ _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08728__A2 _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10233_ _04275_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15211__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10164_ _03992_ _04134_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10095_ _03761_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14972_ _00826_ net3 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08036__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07155__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10299__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13923_ _06641_ _06899_ _06900_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07164__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15361__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11606__S _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13854_ _06847_ _06848_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14929__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12805_ _06026_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13785_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _06753_ _06786_ _06787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09456__A3 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15524_ _01295_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12736_ _05981_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08664__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__A1 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15455_ _01229_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12667_ _05934_ mod.u_cpu.rf_ram.memory\[121\]\[0\] _05935_ _05936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14406_ _00260_ net3 mod.u_cpu.rf_ram.memory\[484\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11618_ _02015_ _05218_ _05219_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_156_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15386_ _01161_ net3 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12598_ _05890_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__A1 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14337_ _00191_ net3 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__A2 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12236__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11549_ _05162_ mod.u_cpu.rf_ram.memory\[275\]\[1\] _05172_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14309__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A2 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14268_ _00122_ net3 mod.u_cpu.rf_ram.memory\[553\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13219_ _06317_ _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13712__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14199_ _03389_ mod.u_cpu.cpu.state.o_cnt\[2\] _07096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14459__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ _02631_ _03059_ _03066_ _02363_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12523__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09144__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ _01956_ _02011_ _02018_ _01989_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08691_ mod.u_cpu.rf_ram.memory\[200\]\[1\] mod.u_cpu.rf_ram.memory\[201\]\[1\] mod.u_cpu.rf_ram.memory\[202\]\[1\]
+ mod.u_cpu.rf_ram.memory\[203\]\[1\] _02349_ _02350_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07642_ mod.u_cpu.rf_ram.memory\[295\]\[0\] _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13079__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09280__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07573_ _01663_ _01880_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ _03557_ _03558_ _03560_ _03561_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08655__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12451__A2 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _03503_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08750__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08407__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09174_ _03457_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08125_ _02405_ _02429_ _02432_ _02415_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15234__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08056_ _02348_ _02351_ _02362_ _02363_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09907__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13703__A2 _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08499__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09383__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15384__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08958_ mod.u_cpu.cpu.decode.opcode\[2\] mod.u_cpu.cpu.decode.opcode\[0\] mod.u_cpu.cpu.decode.opcode\[1\]
+ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07909_ _02216_ mod.u_cpu.rf_ram.memory\[208\]\[0\] _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08889_ mod.u_cpu.rf_ram.memory\[560\]\[1\] mod.u_cpu.rf_ram.memory\[561\]\[1\] mod.u_cpu.rf_ram.memory\[562\]\[1\]
+ mod.u_cpu.rf_ram.memory\[563\]\[1\] _02457_ _02473_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10920_ _04743_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10851_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08646__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13570_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] mod.u_arbiter.i_wb_cpu_dbus_adr\[19\]
+ _06604_ _06605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10782_ _04637_ mod.u_cpu.rf_ram.memory\[396\]\[0\] _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12521_ _05827_ mod.u_cpu.rf_ram.memory\[166\]\[0\] _05839_ _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15240_ _01093_ net3 mod.u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12452_ _03394_ _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10056__I1 mod.u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11253__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _04792_ _05058_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15171_ _01024_ net3 mod.u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12056__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12383_ _05741_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11953__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14122_ _03842_ _05631_ _07047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11334_ _04960_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14601__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09749__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14053_ mod.u_arbiter.i_wb_cpu_rdt\[26\] _06998_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11265_ _04980_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13004_ _01453_ _06172_ _03370_ _06173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10216_ _04262_ _04263_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11196_ _04916_ mod.u_cpu.rf_ram.memory\[331\]\[1\] _04931_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13816__S _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11181__A2 _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10304__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _04068_ _04173_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14751__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14955_ _00809_ net3 mod.u_cpu.rf_ram.memory\[539\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10078_ _04142_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11336__S _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13906_ _06065_ _06490_ _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08885__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14886_ _00740_ net3 mod.u_cpu.rf_ram.memory\[240\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13837_ _06340_ _06832_ _06833_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15107__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13768_ _03674_ _06769_ _06770_ _06411_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08637__A1 _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13630__A1 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15507_ _01278_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12719_ _05970_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08732__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13699_ _03364_ _06704_ _06707_ _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15257__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15438_ _01213_ net3 mod.u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12197__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13933__A2 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15369_ _01144_ net3 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14281__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09930_ _04002_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13697__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13697__B2 _06705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04013_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ mod.u_cpu.rf_ram.memory\[12\]\[1\] mod.u_cpu.rf_ram.memory\[13\]\[1\] mod.u_cpu.rf_ram.memory\[14\]\[1\]
+ mod.u_cpu.rf_ram.memory\[15\]\[1\] _02266_ _02388_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_98_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10214__I _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ _03963_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _02992_ _03011_ _03049_ _02148_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14110__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08674_ _02479_ mod.u_cpu.rf_ram.memory\[212\]\[1\] _02980_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07679__A2 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07625_ mod.u_cpu.rf_ram.memory\[304\]\[0\] mod.u_cpu.rf_ram.memory\[305\]\[0\] mod.u_cpu.rf_ram.memory\[306\]\[0\]
+ mod.u_cpu.rf_ram.memory\[307\]\[0\] _01802_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07556_ _01671_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08628__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13621__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10884__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08723__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07487_ _01728_ mod.u_cpu.rf_ram.memory\[436\]\[0\] _01794_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09226_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14177__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14624__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09157_ mod.u_arbiter.i_wb_cpu_rdt\[8\] _03436_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12983__I0 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08108_ _02405_ _02409_ _02414_ _02415_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08039_ _01630_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13688__A1 _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09185__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12735__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14774__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11050_ _04833_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09356__A2 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09600__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _02529_ _04109_ _04110_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09913__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07861__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14740_ _00594_ net3 mod.u_cpu.rf_ram.memory\[317\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11952_ _03795_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08867__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13860__A1 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__I _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10903_ _04731_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14671_ _00525_ net3 mod.u_cpu.rf_ram.memory\[352\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11883_ _05385_ mod.u_cpu.rf_ram.memory\[227\]\[0\] _05402_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13622_ _01935_ _06636_ _06637_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10834_ _04277_ _04669_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12415__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13553_ _06595_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11474__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09292__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _04621_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10977__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12504_ _05827_ mod.u_cpu.rf_ram.memory\[16\]\[0\] _05828_ _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14168__A2 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13484_ _03605_ _06545_ _06546_ _03610_ _06549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10696_ _04584_ mod.u_cpu.rf_ram.memory\[410\]\[0\] _04591_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15223_ _01076_ net3 mod.u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11226__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13915__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12435_ mod.u_cpu.rf_ram.memory\[173\]\[1\] _05765_ _05774_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11926__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11777__I1 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15154_ _01007_ net3 mod.u_cpu.rf_ram.memory\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _05730_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14105_ _03836_ _05720_ _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11317_ _05007_ mod.u_cpu.rf_ram.memory\[312\]\[0\] _05016_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15085_ _00939_ net3 mod.u_cpu.rf_ram.memory\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12297_ _05139_ _05668_ _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08213__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11529__I1 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07608__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14036_ _06914_ _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11248_ _04968_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11179_ _04921_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08867__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14938_ _00792_ net3 mod.u_cpu.rf_ram.memory\[223\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08858__A1 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07343__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11701__I1 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10665__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14869_ _00723_ net3 mod.u_cpu.rf_ram.memory\[255\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _01703_ _01708_ _01715_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08375__S _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _02272_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07341_ _01647_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14647__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09283__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10968__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07272_ _01578_ _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09011_ mod.u_cpu.cpu.bufreg.lsb\[0\] _03292_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_176_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11217__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13906__A2 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09035__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14797__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07597__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10440__I1 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07518__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12342__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09844_ _03752_ _04003_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08777__C _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14095__A1 _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13255__I _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08726_ _02161_ mod.u_cpu.rf_ram.memory\[244\]\[1\] _03032_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08349__I _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08849__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15422__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13842__A1 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13842__B2 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08657_ _02104_ _02963_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _01581_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08588_ mod.u_cpu.rf_ram.memory\[269\]\[1\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_169_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _01836_ _01846_ _01485_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15572__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11503__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10550_ _04481_ mod.u_cpu.rf_ram.memory\[434\]\[1\] _04491_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09209_ _03477_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11208__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10119__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _04436_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12220_ _05629_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A1 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11384__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12151_ _05583_ mod.u_cpu.rf_ram.memory\[207\]\[1\] _05580_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08880__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08033__B _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11102_ _04868_ _04869_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12082_ _05537_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12333__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08968__B mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _03959_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07591__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12984_ _06157_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12636__A2 _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11935_ _05440_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14723_ _00577_ net3 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11614__S _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14654_ _00508_ net3 mod.u_cpu.rf_ram.memory\[360\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11866_ _05383_ mod.u_cpu.rf_ram.memory\[70\]\[1\] _05389_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13605_ _03362_ _03354_ _06624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _04262_ _04669_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08068__A2 _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14585_ _00439_ net3 mod.u_cpu.rf_ram.memory\[395\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11797_ _03931_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] mod.u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _06584_ _06586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07815__A2 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _04626_ mod.u_cpu.rf_ram.memory\[402\]\[1\] _04624_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13467_ _06537_ _06538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10679_ _04307_ _04570_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15206_ _01059_ net3 mod.u_cpu.rf_ram.memory\[209\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12418_ _05229_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09568__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13398_ _06285_ _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15137_ _00990_ net3 mod.u_cpu.rf_ram.memory\[429\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12349_ _05718_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07338__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15068_ _00922_ net3 mod.u_cpu.rf_ram.memory\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14019_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _06976_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _06977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07890_ _02197_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08623__S0 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15445__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09553__I _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11922__I1 mod.u_cpu.rf_ram.memory\[222\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14077__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13124__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _03749_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08169__I _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ mod.u_cpu.rf_ram.memory\[350\]\[1\] mod.u_cpu.rf_ram.memory\[351\]\[1\] _01664_
+ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11686__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09491_ mod.u_cpu.rf_ram_if.wen1_r mod.u_cpu.rf_ram_if.wen0_r _01418_ _03717_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07503__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15595__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13803__I _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08442_ mod.u_cpu.rf_ram.memory\[392\]\[1\] mod.u_cpu.rf_ram.memory\[393\]\[1\] mod.u_cpu.rf_ram.memory\[394\]\[1\]
+ mod.u_cpu.rf_ram.memory\[395\]\[1\] _02020_ _02748_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07801__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11438__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08373_ _01591_ _02653_ _02679_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09256__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07255_ _01561_ _01562_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__I0 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07186_ mod.u_cpu.raddr\[0\] _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12563__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07248__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08614__S0 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12866__A2 _06066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _03989_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10877__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14812__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08300__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09758_ _03936_ mod.u_cpu.rf_ram.memory\[552\]\[1\] _03934_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08709_ _02594_ _03012_ _03015_ _02764_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09689_ _03862_ mod.u_cpu.rf_ram.memory\[55\]\[1\] _03880_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09495__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11434__S _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11720_ _05037_ _05284_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14962__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13418__I1 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11429__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _05234_ mod.u_cpu.rf_ram.memory\[24\]\[1\] _05240_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09839__S _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10602_ _03892_ _04225_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_14370_ _00224_ net3 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11582_ _05110_ _03797_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13321_ _06417_ _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15318__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10533_ _04481_ mod.u_cpu.rf_ram.memory\[437\]\[1\] _04479_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08470__A2 _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12929__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13252_ _04984_ _06344_ _06352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10464_ _04434_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12203_ _05343_ _05611_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13183_ _03500_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_135_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10395_ _03727_ _03807_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__14342__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15468__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _05334_ _05543_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07981__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12065_ _02395_ _05525_ _05526_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11016_ _04803_ mod.u_cpu.rf_ram.memory\[35\]\[0\] _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14492__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13806__B2 _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12967_ _03338_ _03375_ _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14706_ _00560_ net3 mod.u_cpu.rf_ram.memory\[334\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11293__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11918_ _03750_ _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10340__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12898_ _06072_ _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07621__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14637_ _00491_ net3 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11849_ _05366_ mod.u_cpu.rf_ram.memory\[149\]\[0\] _05378_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10891__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09749__S _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14568_ _00422_ net3 mod.u_cpu.rf_ram.memory\[403\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12093__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13519_ _06568_ _03691_ _06572_ _06573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10643__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14499_ _00353_ net3 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09548__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__I _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09410__A1 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _03260_ _03294_ _03295_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14835__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07942_ mod.u_cpu.rf_ram.memory\[239\]\[0\] _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10859__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ mod.u_cpu.rf_ram.memory\[207\]\[0\] _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07724__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _03821_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14985__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09543_ _03765_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09477__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13533__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09474_ _01418_ _01645_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08425_ _02687_ _02723_ _02731_ _01678_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_169_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09229__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13025__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ _02631_ _02662_ _01618_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07307_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08287_ _02030_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14365__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07238_ mod.u_cpu.rf_ram.memory\[463\]\[0\] _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15610__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12536__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08204__A2 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07169_ _01477_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _03910_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07963__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__S _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12839__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11228__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13870_ _06861_ _06862_ _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12821_ _06037_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15540_ _01311_ net3 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12752_ _05991_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07441__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11703_ _05271_ mod.u_cpu.rf_ram.memory\[252\]\[1\] _05276_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15140__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15471_ _01245_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12683_ _05946_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14422_ _00276_ net3 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14708__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11634_ mod.u_cpu.rf_ram.memory\[261\]\[1\] _05230_ _05227_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14353_ _00207_ net3 mod.u_cpu.rf_ram.memory\[511\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13972__B1 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11822__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11565_ _05180_ mod.u_cpu.rf_ram.memory\[272\]\[0\] _05184_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08443__A2 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13304_ _06118_ _06300_ _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15290__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10516_ _04471_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14284_ _00138_ net3 mod.u_cpu.rf_ram.memory\[545\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ _05138_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12527__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14858__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13235_ _03751_ _06193_ _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10447_ _04347_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13166_ _06275_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10378_ _04376_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07954__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12117_ _05559_ mod.u_cpu.rf_ram.memory\[210\]\[0\] _05560_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10243__S _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13097_ _06233_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07616__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12048_ _05514_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13781__C _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14238__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13999_ _06960_ _06961_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13353__I _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10313__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07351__I mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13007__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14388__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08210_ _02291_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12066__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09190_ mod.u_arbiter.i_wb_cpu_rdt\[21\] mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] _03464_
+ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15633__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ _02124_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13302__B _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11813__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08434__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__I0 mod.u_cpu.rf_ram.memory\[440\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _01485_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08198__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__A1 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08974_ mod.u_cpu.cpu.bufreg.lsb\[0\] _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15013__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ mod.u_cpu.rf_ram.memory\[224\]\[0\] mod.u_cpu.rf_ram.memory\[225\]\[0\] mod.u_cpu.rf_ram.memory\[226\]\[0\]
+ mod.u_cpu.rf_ram.memory\[227\]\[0\] _02151_ _02172_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _01820_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07173__A2 _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15163__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _02090_ _02094_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09526_ _03745_ _03749_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09170__I0 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09457_ _03356_ _03680_ _03682_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _02462_ mod.u_cpu.rf_ram.memory\[444\]\[1\] _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11009__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _03606_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_61_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08339_ _02421_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11350_ _05028_ mod.u_cpu.rf_ram.memory\[307\]\[0\] _05039_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11280__I1 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12509__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ _04324_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08025__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11281_ _04992_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13020_ _06183_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10232_ _04267_ mod.u_cpu.rf_ram.memory\[484\]\[1\] _04273_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09925__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10163_ _04223_ _04224_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09852__S _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ _01597_ _04174_ _04175_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14971_ _00825_ net3 mod.u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15506__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13922_ _06166_ _06649_ _06900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07164__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13853_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[2\]
+ _06848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12804_ _06019_ mod.u_cpu.rf_ram.memory\[128\]\[1\] _06024_ _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14530__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13784_ _06065_ _06783_ _06785_ _06786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07171__I mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10996_ _03761_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15523_ _01294_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09456__A4 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12735_ _05966_ mod.u_cpu.rf_ram.memory\[136\]\[1\] _05979_ _05981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09861__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__A2 mod.u_cpu.rf_ram.memory\[222\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12718__S _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15454_ _01228_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12666_ _05896_ _05721_ _05935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12748__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14405_ _00259_ net3 mod.u_cpu.rf_ram.memory\[485\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14680__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11617_ _05133_ _05218_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__I _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12597_ _05887_ mod.u_cpu.rf_ram.memory\[155\]\[0\] _05889_ _05890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15385_ _01160_ net3 mod.u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10223__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11420__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14336_ _00190_ net3 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11548_ _05173_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13549__S _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14267_ _00121_ net3 mod.u_cpu.rf_ram.memory\[554\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11479_ _05114_ mod.u_cpu.rf_ram.memory\[286\]\[0\] _05126_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15036__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13173__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13218_ _06307_ _06315_ _06319_ _06324_ _06325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14198_ _07076_ _03320_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07927__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12920__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13149_ _06265_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12771__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10782__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15186__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07710_ _01961_ _02014_ _02017_ _02005_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08690_ _02578_ _02993_ _02996_ _02660_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08352__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09561__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07641_ _01758_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07572_ mod.u_cpu.rf_ram.memory\[375\]\[0\] _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07538__S0 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _03486_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08655__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _03502_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09173_ _03456_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] _03452_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ _02410_ mod.u_cpu.rf_ram.memory\[38\]\[0\] _02431_ _01828_ _02432_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_147_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ _01586_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13164__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09368__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14403__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15529__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08957_ mod.u_cpu.cpu.decode.co_ebreak _01423_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11478__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07908_ _01681_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10525__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08888_ _02449_ _03187_ _03194_ _02505_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14553__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09471__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07839_ _02103_ _02146_ _01475_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14089__I _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _04620_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12278__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09509_ _03733_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10781_ _04233_ _04648_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08646__A2 _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12520_ _05355_ _05831_ _05839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10453__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07859__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12451_ _03700_ _05788_ _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10058__S _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12337__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15059__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11402_ _05074_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15170_ _01023_ net3 mod.u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12382_ _05729_ mod.u_cpu.rf_ram.memory\[178\]\[1\] _05739_ _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__A2 _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14121_ _07046_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11953__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ _05027_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14052_ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] _07000_ _07001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11264_ _04978_ mod.u_cpu.rf_ram.memory\[320\]\[0\] _04979_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07909__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13003_ _01435_ _01420_ _01424_ _06172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10215_ _04136_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11195_ _04932_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07166__I _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08582__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10146_ _04212_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14954_ _00808_ net3 mod.u_cpu.rf_ram.memory\[539\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10077_ _04025_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08334__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13905_ _06481_ _06660_ _06887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14885_ _00739_ net3 mod.u_cpu.rf_ram.memory\[241\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13836_ mod.u_cpu.cpu.immdec.imm30_25\[5\] _06774_ _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13767_ _06764_ _03391_ _06416_ _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10979_ _04783_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15506_ _01277_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12718_ _05966_ mod.u_cpu.rf_ram.memory\[138\]\[1\] _05968_ _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13698_ _06421_ _06706_ _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15437_ _01212_ net3 mod.u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12649_ _05924_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13394__A1 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12197__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15368_ _01143_ net3 mod.u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14426__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14319_ _00173_ net3 mod.u_cpu.rf_ram.memory\[528\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15299_ _00059_ net4 mod.u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09860_ _03836_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14576__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ mod.u_cpu.rf_ram.memory\[0\]\[1\] mod.u_cpu.rf_ram.memory\[1\]\[1\] mod.u_cpu.rf_ram.memory\[2\]\[1\]
+ mod.u_cpu.rf_ram.memory\[3\]\[1\] _02211_ _02386_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09791_ _03958_ mod.u_cpu.rf_ram.memory\[548\]\[0\] _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _01848_ _03029_ _03048_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07128__A2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08673_ _02202_ _02979_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ _01827_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07555_ _01862_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15201__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ _01774_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12680__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13909__B1 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09225_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09156_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08107_ _01765_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15351__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10994__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09466__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14919__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14185__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08370__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _02339_ _02341_ _02343_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13688__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10000_ _03899_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08564__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__A2 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09989_ _04091_ mod.u_cpu.rf_ram.memory\[51\]\[1\] _04100_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13716__I _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08316__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10123__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11951_ _05451_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13860__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11236__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ _04720_ mod.u_cpu.rf_ram.memory\[377\]\[1\] _04729_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14670_ _00524_ net3 mod.u_cpu.rf_ram.memory\[352\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11882_ _04965_ _05401_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13621_ _06249_ _06636_ _06637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10833_ _04683_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11172__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11623__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13552_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] mod.u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _06594_ _06595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08545__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12671__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10764_ _04636_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14449__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12503_ _05563_ _03873_ _05828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13483_ _06548_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10695_ _04322_ _04575_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12434_ _02112_ _05774_ _05775_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15222_ _01075_ net3 mod.u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12423__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11226__I1 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11926__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15153_ _01006_ net3 mod.u_cpu.rf_ram.memory\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12365_ _05729_ mod.u_cpu.rf_ram.memory\[180\]\[1\] _05727_ _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14599__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09376__I _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _04732_ _05011_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14104_ _07035_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15084_ _00938_ net3 mod.u_cpu.rf_ram.memory\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12296_ _05682_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13679__A2 _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14035_ _06986_ _06988_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _04952_ mod.u_cpu.rf_ram.memory\[323\]\[1\] _04966_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08555__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11178_ _04916_ mod.u_cpu.rf_ram.memory\[334\]\[1\] _04919_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10362__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10129_ _03858_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14937_ _00791_ net3 mod.u_cpu.rf_ram.memory\[224\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08858__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13851__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10665__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15224__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14868_ _00722_ net3 mod.u_cpu.rf_ram.memory\[255\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13819_ _06363_ _06465_ _06668_ _06779_ _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14799_ _00653_ net3 mod.u_cpu.rf_ram.memory\[288\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08166__S0 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07340_ mod.u_cpu.rf_ram.memory\[495\]\[0\] _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_189_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07271_ mod.u_cpu.rf_ram.memory\[471\]\[0\] _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15374__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09010_ _01428_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07597__A2 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09912_ _03738_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10728__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08546__A1 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12342__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09774_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14095__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08725_ _02197_ _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11153__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13842__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ _02105_ _02953_ _02962_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11853__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07607_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ mod.u_cpu.rf_ram.memory\[270\]\[1\] mod.u_cpu.rf_ram.memory\[271\]\[1\] _02106_
+ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08365__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07538_ _01839_ _01840_ _01842_ _01845_ _01832_ _01833_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11605__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07469_ _01728_ mod.u_cpu.rf_ram.memory\[428\]\[0\] _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12816__S _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13358__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] _03474_
+ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14741__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _04446_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12405__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A2 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12150_ _05549_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _04847_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14891__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12551__S _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12081_ _05521_ mod.u_cpu.rf_ram.memory\[212\]\[0\] _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10719__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11032_ _04820_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12333__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10344__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11392__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13446__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08632__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15247__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07444__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12097__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12983_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie mod.u_cpu.cpu.genblk3.csr.mstatus_mpie
+ _06143_ _06157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08984__B _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14722_ _00576_ net3 mod.u_cpu.rf_ram.memory\[326\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11934_ mod.u_cpu.rf_ram.memory\[169\]\[0\] _05437_ _05439_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14271__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14653_ _00507_ net3 mod.u_cpu.rf_ram.memory\[361\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15397__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _05390_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13604_ _06623_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10816_ _04672_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11796_ _05310_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14584_ _00438_ net3 mod.u_cpu.rf_ram.memory\[395\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08208__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13535_ _06585_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10747_ _04578_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13349__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10678_ _04580_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13466_ _06509_ _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09017__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15205_ _01058_ net3 mod.u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12417_ _05764_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__I0 mod.u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13397_ _06478_ _06479_ _06481_ _06491_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10958__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15136_ _00989_ net3 mod.u_cpu.rf_ram.memory\[429\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12348_ _05713_ mod.u_cpu.rf_ram.memory\[181\]\[0\] _05717_ _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15067_ _00921_ net3 mod.u_cpu.rf_ram.memory\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12279_ _05671_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09834__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14018_ _06963_ _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08878__C _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14077__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14614__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08510_ _02664_ _02807_ _02816_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09490_ _03664_ _03715_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07503__A2 _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08700__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _01762_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08372_ _02661_ _02663_ _02664_ _02678_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14764__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11438__I1 mod.u_cpu.rf_ram.memory\[292\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07323_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07267__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12260__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07254_ mod.u_cpu.rf_ram.memory\[479\]\[0\] _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07957__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07185_ _01492_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08767__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13760__A1 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12563__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08614__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13266__I _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09826_ _03964_ mod.u_cpu.rf_ram.memory\[544\]\[1\] _03987_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07264__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14294__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _03889_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11826__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ _02209_ _03013_ _03014_ _02633_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ _03881_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09495__A2 _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ mod.u_cpu.rf_ram.memory\[173\]\[1\] _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08095__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _05241_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11429__I1 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _03713_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11581_ _05195_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13320_ _06313_ _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10532_ _04429_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10463_ _04430_ mod.u_cpu.rf_ram.memory\[448\]\[1\] _04432_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13251_ _06204_ _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07439__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08758__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13751__A1 _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12202_ _05618_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13182_ _06288_ _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13751__B2 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ _04388_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10565__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12133_ _05571_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12064_ _05488_ _05525_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14637__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _04808_ _03969_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08930__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14787__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12966_ _01425_ _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14705_ _00559_ net3 mod.u_cpu.rf_ram.memory\[335\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11917_ _05427_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__I1 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12897_ _06087_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14636_ _00490_ net3 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11848_ _04014_ _05374_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12242__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13290__I0 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14567_ _00421_ net3 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11779_ _04930_ _05301_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08836__I2 mod.u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09829__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13518_ _03685_ _03690_ _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_158_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14498_ _00352_ net3 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13449_ _06527_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13042__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07349__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15412__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13742__A1 _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15119_ _00972_ net3 mod.u_cpu.rf_ram.memory\[449\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10704__S _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _03278_ _03293_ _03267_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07941_ _01539_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15562__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__C _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07872_ _01778_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09611_ _03818_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09542_ _03764_ mod.u_cpu.rf_ram.memory\[574\]\[1\] _03759_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09721__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__B1 _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11334__I _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08424_ _02611_ _02726_ _02729_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08355_ mod.u_cpu.rf_ram.memory\[488\]\[1\] mod.u_cpu.rf_ram.memory\[489\]\[1\] mod.u_cpu.rf_ram.memory\[490\]\[1\]
+ mod.u_cpu.rf_ram.memory\[491\]\[1\] _02385_ _02633_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07968__B _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07306_ _01523_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _02116_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_20_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07237_ _01516_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12165__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13033__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15092__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07259__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12536__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ _01447_ _01459_ _01466_ _01476_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__10547__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07963__A2 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__C _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08912__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09809_ _03958_ mod.u_cpu.rf_ram.memory\[546\]\[0\] _03976_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09960__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12820_ _06035_ mod.u_cpu.rf_ram.memory\[126\]\[0\] _06036_ _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07722__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12751_ _05984_ mod.u_cpu.rf_ram.memory\[199\]\[1\] _05989_ _05991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08771__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11702_ _05277_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15470_ _01244_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12682_ _05938_ mod.u_cpu.rf_ram.memory\[142\]\[1\] _05944_ _05946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14421_ _00275_ net3 mod.u_cpu.rf_ram.memory\[477\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11633_ _05229_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14352_ _00206_ net3 mod.u_cpu.rf_ram.memory\[511\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15435__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11822__I1 mod.u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11564_ _04766_ _05171_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13303_ _06130_ _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10515_ _04469_ mod.u_cpu.rf_ram.memory\[440\]\[0\] _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14283_ _00137_ net3 mod.u_cpu.rf_ram.memory\[546\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11495_ _05128_ mod.u_cpu.rf_ram.memory\[284\]\[1\] _05136_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07169__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13724__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09779__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ _04422_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13234_ _06280_ _06340_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15585__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10377_ _04363_ mod.u_cpu.rf_ram.memory\[462\]\[1\] _04374_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13165_ _06273_ mod.u_cpu.rf_ram.memory\[349\]\[0\] _06274_ _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07954__A2 _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ _05293_ _05471_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13096_ _06217_ mod.u_cpu.rf_ram.memory\[59\]\[1\] _06231_ _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12047_ _05501_ mod.u_cpu.rf_ram.memory\[213\]\[1\] _05512_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08903__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13998_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _06952_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12949_ mod.u_cpu.cpu.genblk1.align.ctrl_misal _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13570__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08762__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14619_ _00473_ net3 mod.u_cpu.rf_ram.memory\[378\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12186__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15599_ _01370_ net3 mod.u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08140_ _01469_ _02281_ _02447_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09092__B1 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08071_ _02149_ _02364_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13015__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14802__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10529__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11577__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__A2 _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13191__A2 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14952__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _03256_ _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07924_ _01977_ _02187_ _02231_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ _01819_ _02162_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15308__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10701__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ mod.u_cpu.rf_ram.memory\[184\]\[0\] mod.u_cpu.rf_ram.memory\[185\]\[0\] mod.u_cpu.rf_ram.memory\[186\]\[0\]
+ mod.u_cpu.rf_ram.memory\[187\]\[0\] _02092_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _03746_ _03747_ _03748_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_25_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11501__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14332__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09456_ _03365_ mod.u_cpu.cpu.bufreg.c_r _03680_ _03682_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__15458__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08407_ _02111_ _02713_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09387_ _03624_ _03620_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ mod.u_cpu.rf_ram.memory\[509\]\[1\] _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09622__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14482__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _02551_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _04298_ mod.u_cpu.rf_ram.memory\[474\]\[0\] _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12509__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11280_ _04978_ mod.u_cpu.rf_ram.memory\[318\]\[0\] _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13719__I _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _04274_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12623__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _03662_ _03753_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10093_ _04044_ _04174_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14970_ _00824_ net3 mod.u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13921_ _06456_ _06468_ _06861_ _06452_ _06481_ _06899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13852_ _06842_ _06846_ _06483_ _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12803_ _06025_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13783_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _06455_ _06784_ _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10995_ _04794_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15522_ _01293_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12734_ _05980_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__A2 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14198__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15453_ _01227_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14825__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12665_ _05886_ _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14404_ _00258_ net3 mod.u_cpu.rf_ram.memory\[485\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12748__A2 _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11616_ _04539_ _05130_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15384_ _01159_ net3 mod.u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12596_ _05888_ _05882_ _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14335_ _00189_ net3 mod.u_cpu.rf_ram.memory\[520\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11547_ _05159_ mod.u_cpu.rf_ram.memory\[275\]\[0\] _05172_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11420__A2 _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14975__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14266_ _00120_ net3 mod.u_cpu.rf_ram.memory\[554\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11478_ _04852_ _05125_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13629__I _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13217_ _06321_ _06323_ _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13173__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10429_ _04411_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14197_ _07095_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12920__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13148_ mod.u_arbiter.i_wb_cpu_rdt\[25\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _06263_ _06265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09047__C _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11149__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10782__I1 mod.u_cpu.rf_ram.memory\[396\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10053__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14122__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13079_ mod.u_cpu.rf_ram.memory\[105\]\[1\] _06221_ _06219_ _06222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12684__A1 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11085__S _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__A2 _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14355__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ _01643_ mod.u_cpu.rf_ram.memory\[292\]\[0\] _01947_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07786__S1 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07362__I _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15600__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07571_ _01710_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11813__S _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__S1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09310_ _03549_ _03559_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09241_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13236__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12708__I _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09289__I mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09172_ mod.u_arbiter.i_wb_cpu_rdt\[14\] _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12739__A2 _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ _02411_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10228__I _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ _02352_ _02355_ _02360_ _02361_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09368__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13164__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12443__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11175__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15130__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08591__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ mod.u_arbiter.i_wb_cpu_dbus_we _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09752__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09915__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07907_ mod.u_cpu.rf_ram.memory\[209\]\[0\] _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10898__I _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08887_ _02455_ _03190_ _03193_ _02467_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10525__I1 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A2 mod.u_cpu.rf_ram.memory\[510\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07838_ _02104_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15280__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12427__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07769_ _01677_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14848__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09508_ _03732_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10780_ _04569_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09439_ _03331_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12450_ _05780_ mod.u_cpu.cpu.state.stage_two_req _05787_ _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14998__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11401_ _05069_ mod.u_cpu.rf_ram.memory\[2\]\[1\] _05072_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12381_ _05740_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14120_ _07041_ mod.u_cpu.rf_ram.memory\[11\]\[1\] _07044_ _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11332_ _05014_ mod.u_cpu.rf_ram.memory\[310\]\[1\] _05025_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14228__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07875__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09359__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14051_ _06914_ _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12353__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11263_ _04838_ _04969_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A2 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13002_ _06167_ _06164_ _06171_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08031__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _03950_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11194_ _04918_ mod.u_cpu.rf_ram.memory\[331\]\[0\] _04931_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11961__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _04199_ mod.u_cpu.rf_ram.memory\[496\]\[1\] _04210_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14378__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15623__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14953_ _00807_ net3 mod.u_cpu.rf_ram.memory\[529\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10076_ _04147_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12666__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13904_ _06707_ _06886_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10601__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08278__I _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14884_ _00738_ net3 mod.u_cpu.rf_ram.memory\[241\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07182__I mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13835_ mod.u_cpu.cpu.immdec.imm7 _03682_ _06812_ _06831_ _06832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_46_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13766_ mod.u_cpu.cpu.immdec.imm7 _06753_ _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10978_ mod.u_cpu.rf_ram.memory\[365\]\[1\] _04661_ _04781_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07910__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13630__A3 _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15505_ _01276_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12717_ _05969_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13697_ _06694_ _06431_ _06450_ _06705_ _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15003__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15436_ _01211_ net3 mod.u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12648_ _05923_ mod.u_cpu.rf_ram.memory\[147\]\[1\] _05921_ _05924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15367_ _01142_ net3 mod.u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12579_ _05877_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14318_ _00172_ net3 mod.u_cpu.rf_ram.memory\[528\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15298_ _00058_ net4 mod.u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15153__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12263__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14249_ _00103_ net3 mod.u_cpu.rf_ram.memory\[563\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11157__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07357__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ mod.u_cpu.rf_ram.memory\[4\]\[1\] mod.u_cpu.rf_ram.memory\[5\]\[1\] mod.u_cpu.rf_ram.memory\[6\]\[1\]
+ mod.u_cpu.rf_ram.memory\[7\]\[1\] _02366_ _02383_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _03948_ _03961_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08741_ _01978_ _03038_ _03047_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09522__A1 _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08672_ mod.u_cpu.rf_ram.memory\[213\]\[1\] _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07623_ _01915_ _01917_ _01930_ _01812_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13082__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07554_ _01509_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07485_ mod.u_cpu.rf_ram.memory\[437\]\[0\] _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07836__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13909__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10691__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09224_ _03384_ _03486_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09155_ _03445_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09747__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08106_ _02410_ mod.u_cpu.rf_ram.memory\[22\]\[0\] _02413_ _01830_ _02414_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09086_ _03386_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13269__I _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _01493_ _02344_ _01534_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14520__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15646__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11943__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _04101_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _01464_ _01465_ _03206_ _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_69_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14670__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08316__A2 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11950_ _05450_ mod.u_cpu.rf_ram.memory\[21\]\[1\] _05447_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08098__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10123__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10901_ _04730_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11881_ _05262_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13620_ _05164_ _04989_ _06636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15026__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10832_ _04682_ mod.u_cpu.rf_ram.memory\[388\]\[1\] _04680_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13551_ _06583_ _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_186_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10069__S _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10763_ _04626_ mod.u_cpu.rf_ram.memory\[3\]\[1\] _04634_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12502_ _05812_ _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10682__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13482_ _03602_ _06545_ _06546_ _03605_ _06548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14168__A4 _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10694_ _04590_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15176__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15221_ _01074_ net3 mod.u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12433_ _05642_ _05774_ _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15152_ _01005_ net3 mod.u_cpu.rf_ram.memory\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12364_ _05710_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14103_ _07028_ mod.u_cpu.rf_ram.memory\[110\]\[1\] _07033_ _07035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11315_ _05015_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15083_ _00937_ net3 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12295_ _05677_ mod.u_cpu.rf_ram.memory\[188\]\[1\] _05680_ _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07177__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14034_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _06987_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11246_ _04967_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12887__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12811__I _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11177_ _04920_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10128_ _04200_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08307__A2 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10331__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10059_ _04151_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14936_ _00790_ net3 mod.u_cpu.rf_ram.memory\[224\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14867_ _00721_ net3 mod.u_cpu.rf_ram.memory\[256\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13818_ _06814_ _06816_ _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13064__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14798_ _00652_ net3 mod.u_cpu.rf_ram.memory\[288\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12111__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08166__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13749_ _06335_ _03428_ _06754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15519__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10673__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07270_ _01560_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08491__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15419_ _01194_ net3 mod.u_cpu.rf_ram.memory\[349\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14543__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08471__I _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09991__A1 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10506__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12178__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09911_ _04049_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14693__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09842_ _03994_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09773_ _03856_ _03939_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08724_ mod.u_cpu.rf_ram.memory\[245\]\[1\] _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10241__I _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15049__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12350__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _02124_ _02954_ _02961_ _02143_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11853__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _01850_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _01978_ _02883_ _02892_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07550__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12102__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15199__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ mod.u_cpu.rf_ram.memory\[336\]\[0\] mod.u_cpu.rf_ram.memory\[337\]\[0\] mod.u_cpu.rf_ram.memory\[338\]\[0\]
+ mod.u_cpu.rf_ram.memory\[339\]\[0\] _01843_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_169_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11605__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ _01774_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _03476_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13358__A2 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07399_ _01567_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10416__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ _03431_ _03387_ _03432_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__I _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10041__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__A2 _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09069_ _01433_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11100_ _03795_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12080_ _05535_ _05471_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11916__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10719__I1 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11031_ mod.u_cpu.rf_ram.memory\[357\]\[1\] _04819_ _04816_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10352__S _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11392__I1 mod.u_cpu.rf_ram.memory\[300\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13294__A1 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12097__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12982_ _06146_ _06155_ _06156_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14721_ _00575_ net3 mod.u_cpu.rf_ram.memory\[327\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14416__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11933_ _05078_ _05438_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_73_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14652_ _00506_ net3 mod.u_cpu.rf_ram.memory\[361\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11864_ _05385_ mod.u_cpu.rf_ram.memory\[70\]\[0\] _05389_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07460__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13603_ mod.u_cpu.rf_ram.memory\[329\]\[1\] _06221_ _06621_ _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13597__A2 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ _04666_ mod.u_cpu.rf_ram.memory\[391\]\[1\] _04670_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14583_ _00437_ net3 mod.u_cpu.rf_ram.memory\[396\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11795_ _05341_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10655__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14566__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13534_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] mod.u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _06584_ _06585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10746_ _04625_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10280__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13465_ _06536_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _04579_ mod.u_cpu.rf_ram.memory\[414\]\[1\] _04576_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15204_ _01057_ net3 mod.u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12416_ mod.u_cpu.rf_ram.memory\[489\]\[0\] _05622_ _05763_ _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13396_ _06483_ _06489_ _06490_ _06491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15135_ _00988_ net3 mod.u_cpu.rf_ram.memory\[469\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11080__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12347_ _04014_ _05703_ _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15066_ _00920_ net3 mod.u_cpu.rf_ram.memory\[186\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12278_ _05660_ mod.u_cpu.rf_ram.memory\[191\]\[1\] _05669_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14017_ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] _06966_ _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11229_ _04107_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12580__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10996__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12189__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14919_ _00773_ net3 mod.u_cpu.rf_ram.memory\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15341__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13372__I _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10894__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08440_ _02143_ _02744_ _02746_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08700__A2 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14909__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07370__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I0 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _02665_ _02667_ _02676_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _01490_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15491__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08464__A1 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12260__A2 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07253_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12399__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07184_ _01491_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08134__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12571__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09825_ _03988_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14439__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11067__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09756_ _03935_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10900__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12323__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08707_ _02385_ mod.u_cpu.rf_ram.memory\[236\]\[1\] _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _03877_ mod.u_cpu.rf_ram.memory\[55\]\[0\] _03880_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11826__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13291__A4 _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14589__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08638_ mod.u_cpu.rf_ram.memory\[168\]\[1\] mod.u_cpu.rf_ram.memory\[169\]\[1\] mod.u_cpu.rf_ram.memory\[170\]\[1\]
+ mod.u_cpu.rf_ram.memory\[171\]\[1\] _02106_ _02127_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08569_ mod.u_cpu.rf_ram.memory\[277\]\[1\] _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10600_ _04526_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07258__A2 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08455__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11580_ _05194_ mod.u_cpu.rf_ram.memory\[270\]\[1\] _05192_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09201__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08845__I3 mod.u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10531_ _01793_ _04479_ _04480_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__S _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _06350_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13200__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10462_ _04433_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12201_ mod.u_cpu.rf_ram.memory\[201\]\[1\] _05617_ _05615_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08758__A2 mod.u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13181_ _06286_ _06287_ _06288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13751__A2 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ _04387_ mod.u_cpu.rf_ram.memory\[460\]\[1\] _04385_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10565__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15214__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12132_ _05566_ mod.u_cpu.rf_ram.memory\[208\]\[1\] _05569_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09707__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13457__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12063_ _04983_ _03771_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11014_ _04250_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15364__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12965_ _06135_ _06141_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11705__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08286__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11916_ _05426_ mod.u_cpu.rf_ram.memory\[223\]\[1\] _05424_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14704_ _00558_ net3 mod.u_cpu.rf_ram.memory\[335\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12896_ _06086_ mod.u_cpu.rf_ram.memory\[98\]\[1\] _06084_ _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07190__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14635_ _00489_ net3 mod.u_cpu.rf_ram.memory\[370\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__C _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11847_ _05377_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14566_ _00420_ net3 mod.u_cpu.rf_ram.memory\[404\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11778_ _05330_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08836__I3 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13517_ _03425_ _06570_ _06571_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10729_ _04613_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14497_ _00351_ net3 mod.u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13448_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _06525_ _06526_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A1 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08749__A2 _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13742__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13379_ _06454_ _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11753__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15118_ _00971_ net3 mod.u_cpu.rf_ram.memory\[449\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07972__A3 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07940_ _02244_ mod.u_cpu.rf_ram.memory\[236\]\[0\] _02247_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15049_ _00903_ net3 mod.u_cpu.rf_ram.memory\[195\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11505__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07871_ _01646_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10859__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09610_ _03746_ _03819_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13258__A1 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14731__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09541_ _03763_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09721__I1 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09472_ _03697_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12481__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08423_ _01914_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14881__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _02654_ _02655_ _02659_ _02660_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08437__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13430__A1 _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07968__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07305_ _01578_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12446__I _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08988__A2 _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _02591_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11992__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15237__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07236_ _01508_ mod.u_cpu.rf_ram.memory\[460\]\[0\] _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13033__I1 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07167_ _01469_ _01471_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11744__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14261__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15387__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12544__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09808_ _03948_ _03975_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _03890_ mod.u_cpu.rf_ram.memory\[554\]\[1\] _03920_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09712__I1 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12750_ _02162_ _05989_ _05990_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08676__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10483__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11701_ _05268_ mod.u_cpu.rf_ram.memory\[252\]\[0\] _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08771__S1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12681_ _05945_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14420_ _00274_ net3 mod.u_cpu.rf_ram.memory\[477\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11632_ _03733_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12224__A2 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07878__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14351_ _00205_ net3 mod.u_cpu.rf_ram.memory\[512\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13972__A2 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11563_ _05183_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13302_ _06366_ _06376_ _06381_ _06399_ _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10514_ _04168_ _04464_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14282_ _00136_ net3 mod.u_cpu.rf_ram.memory\[546\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11494_ _05137_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13233_ _06325_ _06333_ _06336_ _06339_ _06340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13724__A2 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10445_ _04410_ mod.u_cpu.rf_ram.memory\[451\]\[1\] _04420_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13164_ _05515_ _04969_ _06274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08600__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ _04375_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12091__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12115_ _05520_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13095_ _06232_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07185__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14754__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12046_ _02226_ _05512_ _05513_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12160__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08903__A2 mod.u_cpu.rf_ram.memory\[516\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13997_ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] _06954_ _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12948_ _06122_ _06123_ _06124_ _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08762__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12879_ _06070_ mod.u_cpu.rf_ram.memory\[246\]\[1\] _06074_ _06076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14618_ _00472_ net3 mod.u_cpu.rf_ram.memory\[378\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13412__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15598_ _01369_ net3 mod.u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11274__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14549_ _00403_ net3 mod.u_cpu.rf_ram.memory\[413\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12266__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09092__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09092__B2 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11974__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08070_ _02365_ _02368_ _02376_ _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14284__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10529__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11726__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11577__I1 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08442__I1 mod.u_cpu.rf_ram.memory\[393\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08412__C _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07309__B _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ _03268_ _03270_ _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07923_ _02195_ _02208_ _02229_ _02230_ _01978_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07158__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07854_ mod.u_cpu.rf_ram.memory\[199\]\[0\] _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10701__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _02042_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _03709_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08658__A1 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13651__A1 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09455_ _03349_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13560__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08406_ mod.u_cpu.rf_ram.memory\[445\]\[1\] _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13403__A1 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07698__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14627__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08337_ mod.u_cpu.rf_ram.memory\[504\]\[1\] mod.u_cpu.rf_ram.memory\[505\]\[1\] mod.u_cpu.rf_ram.memory\[506\]\[1\]
+ mod.u_cpu.rf_ram.memory\[507\]\[1\] _02385_ _02633_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_177_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08268_ mod.u_cpu.rf_ram.memory\[543\]\[0\] _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07633__A2 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _01490_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12904__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _02209_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_152_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__B _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14777__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10230_ _04249_ mod.u_cpu.rf_ram.memory\[484\]\[0\] _04273_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10161_ _04222_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_161_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10092_ _04172_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13920_ _06898_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07733__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13851_ _06451_ _06672_ _06844_ _06845_ _06846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11255__I _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12802_ _06010_ mod.u_cpu.rf_ram.memory\[128\]\[0\] _06024_ _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13782_ _03509_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _06784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08649__A1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10994_ _04774_ mod.u_cpu.rf_ram.memory\[362\]\[0\] _04793_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15402__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15521_ _01292_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12733_ _05963_ mod.u_cpu.rf_ram.memory\[136\]\[0\] _05979_ _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15452_ _01226_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12664_ _05933_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14403_ _00257_ net3 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11615_ _05217_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15552__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15383_ _01158_ net3 mod.u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12595_ _03789_ _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14334_ _00188_ net3 mod.u_cpu.rf_ram.memory\[520\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11546_ _05037_ _05171_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14265_ _00119_ net3 mod.u_cpu.rf_ram.memory\[555\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11477_ _05124_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11708__A1 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13216_ _06322_ _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _04410_ mod.u_cpu.rf_ram.memory\[454\]\[1\] _04408_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14196_ _06057_ _03388_ _07095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_152_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08232__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13147_ _06264_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _04363_ mod.u_cpu.rf_ram.memory\[465\]\[1\] _04361_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13078_ _03734_ _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12029_ _05239_ _03851_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08888__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10695__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07570_ _01875_ mod.u_cpu.rf_ram.memory\[372\]\[0\] _01877_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15082__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11495__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07312__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09240_ _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13397__B1 _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11247__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09171_ _03455_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07311__C _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09065__A1 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11947__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08122_ mod.u_cpu.rf_ram.memory\[39\]\[0\] _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07615__A2 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08053_ _01528_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08955_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07981__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07906_ _02209_ _02210_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ _02461_ mod.u_cpu.rf_ram.memory\[574\]\[1\] _03192_ _02465_ _03193_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08879__A1 _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13872__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15425__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07837_ _02105_ _02123_ _02144_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12427__A2 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ _02074_ _02075_ _01602_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09507_ _01462_ _03352_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10289__I1 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15575__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07303__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _01787_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09438_ _03668_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09369_ _03568_ _03607_ _03608_ _03609_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11400_ _05073_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12380_ _05731_ mod.u_cpu.rf_ram.memory\[178\]\[0\] _05739_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08803__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11331_ _05026_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14050_ _06997_ _06999_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11262_ _04960_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08052__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13001_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _03353_ _06163_ _06170_ _06171_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10213_ _04261_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10154__I _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11193_ _04930_ _04926_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08031__A2 _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10144_ _04211_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10075_ _04161_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14952_ _00806_ net3 mod.u_cpu.rf_ram.memory\[529\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13863__A1 mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12666__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07463__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13863__B2 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13903_ _03355_ _06140_ _06886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14883_ _00737_ net3 mod.u_cpu.rf_ram.memory\[242\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13834_ _06651_ _06829_ _06830_ _03682_ _06831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13615__A1 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13765_ _06768_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10977_ _01894_ _04781_ _04782_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15504_ _01275_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12716_ _05963_ mod.u_cpu.rf_ram.memory\[138\]\[0\] _05968_ _05969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13696_ _06295_ _06306_ _06464_ _06682_ _06493_ _06323_ _06705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__14942__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13918__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15435_ _01210_ net3 mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09047__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12647_ _05873_ _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14040__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15366_ _01141_ net3 mod.u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12578_ _05869_ mod.u_cpu.rf_ram.memory\[158\]\[0\] _05876_ _05877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14317_ _00171_ net3 mod.u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11529_ _05159_ mod.u_cpu.rf_ram.memory\[278\]\[0\] _05160_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15297_ _00057_ net4 mod.u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12729__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14248_ _00102_ net3 mod.u_cpu.rf_ram.memory\[563\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12354__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13576__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11401__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14179_ _07084_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14322__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15448__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08897__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13375__I _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12106__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11096__S _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07781__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08740_ _03017_ _03039_ _03046_ _01870_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08405__S0 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13854__A1 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09522__A2 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14472__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08671_ _02606_ _02977_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15598__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__S _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07622_ _01918_ _01923_ _01928_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07553_ _01857_ mod.u_cpu.rf_ram.memory\[380\]\[0\] _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09286__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13082__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07484_ mod.u_cpu.rf_ram.memory\[432\]\[0\] mod.u_cpu.rf_ram.memory\[433\]\[0\] mod.u_cpu.rf_ram.memory\[434\]\[0\]
+ mod.u_cpu.rf_ram.memory\[435\]\[0\] _01745_ _01747_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07836__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08137__C _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09223_ _03406_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13909__A2 _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10840__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09154_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _03444_ _03442_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09589__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _02411_ _02412_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11640__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09085_ _03385_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08261__A2 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07548__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ mod.u_cpu.rf_ram.memory\[92\]\[0\] mod.u_cpu.rf_ram.memory\[93\]\[0\] mod.u_cpu.rf_ram.memory\[94\]\[0\]
+ mod.u_cpu.rf_ram.memory\[95\]\[0\] _01636_ _01638_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09987_ _04096_ mod.u_cpu.rf_ram.memory\[51\]\[0\] _04100_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14815__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08600__C _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ _01459_ _03225_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_153_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ _02542_ _03168_ _03175_ _02518_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_18_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10900_ _04728_ mod.u_cpu.rf_ram.memory\[377\]\[0\] _04729_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11880_ _05400_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14965__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09204__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _04640_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13550_ _06593_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10762_ _04635_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09003__I mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12501_ _05826_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13481_ _06547_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _04579_ mod.u_cpu.rf_ram.memory\[411\]\[1\] _04588_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15220_ _01073_ net3 mod.u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12432_ _05593_ _05438_ _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__I0 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07886__C _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11387__A2 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15151_ _01004_ net3 mod.u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12363_ _05728_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12364__I _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14345__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07458__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14102_ _07034_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11314_ _05014_ mod.u_cpu.rf_ram.memory\[313\]\[1\] _05012_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15082_ _00936_ net3 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12294_ _05681_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14033_ _06963_ _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11245_ _04961_ mod.u_cpu.rf_ram.memory\[323\]\[0\] _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10813__S _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12887__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11934__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ _04918_ mod.u_cpu.rf_ram.memory\[334\]\[0\] _04919_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14495__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10127_ _04199_ mod.u_cpu.rf_ram.memory\[4\]\[1\] _04197_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10058_ _04140_ mod.u_cpu.rf_ram.memory\[50\]\[1\] _04149_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11698__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14935_ _00789_ net3 mod.u_cpu.rf_ram.memory\[225\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14866_ _00720_ net3 mod.u_cpu.rf_ram.memory\[256\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13817_ _06423_ _06449_ _06459_ _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13064__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14797_ _00651_ net3 mod.u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12111__I1 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13748_ _06482_ _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15120__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13679_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _06678_ _06690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15418_ _01193_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12274__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15349_ _01124_ net3 mod.u_cpu.rf_ram.memory\[369\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15270__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09991__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14838__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09910_ _04036_ mod.u_cpu.rf_ram.memory\[532\]\[1\] _04047_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09841_ _03915_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10889__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09772_ _03766_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08199__I _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13827__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14988__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08723_ mod.u_cpu.rf_ram.memory\[240\]\[1\] mod.u_cpu.rf_ram.memory\[241\]\[1\] mod.u_cpu.rf_ram.memory\[242\]\[1\]
+ mod.u_cpu.rf_ram.memory\[243\]\[1\] _01647_ _01732_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_152_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07506__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _02110_ _02957_ _02960_ _02141_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07831__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07605_ _01835_ _01847_ _01912_ _01482_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12449__I _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08585_ _01992_ _02884_ _02891_ _02007_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07536_ _01503_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07467_ mod.u_cpu.rf_ram.memory\[429\]\[0\] _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14368__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] _03474_
+ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15613__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07398_ mod.u_cpu.rf_ram.memory\[413\]\[0\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09137_ mod.u_arbiter.i_wb_cpu_rdt\[3\] _03410_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07278__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09068_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11729__S _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08019_ _02298_ _02326_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S0 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__B _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11030_ _04531_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13118__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12981_ mod.u_cpu.cpu.genblk3.csr.mie_mtie _06155_ _06056_ _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11464__S _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14720_ _00574_ net3 mod.u_cpu.rf_ram.memory\[327\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09442__B _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11932_ _03892_ _05319_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07741__I _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15143__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12359__I _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14651_ _00505_ net3 mod.u_cpu.rf_ram.memory\[362\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11863_ _05355_ _05388_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13602_ _06622_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10814_ _04671_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10104__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11794_ mod.u_cpu.rf_ram.memory\[233\]\[1\] _05230_ _05339_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14582_ _00436_ net3 mod.u_cpu.rf_ram.memory\[396\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10804__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13533_ _06583_ _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10745_ _04622_ mod.u_cpu.rf_ram.memory\[402\]\[0\] _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09668__I _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15293__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10280__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13464_ _03574_ _06531_ _06532_ _03578_ _06536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10676_ _04578_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12415_ _05588_ _04228_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15203_ _01056_ net3 mod.u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10607__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13395_ _06310_ _06329_ _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07188__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15134_ _00987_ net3 mod.u_cpu.rf_ram.memory\[469\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12346_ _05716_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15065_ _00919_ net3 mod.u_cpu.rf_ram.memory\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12277_ _05670_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__S0 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14016_ _06973_ _06974_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11228_ _03924_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__S1 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10342__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11159_ _04908_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13285__A2 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14918_ _00772_ net3 mod.u_cpu.rf_ram.memory\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09352__B _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14849_ _00703_ net3 mod.u_cpu.rf_ram.memory\[263\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11048__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08370_ _01886_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14510__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15636__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__I1 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07321_ _01602_ _01621_ _01628_ _01587_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12796__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08464__A2 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07252_ mod.u_cpu.raddr\[0\] _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14660__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07183_ _01490_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09413__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08847__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15016__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12020__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07727__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11348__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09824_ _03958_ mod.u_cpu.rf_ram.memory\[544\]\[0\] _03987_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10582__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09755_ _03916_ mod.u_cpu.rf_ram.memory\[552\]\[0\] _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09024__S0 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15166__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12323__I1 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11287__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08706_ mod.u_cpu.rf_ram.memory\[237\]\[1\] _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09686_ _03878_ _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08152__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08637_ _02938_ _02943_ _02102_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12087__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ mod.u_cpu.rf_ram.memory\[272\]\[1\] mod.u_cpu.rf_ram.memory\[273\]\[1\] mod.u_cpu.rf_ram.memory\[274\]\[1\]
+ mod.u_cpu.rf_ram.memory\[275\]\[1\] _01957_ _01958_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07519_ _01700_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08499_ _02668_ _02802_ _02805_ _02096_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09488__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10530_ _04439_ _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10262__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13736__B1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ _04423_ mod.u_cpu.rf_ram.memory\[448\]\[0\] _04432_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10427__I _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09404__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13200__A2 _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08838__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12200_ _05229_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13180_ _05783_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _06287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10392_ _04344_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07966__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ _05570_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12642__I _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09707__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12062_ _05524_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15509__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11013_ _04807_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10573__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15821_ net4 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12964_ mod.u_cpu.cpu.ctrl.i_iscomp _06140_ _06141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14533__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07471__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14703_ _00557_ net3 mod.u_cpu.rf_ram.memory\[336\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _05405_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12895_ _06018_ _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14634_ _00488_ net3 mod.u_cpu.rf_ram.memory\[370\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11846_ _05364_ mod.u_cpu.rf_ram.memory\[159\]\[1\] _05375_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10628__I1 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14683__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13422__B net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14565_ _00419_ net3 mod.u_cpu.rf_ram.memory\[405\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11777_ _05329_ mod.u_cpu.rf_ram.memory\[236\]\[1\] _05326_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13516_ _03426_ _06570_ _06571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10728_ _04608_ mod.u_cpu.rf_ram.memory\[405\]\[1\] _04610_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14496_ _00350_ net3 mod.u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10659_ _04566_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13447_ _06513_ _06526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15039__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10005__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A2 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13378_ _06462_ _06467_ _06469_ _06473_ _06474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__12250__I0 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07957__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12950__A1 _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11753__A2 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15117_ _00970_ net3 mod.u_cpu.rf_ram.memory\[519\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12329_ _05696_ mod.u_cpu.rf_ram.memory\[184\]\[0\] _05704_ _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12002__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15048_ _00902_ net3 mod.u_cpu.rf_ram.memory\[195\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15189__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12702__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07870_ _02175_ mod.u_cpu.rf_ram.memory\[204\]\[0\] _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13258__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09540_ _03762_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10800__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08134__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07381__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_180 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14207__A1 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09882__A1 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__A2 _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08422_ _02692_ mod.u_cpu.rf_ram.memory\[414\]\[1\] _02728_ _01773_ _02729_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12069__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08353_ _01679_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__A2 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ mod.u_cpu.rf_ram.memory\[511\]\[0\] _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08284_ _01851_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09101__I _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ _01511_ _01542_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11992__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__I _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13194__A1 _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _01474_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14406__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11744__A2 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07556__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14556__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08373__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09807_ _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07999_ _02302_ mod.u_cpu.rf_ram.memory\[110\]\[0\] _02305_ _02306_ _02307_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10307__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09738_ _03921_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09173__I0 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _03855_ _03866_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11700_ _04859_ _05255_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10483__A2 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12680_ _05934_ mod.u_cpu.rf_ram.memory\[142\]\[0\] _05944_ _05945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11631_ _02012_ _05227_ _05228_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14350_ _00204_ net3 mod.u_cpu.rf_ram.memory\[512\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11562_ _05178_ mod.u_cpu.rf_ram.memory\[273\]\[1\] _05181_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11432__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _04452_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13301_ _06383_ _06362_ _06375_ _06396_ _06398_ _06399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_14281_ _00135_ net3 mod.u_cpu.rf_ram.memory\[547\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11493_ _05114_ mod.u_cpu.rf_ram.memory\[284\]\[0\] _05136_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13232_ _06338_ _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _04421_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13468__I _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15331__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13163_ _06204_ _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10375_ _04365_ mod.u_cpu.rf_ram.memory\[462\]\[0\] _04374_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08600__A2 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10794__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12114_ _05558_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13094_ _06230_ mod.u_cpu.rf_ram.memory\[59\]\[0\] _06231_ _06232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12045_ _05488_ _05512_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08364__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15481__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11716__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13996_ _06957_ _06959_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12947_ _03500_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _06124_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13931__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12878_ _06075_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14617_ _00471_ net3 mod.u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11829_ _05328_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13412__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15597_ _01368_ net3 mod.u_cpu.rf_ram.memory\[245\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11451__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14548_ _00402_ net3 mod.u_cpu.rf_ram.memory\[413\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14429__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11974__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14479_ _00333_ net3 mod.u_cpu.rf_ram.memory\[448\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12774__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14579__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ mod.u_cpu.cpu.bufreg2.i_cnt_done _03272_ _03273_ _03275_ _03276_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_130_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07922_ _01719_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07158__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09591__I _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _01646_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14002__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07784_ _02091_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09523_ _03271_ _03715_ _03705_ _01461_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13651__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _03255_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15204__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08405_ mod.u_cpu.rf_ram.memory\[440\]\[1\] mod.u_cpu.rf_ram.memory\[441\]\[1\] mod.u_cpu.rf_ram.memory\[442\]\[1\]
+ mod.u_cpu.rf_ram.memory\[443\]\[1\] _02711_ _01703_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09385_ _03563_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13403__A2 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ _02631_ _02634_ _02642_ _01587_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11414__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07713__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15354__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ _02546_ mod.u_cpu.rf_ram.memory\[540\]\[0\] _02574_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09766__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ _01517_ mod.u_cpu.rf_ram.memory\[454\]\[0\] _01522_ _01525_ _01526_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_165_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08198_ _02449_ _02496_ _02504_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_180_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10160_ mod.u_cpu.cpu.immdec.imm11_7\[4\] _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10091_ _04136_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10641__S _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08346__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13850_ _06472_ _06443_ _06466_ _06845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12801_ _03985_ _06011_ _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13781_ _06381_ _06372_ _06781_ _06782_ _06432_ _06783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10993_ _04792_ _04788_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15520_ _01291_ net3 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12732_ _03932_ _05978_ _05979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A2 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15451_ _01225_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12367__I _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12663_ _05923_ mod.u_cpu.rf_ram.memory\[144\]\[1\] _05931_ _05933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14402_ _00256_ net3 mod.u_cpu.rf_ram.memory\[486\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11614_ _05208_ mod.u_cpu.rf_ram.memory\[264\]\[1\] _05215_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15382_ _01157_ net3 mod.u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12594_ _05886_ _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14333_ _00187_ net3 mod.u_cpu.rf_ram.memory\[521\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11545_ _05124_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08821__A2 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09676__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14721__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14264_ _00118_ net3 mod.u_cpu.rf_ram.memory\[555\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11476_ _05118_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12905__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13215_ _06286_ _06287_ _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10427_ _04344_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14195_ _07076_ _07094_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07196__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08585__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _04344_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13146_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _06263_ _06264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14871__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13077_ _06220_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10289_ _04298_ mod.u_cpu.rf_ram.memory\[476\]\[0\] _04316_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08188__I1 mod.u_cpu.rf_ram.memory\[569\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12028_ _05502_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08888__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15227__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14130__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13979_ _06910_ _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14251__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15377__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ mod.u_arbiter.i_wb_cpu_rdt\[13\] mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _03452_
+ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13397__B2 _06491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08112__I1 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08121_ _02329_ mod.u_cpu.rf_ram.memory\[36\]\[0\] _02428_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11947__A2 _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ _02356_ mod.u_cpu.rf_ram.memory\[70\]\[0\] _02358_ _02359_ _02360_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10758__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08576__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12740__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08954_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07905_ _02211_ mod.u_cpu.rf_ram.memory\[210\]\[0\] _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08885_ _02500_ _03191_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13872__A2 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10260__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07836_ _02124_ _02128_ _02142_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_186_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07767_ mod.u_cpu.rf_ram.memory\[156\]\[0\] mod.u_cpu.rf_ram.memory\[157\]\[0\] mod.u_cpu.rf_ram.memory\[158\]\[0\]
+ mod.u_cpu.rf_ram.memory\[159\]\[0\] _01925_ _02071_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09828__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ _01462_ mod.u_cpu.rf_ram_if.wdata1_r\[1\] _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07698_ _01997_ _02001_ _02004_ _02005_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07303__A2 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ _03289_ _03667_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11091__I _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14744__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09368_ _03386_ mod.u_scanchain_local.module_data_in\[59\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_166_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08319_ _02198_ mod.u_cpu.rf_ram.memory\[470\]\[1\] _02625_ _01751_ _02626_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09299_ _03535_ mod.u_scanchain_local.module_data_in\[48\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_126_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11330_ _05007_ mod.u_cpu.rf_ram.memory\[310\]\[0\] _05025_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14188__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14894__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11261_ _04977_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08567__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10212_ _04245_ mod.u_cpu.rf_ram.memory\[487\]\[1\] _04259_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13000_ _06113_ _06166_ _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11410__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11192_ _03909_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10374__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _04193_ mod.u_cpu.rf_ram.memory\[496\]\[0\] _04210_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10371__S _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08319__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10074_ _04157_ mod.u_cpu.rf_ram.memory\[506\]\[1\] _04159_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14951_ _00805_ net3 mod.u_cpu.rf_ram.memory\[218\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13863__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13902_ _03359_ _06422_ _06693_ _06463_ _06699_ _06135_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_43_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14882_ _00736_ net3 mod.u_cpu.rf_ram.memory\[242\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10921__I0 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14274__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13833_ _06764_ _06829_ _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13764_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _06767_ _06709_ _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _04414_ _04781_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15503_ _01274_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07925__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12715_ _03918_ _05940_ _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08508__C _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13695_ _05787_ _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15434_ _01209_ net3 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12646_ _05922_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15365_ _01140_ net3 mod.u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12577_ _05428_ _05374_ _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10988__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14316_ _00170_ net3 mod.u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11528_ _04741_ _05149_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15296_ _00056_ net4 mod.u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12729__I1 mod.u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14247_ _00101_ net3 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11459_ _05112_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12354__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11401__I1 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14178_ _07057_ mod.u_cpu.rf_ram.memory\[8\]\[0\] _07083_ _07084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13129_ _06254_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12106__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07654__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08405__S1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11165__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14617__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08670_ _02759_ _02973_ _02976_ _01872_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08686__S _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14103__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08730__A1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07621_ _01686_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07552_ _01858_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11617__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14767__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ _01445_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _03435_ mod.u_scanchain_local.module_data_in\[37\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10840__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13090__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08104_ mod.u_cpu.rf_ram.memory\[23\]\[0\] _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _03384_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11640__I1 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08035_ _01662_ _02342_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12470__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09986_ _04013_ _03851_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14297__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08937_ _03234_ _03243_ _02520_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15542__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ _02455_ _03171_ _03174_ _02555_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_45_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08721__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13515__B _06569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07819_ _02126_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15433__D _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ mod.u_cpu.rf_ram.memory\[69\]\[1\] _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10830_ _04681_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07288__A1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10761_ _04622_ mod.u_cpu.rf_ram.memory\[3\]\[0\] _04634_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12500_ _05822_ mod.u_cpu.rf_ram.memory\[459\]\[1\] _05824_ _05826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10692_ _04589_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13480_ _03598_ _06545_ _06546_ _03602_ _06547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14022__A2 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12431_ _05773_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07739__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13781__A1 _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15150_ _01003_ net3 mod.u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12362_ _05713_ mod.u_cpu.rf_ram.memory\[180\]\[0\] _05727_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14101_ _07021_ mod.u_cpu.rf_ram.memory\[110\]\[0\] _07033_ _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10165__I _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ _04951_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15081_ _00935_ net3 mod.u_cpu.rf_ram.memory\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12293_ _05679_ mod.u_cpu.rf_ram.memory\[188\]\[0\] _05680_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15072__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14032_ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] _06978_ _06986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11244_ _04965_ _04945_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11395__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11175_ _04775_ _04906_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07474__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _04177_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07407__C _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13836__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04150_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14934_ _00788_ net3 mod.u_cpu.rf_ram.memory\[225\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11698__I1 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08712__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14865_ _00719_ net3 mod.u_cpu.rf_ram.memory\[250\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13816_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_arbiter.i_wb_cpu_rdt\[12\] _03510_
+ _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09268__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14796_ _00650_ net3 mod.u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13747_ _06752_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10959_ _04769_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10822__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13678_ _06421_ _06688_ _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15417_ _01192_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12629_ _05907_ mod.u_cpu.rf_ram.memory\[150\]\[1\] _05909_ _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07649__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15415__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15348_ _01123_ net3 mod.u_cpu.rf_ram.memory\[379\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15279_ _00037_ net4 mod.u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09864__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15565__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__C _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _04000_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09771_ _03947_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13827__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ _03016_ _03019_ _02074_ _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08653_ _02135_ mod.u_cpu.rf_ram.memory\[166\]\[1\] _02959_ _02139_ _02960_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14010__I _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07604_ _01848_ _01889_ _01911_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08584_ _01997_ _02887_ _02890_ _02005_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09104__I _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _01825_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ _01744_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ _03475_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15095__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13763__A1 _06761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ _03353_ _03369_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ mod.u_cpu.rf_ram.memory\[117\]\[0\] _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07993__A2 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07508__B _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07294__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14932__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ _04073_ mod.u_cpu.rf_ram.memory\[522\]\[0\] _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07227__C _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12980_ mod.u_cpu.cpu.decode.op22 _03343_ _06151_ _06154_ _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__12877__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13294__A3 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09215__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11931_ _03698_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09442__C _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10501__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14650_ _00504_ net3 mod.u_cpu.rf_ram.memory\[362\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12629__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11862_ _05387_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13601_ mod.u_cpu.rf_ram.memory\[329\]\[0\] _03899_ _06621_ _06622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _04663_ mod.u_cpu.rf_ram.memory\[391\]\[0\] _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12254__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14581_ _00435_ net3 mod.u_cpu.rf_ram.memory\[397\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10104__I1 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11301__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11793_ _05340_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14312__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15438__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13532_ _03292_ _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10744_ _04201_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13463_ _06535_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _04496_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09885__S _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15202_ _01055_ net3 mod.u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13754__A1 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12414_ _05762_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13394_ _06485_ _06488_ _06489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14462__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15588__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15133_ _00986_ net3 mod.u_cpu.rf_ram.memory\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12345_ _05711_ mod.u_cpu.rf_ram.memory\[182\]\[1\] _05714_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09684__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13506__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07984__A2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15064_ _00918_ net3 mod.u_cpu.rf_ram.memory\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _05662_ mod.u_cpu.rf_ram.memory\[191\]\[0\] _05669_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08608__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11719__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14015_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _06964_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11227_ _04953_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08933__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11158_ _04901_ mod.u_cpu.rf_ram.memory\[337\]\[0\] _04907_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10109_ _04186_ _04185_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11089_ _04843_ mod.u_cpu.rf_ram.memory\[348\]\[0\] _04860_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09489__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14917_ _00771_ net3 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13690__B1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14848_ _00702_ net3 mod.u_cpu.rf_ram.memory\[263\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13293__I0 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14779_ _00633_ net3 mod.u_cpu.rf_ram.memory\[298\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__I2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09859__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07320_ _01572_ _01624_ _01627_ _01584_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12796__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07251_ _01556_ mod.u_cpu.rf_ram.memory\[476\]\[0\] _01558_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13045__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14805__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07600__C _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07379__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07182_ mod.u_cpu.raddr\[2\] _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08847__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08712__B _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14955__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14170__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14005__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__I1 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09823_ _03767_ _03986_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09754_ _03902_ _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__S1 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07842__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08705_ mod.u_cpu.rf_ram.memory\[238\]\[1\] mod.u_cpu.rf_ram.memory\[239\]\[1\] _01807_
+ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11287__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _03822_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08152__A2 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14335__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08636_ _01836_ _02940_ _02942_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08567_ _01848_ _02854_ _02873_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_154_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10098__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08535__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07518_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _01875_ mod.u_cpu.rf_ram.memory\[334\]\[1\] _02804_ _02453_ _02805_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14485__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07449_ _01515_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13736__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _04290_ _04309_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13736__B2 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09404__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08838__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _03416_ _03392_ _03417_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10391_ _04386_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12923__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12130_ _05559_ mod.u_cpu.rf_ram.memory\[208\]\[0\] _05569_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12061_ _05518_ mod.u_cpu.rf_ram.memory\[62\]\[1\] _05522_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08915__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11012_ _04797_ mod.u_cpu.rf_ram.memory\[360\]\[1\] _04805_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15110__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__I1 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__A2 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12475__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12963_ _06139_ _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14702_ _00556_ net3 mod.u_cpu.rf_ram.memory\[336\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _05425_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15260__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12894_ _06085_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14633_ _00487_ net3 mod.u_cpu.rf_ram.memory\[371\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14828__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11845_ _05376_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14564_ _00418_ net3 mod.u_cpu.rf_ram.memory\[405\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _05328_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13515_ _03693_ _06568_ _06569_ _06570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_186_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10727_ _01725_ _04610_ _04612_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14495_ _00349_ net3 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13727__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14978__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13446_ _06510_ _06525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ _04557_ mod.u_cpu.rf_ram.memory\[416\]\[0\] _04565_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13377_ _06471_ _06464_ _06458_ _06395_ _06472_ _06473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_127_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _04238_ _04507_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15116_ _00969_ net3 mod.u_cpu.rf_ram.memory\[519\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07957__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12950__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12328_ _05283_ _05703_ _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10961__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15047_ _00901_ net3 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12259_ _03979_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12702__A2 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10713__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11761__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14358__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07662__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15603__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11513__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_170 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_181 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _03695_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14207__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09882__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08421_ _02244_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07893__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08352_ _02656_ _02657_ _02658_ _02067_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_51_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09634__A2 _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ _01607_ mod.u_cpu.rf_ram.memory\[508\]\[0\] _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08283_ _02561_ _02586_ _02589_ _02080_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_165_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ mod.u_cpu.rf_ram.memory\[461\]\[0\] _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09398__A1 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07165_ _01472_ _01473_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08445__I0 mod.u_cpu.rf_ram.memory\[396\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10252__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08070__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15133__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08373__A2 _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15283__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _01569_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09737_ _03916_ mod.u_cpu.rf_ram.memory\[554\]\[0\] _03920_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07505__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11094__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09668_ _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08619_ mod.u_cpu.rf_ram.memory\[152\]\[1\] mod.u_cpu.rf_ram.memory\[153\]\[1\] mod.u_cpu.rf_ram.memory\[154\]\[1\]
+ mod.u_cpu.rf_ram.memory\[155\]\[1\] _02066_ _02067_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12209__A1 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13406__B1 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09599_ _03812_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _04817_ _05227_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07240__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ _05182_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11432__A2 _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13300_ _06397_ _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13709__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10512_ _04468_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10491__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14280_ _00134_ net3 mod.u_cpu.rf_ram.memory\[547\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11492_ _04859_ _05125_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13231_ _06337_ _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10443_ _04400_ mod.u_cpu.rf_ram.memory\[451\]\[0\] _04420_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12232__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13162_ _06272_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _04218_ _04373_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11269__I _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12113_ _05550_ mod.u_cpu.rf_ram.memory\[68\]\[1\] _05556_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13093_ _05888_ _03878_ _06231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14500__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15626__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07247__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12044_ _05164_ _05433_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07167__A3 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12448__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13995_ mod.u_arbiter.i_wb_cpu_rdt\[11\] _06952_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14650__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12946_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12877_ _06073_ mod.u_cpu.rf_ram.memory\[246\]\[0\] _06074_ _06075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08527__B _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15006__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14616_ _00470_ net3 mod.u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11828_ _02430_ _05362_ _05363_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14070__B1 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15596_ _01367_ net3 mod.u_cpu.rf_ram.memory\[245\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08246__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14547_ _00401_ net3 mod.u_cpu.rf_ram.memory\[414\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12620__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11759_ _05265_ _05316_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14478_ _00332_ net3 mod.u_cpu.rf_ram.memory\[448\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15156__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13429_ _06515_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13420__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08970_ mod.u_cpu.cpu.bufreg2.i_cnt_done mod.u_cpu.cpu.immdec.imm31 _03274_ _03275_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07921_ _02120_ _02214_ _02219_ _02224_ _02228_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_111_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11734__I0 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10811__I _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07852_ _02156_ mod.u_cpu.rf_ram.memory\[196\]\[0\] _02159_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07392__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07783_ _01671_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09522_ _01850_ _03703_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09453_ _03395_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ _01518_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09384_ _03613_ _03622_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08335_ _02597_ _02637_ _02641_ _01651_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__I0 mod.u_cpu.rf_ram.memory\[218\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11414__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07713__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ _02472_ _02573_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13569__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07217_ _01524_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08197_ _02122_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07567__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14523__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07148_ _01450_ _01456_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10925__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10776__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10090_ _03821_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14673__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12800_ _06023_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15029__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13780_ _06494_ _06324_ _06380_ _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11102__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _03917_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12731_ _05919_ _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07857__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12850__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15450_ _01224_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12662_ _05932_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14401_ _00255_ net3 mod.u_cpu.rf_ram.memory\[487\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15179__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11613_ _05216_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10168__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12602__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15381_ _01156_ net3 mod.u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12593_ _05694_ _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14332_ _00186_ net3 mod.u_cpu.rf_ram.memory\[521\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08282__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11544_ _05170_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13479__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14263_ _00117_ net3 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _05123_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07477__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13214_ _06320_ _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _04409_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12905__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14194_ _07067_ _03389_ _03674_ _07093_ _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13145_ _06252_ _06263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10357_ _04362_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13076_ mod.u_cpu.rf_ram.memory\[105\]\[0\] _05971_ _06219_ _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10288_ _04315_ _04303_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12027_ _05501_ mod.u_cpu.rf_ram.memory\[58\]\[1\] _05499_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14130__I1 mod.u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13978_ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _06943_ _06946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09837__A2 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12929_ _06107_ mod.u_cpu.rf_ram.memory\[369\]\[0\] _06108_ _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11462__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10078__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15579_ _01350_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14546__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _02406_ _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _01820_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10207__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14696__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__A2 _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10383__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ mod.u_cpu.cpu.mem_bytecnt\[0\] mod.u_cpu.cpu.state.o_cnt\[2\] mod.u_cpu.cpu.mem_bytecnt\[1\]
+ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10541__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07904_ _01701_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ mod.u_cpu.rf_ram.memory\[575\]\[1\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12380__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ _01533_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08946__I _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07766_ _01890_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12132__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09828__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _03730_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07839__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15321__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ _01491_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08500__A2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09978__S _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ mod.u_cpu.cpu.state.init_done _01434_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _03605_ _03606_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12435__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ _02115_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15471__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09298_ _03547_ _03548_ _03549_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10071__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08249_ _02542_ _02544_ _02556_ _02491_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14188__I1 mod.u_cpu.rf_ram.memory\[244\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11260_ _04976_ mod.u_cpu.rf_ram.memory\[321\]\[1\] _04974_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12899__A1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10211_ _01625_ _04259_ _04260_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11191_ _04929_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11571__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _04209_ _04202_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08319__A2 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10073_ _04160_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14950_ _00804_ net3 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11323__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13901_ _03306_ _06881_ _06689_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14419__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14881_ _00735_ net3 mod.u_cpu.rf_ram.memory\[243\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10921__I1 mod.u_cpu.rf_ram.memory\[374\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13832_ _05790_ _03670_ _03679_ _06829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12123__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13763_ _06761_ _06763_ _06765_ _06766_ _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10975_ _04377_ _04780_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14569__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15502_ _01273_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12714_ _05967_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07925__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13694_ _06703_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15433_ _01208_ net3 mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12645_ _05918_ mod.u_cpu.rf_ram.memory\[147\]\[0\] _05921_ _05922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13623__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15364_ _01139_ net3 mod.u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12576_ _05875_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14315_ _00169_ net3 mod.u_cpu.rf_ram.memory\[530\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08524__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11527_ _05143_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15295_ _00055_ net4 mod.u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14246_ _00100_ net3 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11458_ _05096_ mod.u_cpu.rf_ram.memory\[28\]\[0\] _05111_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13000__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13937__I _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10409_ _04398_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14177_ _06181_ _03933_ _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11389_ mod.u_cpu.rf_ram.memory\[301\]\[1\] _05065_ _05063_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13128_ mod.u_arbiter.i_wb_cpu_rdt\[16\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _06253_ _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09507__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10361__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13059_ _04107_ _05589_ _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12362__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15344__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07620_ _01925_ mod.u_cpu.rf_ram.memory\[318\]\[0\] _01927_ _01783_ _01928_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07670__I _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07551_ mod.u_cpu.rf_ram.memory\[381\]\[0\] _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12288__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12814__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ _01740_ _01769_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08494__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15494__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _03483_ _03435_ _03484_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08246__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09152_ _03443_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08434__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08103_ _01778_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08797__A2 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09083_ net2 _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08034_ mod.u_cpu.rf_ram.memory\[88\]\[0\] mod.u_cpu.rf_ram.memory\[89\]\[0\] mod.u_cpu.rf_ram.memory\[90\]\[0\]
+ mod.u_cpu.rf_ram.memory\[91\]\[0\] _01673_ _01666_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08450__B _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _04099_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10271__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08936_ _02542_ _03235_ _03242_ _02518_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08867_ _02461_ mod.u_cpu.rf_ram.memory\[550\]\[1\] _03173_ _02578_ _03174_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08721__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07818_ _01568_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14711__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08798_ mod.u_cpu.rf_ram.memory\[64\]\[1\] mod.u_cpu.rf_ram.memory\[65\]\[1\] mod.u_cpu.rf_ram.memory\[66\]\[1\]
+ mod.u_cpu.rf_ram.memory\[67\]\[1\] _01561_ _01714_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _01487_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07288__A2 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10760_ _04196_ _03969_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14007__B1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09419_ _03439_ mod.u_scanchain_local.module_data_in\[66\] _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10691_ _04584_ mod.u_cpu.rf_ram.memory\[411\]\[0\] _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14861__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12430_ _05761_ mod.u_cpu.rf_ram.memory\[439\]\[1\] _05771_ _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13230__A1 _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08344__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13781__A2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12361_ _05535_ _05726_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15217__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14100_ _03885_ _07014_ _07033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11312_ _05013_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15080_ _00934_ net3 mod.u_cpu.rf_ram.memory\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12292_ _05443_ _05668_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14031_ _06984_ _06985_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11243_ _03967_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08096__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07755__I _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11395__I1 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11174_ _04882_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14241__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15367__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11277__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10125_ _04198_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11147__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10056_ _04148_ mod.u_cpu.rf_ram.memory\[50\]\[0\] _04149_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14933_ _00787_ net3 mod.u_cpu.rf_ram.memory\[226\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14391__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14864_ _00718_ net3 mod.u_cpu.rf_ram.memory\[250\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13815_ _06431_ _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14795_ _00649_ net3 mod.u_cpu.rf_ram.memory\[290\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10658__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13746_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _06658_ _06749_ _06751_ _06752_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10958_ _04756_ mod.u_cpu.rf_ram.memory\[368\]\[1\] _04767_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10283__A1 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13677_ _06451_ _06685_ _06687_ _06688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10889_ _04414_ _04722_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15416_ _01191_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08228__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12628_ _05910_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10035__A1 mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15347_ _01122_ net3 mod.u_cpu.rf_ram.memory\[379\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11083__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A2 _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12559_ _05855_ mod.u_cpu.rf_ram.memory\[161\]\[0\] _05863_ _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15278_ _00036_ net4 mod.u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14229_ _00083_ net3 mod.u_cpu.rf_ram.memory\[573\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11535__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12583__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08400__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10091__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09770_ _03936_ mod.u_cpu.rf_ram.memory\[551\]\[1\] _03943_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14734__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13827__A3 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08721_ _02591_ _03020_ _03027_ _01657_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11915__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09900__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08652_ _02136_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07603_ _01891_ _01901_ _01910_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08583_ _01722_ mod.u_cpu.rf_ram.memory\[286\]\[1\] _02889_ _02030_ _02890_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14884__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07534_ mod.u_cpu.rf_ram.memory\[320\]\[0\] mod.u_cpu.rf_ram.memory\[321\]\[0\] mod.u_cpu.rf_ram.memory\[322\]\[0\]
+ mod.u_cpu.rf_ram.memory\[323\]\[0\] _01841_ _01763_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07465_ _01750_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09204_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _03474_
+ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07396_ _01538_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09135_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11074__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10266__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _03361_ _03368_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14264__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ _02109_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13515__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07508__C _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09968_ _03919_ _04087_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08919_ mod.u_cpu.rf_ram.memory\[536\]\[1\] mod.u_cpu.rf_ram.memory\[537\]\[1\] mod.u_cpu.rf_ram.memory\[538\]\[1\]
+ mod.u_cpu.rf_ram.memory\[539\]\[1\] _02560_ _02495_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09899_ _04041_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11930_ _05436_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11861_ _05386_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13600_ _03713_ _04922_ _06621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _04668_ _04669_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08458__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14580_ _00434_ net3 mod.u_cpu.rf_ram.memory\[397\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11792_ mod.u_cpu.rf_ram.memory\[233\]\[0\] _04954_ _05339_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12254__A2 _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13531_ _06582_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _04574_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10377__S _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13462_ _03569_ _06531_ _06532_ _03574_ _06535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10674_ _04577_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15201_ _01054_ net3 mod.u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12413_ _05761_ mod.u_cpu.rf_ram.memory\[175\]\[1\] _05758_ _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14607__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13754__A2 _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13393_ _06442_ _06398_ _06486_ _06487_ _06488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11765__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15132_ _00985_ net3 mod.u_cpu.rf_ram.memory\[166\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12344_ _05715_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08630__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13506__A2 _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15063_ _00917_ net3 mod.u_cpu.rf_ram.memory\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10904__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12275_ _04984_ _05668_ _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14757__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11517__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14014_ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] _06966_ _06973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11226_ _04952_ mod.u_cpu.rf_ram.memory\[326\]\[1\] _04949_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11936__S _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11157_ _04360_ _04906_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10108_ _04043_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11088_ _04859_ _04848_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10879__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10039_ _04136_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14916_ _00770_ net3 mod.u_cpu.rf_ram.memory\[228\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08697__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13690__A1 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14847_ _00701_ net3 mod.u_cpu.rf_ram.memory\[264\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08449__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14778_ _00632_ net3 mod.u_cpu.rf_ram.memory\[298\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13729_ _06429_ _06732_ _06734_ _06735_ _06736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__11470__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07250_ _01511_ _01557_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14287__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15532__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07181_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07395__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13902__C1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _03985_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ _01486_ _03010_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14021__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09684_ _03809_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08688__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09115__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02097_ _02941_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15062__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08566_ _01791_ _02863_ _02872_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07517_ _01743_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08535__S1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08497_ _02672_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07448_ _01728_ mod.u_cpu.rf_ram.memory\[420\]\[0\] _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08860__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__A2 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13736__A2 _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _01686_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _03413_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10390_ _04365_ mod.u_cpu.rf_ram.memory\[460\]\[0\] _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09049_ _03352_ mod.u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12060_ _05523_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12172__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11011_ _04806_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__A2 mod.u_cpu.rf_ram.memory\[526\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12962_ _06138_ _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15405__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11913_ _05413_ mod.u_cpu.rf_ram.memory\[223\]\[0\] _05424_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14701_ _00555_ net3 mod.u_cpu.rf_ram.memory\[337\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12893_ _06073_ mod.u_cpu.rf_ram.memory\[98\]\[0\] _06084_ _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14632_ _00486_ net3 mod.u_cpu.rf_ram.memory\[371\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11844_ _05366_ mod.u_cpu.rf_ram.memory\[159\]\[0\] _05375_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14563_ _00417_ net3 mod.u_cpu.rf_ram.memory\[406\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13975__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15555__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11775_ _05106_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10726_ _04611_ _04610_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13514_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03388_ _03337_ _06568_ _06569_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14494_ _00348_ net3 mod.u_cpu.rf_ram.memory\[440\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13445_ _06524_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10657_ _04290_ _04437_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11738__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12786__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11589__I1 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13376_ _06130_ _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10588_ _04518_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15115_ _00968_ net3 mod.u_cpu.rf_ram.memory\[419\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12327_ _05667_ _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15046_ _00900_ net3 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12258_ _05656_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11209_ _04941_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12189_ _05609_ mod.u_cpu.rf_ram.memory\[203\]\[1\] _05607_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10713__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07590__A1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15085__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13663__A1 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_160 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12466__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12710__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_171 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08420_ mod.u_cpu.rf_ram.memory\[415\]\[1\] _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10229__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08351_ _02085_ mod.u_cpu.rf_ram.memory\[492\]\[1\] _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09095__A1 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ _01608_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08282_ _02560_ _02587_ _02588_ _02188_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08842__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14215__I0 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14922__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07233_ mod.u_cpu.rf_ram.memory\[456\]\[0\] mod.u_cpu.rf_ram.memory\[457\]\[0\] mod.u_cpu.rf_ram.memory\[458\]\[0\]
+ mod.u_cpu.rf_ram.memory\[459\]\[0\] _01540_ _01501_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13718__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__S _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12777__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _01462_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10401__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__A2 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12529__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14302__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15428__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07853__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09805_ _03856_ _03966_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ _02303_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07581__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09736_ _03902_ _03919_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13654__A1 _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10468__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09322__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14452__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09667_ _03864_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15578__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07333__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _01849_ _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09598_ _03802_ mod.u_cpu.rf_ram.memory\[56\]\[0\] _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13406__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12209__A2 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ mod.u_cpu.rf_ram.memory\[317\]\[1\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11968__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11560_ _05180_ mod.u_cpu.rf_ram.memory\[273\]\[0\] _05181_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08833__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10511_ _04467_ mod.u_cpu.rf_ram.memory\[441\]\[1\] _04465_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13709__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10640__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11491_ _05135_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12768__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13230_ _06137_ _06133_ _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10442_ _04277_ _04407_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__C _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13161_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _06268_ _06272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11440__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10373_ _04308_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ _05557_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13092_ _06204_ _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12043_ _05511_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11285__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12448__A2 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13994_ _06910_ _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12945_ _03498_ _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14945__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12876_ _05494_ _05263_ _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14615_ _00469_ net3 mod.u_cpu.rf_ram.memory\[380\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _05348_ _05362_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_187_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15595_ _01366_ net3 mod.u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14546_ _00400_ net3 mod.u_cpu.rf_ram.memory\[414\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11758_ _05187_ _05279_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12620__A2 _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10631__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ _04598_ mod.u_cpu.rf_ram.memory\[408\]\[0\] _04600_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14477_ _00331_ net3 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11689_ _05139_ _05255_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13428_ _03371_ _06511_ _06514_ _03492_ _06515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13420__I1 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08262__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13359_ _06454_ _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__A2 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14325__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07920_ _02225_ _02226_ _02227_ _01683_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15029_ _00883_ net3 mod.u_cpu.rf_ram.memory\[203\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13884__A1 _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12687__A2 _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07673__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12931__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07851_ _02157_ _02158_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14475__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07782_ _01661_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _03744_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07315__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09452_ mod.u_cpu.cpu.decode.opcode\[1\] _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12020__S _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08403_ _02687_ _02702_ _02709_ _02606_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10870__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09383_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] _03615_ _03621_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08334_ _02638_ mod.u_cpu.rf_ram.memory\[502\]\[1\] _02640_ _01615_ _02641_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15100__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ mod.u_cpu.rf_ram.memory\[541\]\[0\] _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07216_ _01523_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _02455_ _02499_ _02503_ _02467_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _01451_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15250__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14818__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08426__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14968__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09504__S _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09719_ _03877_ mod.u_cpu.rf_ram.memory\[556\]\[0\] _03906_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10991_ _04791_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11833__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12730_ _05977_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07857__A2 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09303__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12661_ _05918_ mod.u_cpu.rf_ram.memory\[144\]\[0\] _05931_ _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14400_ _00254_ net3 mod.u_cpu.rf_ram.memory\[487\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _05199_ mod.u_cpu.rf_ram.memory\[264\]\[0\] _05215_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12592_ _05885_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15380_ _01155_ net3 mod.u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08806__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12602__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14331_ _00185_ net3 mod.u_cpu.rf_ram.memory\[522\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11543_ _05162_ mod.u_cpu.rf_ram.memory\[276\]\[1\] _05168_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14348__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14262_ _00116_ net3 mod.u_cpu.rf_ram.memory\[556\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09606__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11474_ _05108_ mod.u_cpu.rf_ram.memory\[287\]\[1\] _05121_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13213_ _06118_ _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10425_ _04400_ mod.u_cpu.rf_ram.memory\[454\]\[0\] _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14193_ _07092_ _05803_ _07093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13144_ _06262_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10356_ _04348_ mod.u_cpu.rf_ram.memory\[465\]\[0\] _04361_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14498__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13075_ _03713_ _05640_ _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10287_ _03781_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13866__A1 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12913__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12026_ _05483_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07426__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13977_ _06944_ _06945_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12928_ _05742_ _04704_ _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15123__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10852__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12859_ mod.u_cpu.rf_ram_if.rtrig1 mod.u_cpu.rf_ram.rdata\[1\] _06061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09845__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15578_ _01349_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14529_ _00383_ net3 mod.u_cpu.rf_ram.memory\[423\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12574__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15273__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _01823_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09222__A1 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08025__A2 _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13157__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11918__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08720__C _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07903_ _01924_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09525__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08883_ _02456_ mod.u_cpu.rf_ram.memory\[572\]\[1\] _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11854__S _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07834_ _02110_ _02133_ _02140_ _02141_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ _02053_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11653__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12132__I1 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ mod.u_cpu.rf_ram.memory\[9\]\[0\] _03699_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10143__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07696_ _01722_ mod.u_cpu.rf_ram.memory\[286\]\[0\] _02003_ _01970_ _02004_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09435_ mod.u_cpu.cpu.immdec.imm11_7\[0\] mod.u_cpu.cpu.immdec.imm11_7\[1\] _03664_
+ _03665_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14034__A1 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09366_ _03605_ _03606_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15616__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12596__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08317_ mod.u_cpu.rf_ram.memory\[471\]\[1\] _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11643__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__A1 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09297_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03543_
+ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_21_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07578__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08248_ _02545_ _02549_ _02554_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14640__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08179_ _02010_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08647__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09793__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12899__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10210_ _04186_ _04259_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11190_ _04916_ mod.u_cpu.rf_ram.memory\[332\]\[1\] _04927_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08567__A3 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13148__I0 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10141_ _03872_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14790__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10072_ _04148_ mod.u_cpu.rf_ram.memory\[506\]\[0\] _04159_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12520__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13900_ _06677_ _06885_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14880_ _00734_ net3 mod.u_cpu.rf_ram.memory\[243\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13831_ _06135_ _06826_ _06828_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15146__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10134__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13762_ _03298_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _06421_ _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10974_ _04227_ _04779_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15501_ _01272_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12713_ _05966_ mod.u_cpu.rf_ram.memory\[7\]\[1\] _05964_ _05967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10834__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13693_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _06658_ _06700_ _06702_ _06703_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15432_ _01207_ net3 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15296__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12644_ _05732_ _05920_ _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08805__C _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15363_ _01138_ net3 mod.u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12575_ _05874_ mod.u_cpu.rf_ram.memory\[15\]\[1\] _05871_ _05875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08093__B _02400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11004__S _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14314_ _00168_ net3 mod.u_cpu.rf_ram.memory\[530\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11526_ _05158_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15294_ _00054_ net4 mod.u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14245_ _00099_ net3 mod.u_cpu.rf_ram.memory\[565\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11457_ _05110_ _03782_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08638__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13000__A2 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10408_ mod.u_cpu.rf_ram.memory\[457\]\[0\] _04396_ _04397_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14176_ _07082_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11388_ _04531_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13139__I0 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _04350_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13127_ _06252_ _06253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A2 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13058_ _06208_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12009_ _05484_ mod.u_cpu.rf_ram.memory\[575\]\[1\] _05486_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12997__C _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08191__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12569__I _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _01758_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14513__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15639__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12814__A2 _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ _01770_ _01772_ _01786_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09220_ _03410_ mod.u_scanchain_local.module_data_in\[36\] _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07900__B _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09151_ mod.u_arbiter.i_wb_cpu_rdt\[6\] _03441_ _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14663__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10428__I1 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08246__A2 mod.u_cpu.rf_ram.memory\[526\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08102_ _01646_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09082_ net1 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11250__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _01696_ _02340_ _02321_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15019__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07757__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12750__A1 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _04091_ mod.u_cpu.rf_ram.memory\[520\]\[1\] _04097_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09118__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08935_ _02545_ _03238_ _03241_ _02555_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15169__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08866_ _02462_ _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12479__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07817_ _01672_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_57_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08797_ _02348_ _03103_ _01618_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09989__S _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07748_ _02053_ _02055_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11864__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14007__A1 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07679_ _01938_ mod.u_cpu.rf_ram.memory\[278\]\[0\] _01986_ _01952_ _01987_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08906__B _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09788__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] _03615_ _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09809__I0 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10690_ _04457_ _04575_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08625__C _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09349_ _03588_ _03590_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13230__A2 _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12360_ _05725_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__I1 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11311_ _05007_ mod.u_cpu.rf_ram.memory\[313\]\[0\] _05012_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12291_ _05604_ _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14030_ mod.u_arbiter.i_wb_cpu_rdt\[20\] _06976_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11242_ _04964_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08096__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11558__I _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11173_ _04917_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10124_ _04193_ mod.u_cpu.rf_ram.memory\[4\]\[0\] _04197_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10055_ _04013_ _03859_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14932_ _00786_ net3 mod.u_cpu.rf_ram.memory\[226\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14536__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08173__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14863_ _00717_ net3 mod.u_cpu.rf_ram.memory\[257\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13814_ _06810_ _06813_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14794_ _00648_ net3 mod.u_cpu.rf_ram.memory\[290\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07359__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13745_ _06656_ _06750_ _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14686__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10957_ _04768_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09698__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10283__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13676_ _06437_ _06448_ _06686_ _06372_ _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10888_ _04389_ _04108_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_31_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15415_ _01190_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13757__B1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12627_ _05904_ mod.u_cpu.rf_ram.memory\[150\]\[0\] _05909_ _05910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08079__I2 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13221__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08107__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15346_ _01121_ net3 mod.u_cpu.rf_ram.memory\[389\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12558_ _05657_ _05757_ _05863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11509_ _05147_ mod.u_cpu.rf_ram.memory\[282\]\[1\] _05145_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15277_ _00035_ net4 mod.u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12489_ _05807_ mod.u_cpu.rf_ram.memory\[171\]\[1\] _05817_ _05819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14228_ _00082_ net3 mod.u_cpu.rf_ram.memory\[573\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12032__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12732__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11535__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15311__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14159_ _06153_ _03270_ _01407_ _07070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13288__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09382__B _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08720_ _01698_ _03023_ _03026_ _02347_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15461__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08651_ mod.u_cpu.rf_ram.memory\[167\]\[1\] _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07911__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07602_ _01872_ _01902_ _01909_ _01657_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08582_ _02027_ _02888_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07533_ _01710_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11846__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10748__S _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__A2 mod.u_cpu.rf_ram.memory\[374\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11931__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07464_ mod.u_cpu.rf_ram.memory\[424\]\[0\] mod.u_cpu.rf_ram.memory\[425\]\[0\] mod.u_cpu.rf_ram.memory\[426\]\[0\]
+ mod.u_cpu.rf_ram.memory\[427\]\[0\] _01753_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09203_ _03414_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07395_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _03428_ _03387_ _03421_ _03429_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08017__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14409__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07978__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _03300_ _03367_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12762__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08016_ mod.u_cpu.rf_ram.memory\[112\]\[0\] mod.u_cpu.rf_ram.memory\[113\]\[0\] mod.u_cpu.rf_ram.memory\[114\]\[0\]
+ mod.u_cpu.rf_ram.memory\[115\]\[0\] _01664_ _02323_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11378__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08180__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14559__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09967_ _03995_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08918_ _03215_ _03224_ _01447_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09898_ _04036_ mod.u_cpu.rf_ram.memory\[534\]\[1\] _04039_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _03001_ _03155_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _03726_ _04378_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13987__B1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11837__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ _04569_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11791_ _05078_ _05320_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11841__I _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13530_ _06581_ mod.u_cpu.rf_ram.memory\[129\]\[1\] _06579_ _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10742_ _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10673_ _04557_ mod.u_cpu.rf_ram.memory\[414\]\[0\] _04576_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13461_ _06534_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15200_ _01053_ net3 mod.u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12412_ _05710_ _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13392_ _06470_ _06397_ _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15131_ _00984_ net3 mod.u_cpu.rf_ram.memory\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15334__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11765__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12343_ _05713_ mod.u_cpu.rf_ram.memory\[182\]\[0\] _05714_ _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12014__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12274_ _05667_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15062_ _00916_ net3 mod.u_cpu.rf_ram.memory\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11517__A2 _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14013_ _06969_ _06972_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ _04951_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15484__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11156_ _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10107_ _04184_ _04173_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11087_ _03780_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10038_ _04135_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14915_ _00769_ net3 mod.u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08697__A2 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13690__A2 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14846_ _00700_ net3 mod.u_cpu.rf_ram.memory\[264\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__A2 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14777_ _00631_ net3 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11989_ _02485_ _05475_ _05476_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11751__I _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13728_ _06494_ _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07752__S0 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10367__I _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13659_ _06371_ _06670_ _06671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11205__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07180_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15329_ mod.u_cpu.cpu.o_wen1 net3 mod.u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14701__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13902__B1 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__C2 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09891__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09821_ _03984_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14851__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _03931_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08137__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09334__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08703_ _02997_ _02999_ _01891_ _03009_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09683_ _03739_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07344__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15207__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ mod.u_cpu.rf_ram.memory\[188\]\[1\] mod.u_cpu.rf_ram.memory\[189\]\[1\] mod.u_cpu.rf_ram.memory\[190\]\[1\]
+ mod.u_cpu.rf_ram.memory\[191\]\[1\] _02092_ _02098_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07360__A2 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11819__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ _01956_ _02864_ _02871_ _01989_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15280__D _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ mod.u_cpu.rf_ram.memory\[348\]\[0\] mod.u_cpu.rf_ram.memory\[349\]\[0\] mod.u_cpu.rf_ram.memory\[350\]\[0\]
+ mod.u_cpu.rf_ram.memory\[351\]\[0\] _01823_ _01821_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12492__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08496_ mod.u_cpu.rf_ram.memory\[335\]\[1\] _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14231__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07447_ _01753_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10277__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15357__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12693__S _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ _01527_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09117_ _03279_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14381__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09048_ _03250_ _03348_ _03351_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10558__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _04803_ mod.u_cpu.rf_ram.memory\[360\]\[0\] _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12172__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10740__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08210__I _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12961_ _06137_ _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08518__I3 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14700_ _00554_ net3 mod.u_cpu.rf_ram.memory\[337\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11912_ _04845_ _05423_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12892_ _03974_ _06048_ _06084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14631_ _00485_ net3 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11843_ _04845_ _05374_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14562_ _00416_ net3 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11774_ _05327_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13513_ _05791_ _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10725_ _04541_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14493_ _00347_ net3 mod.u_cpu.rf_ram.memory\[441\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14724__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13444_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _06519_ _06520_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10656_ _04564_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11738__A2 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13498__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12786__I1 mod.u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13375_ _06470_ _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10587_ _04514_ mod.u_cpu.rf_ram.memory\[428\]\[1\] _04516_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12108__S _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08603__A2 _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09800__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15114_ _00967_ net3 mod.u_cpu.rf_ram.memory\[419\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12326_ _05702_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14874__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15045_ _00899_ net3 mod.u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12257_ _05635_ mod.u_cpu.rf_ram.memory\[194\]\[1\] _05654_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11208_ _04936_ mod.u_cpu.rf_ram.memory\[32\]\[1\] _04939_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12188_ _05549_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11139_ _04883_ mod.u_cpu.rf_ram.memory\[340\]\[0\] _04894_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13663__A2 _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_150 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_161 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_172 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14254__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14829_ _00683_ net3 mod.u_cpu.rf_ram.memory\[273\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09619__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11481__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10229__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ mod.u_cpu.rf_ram.memory\[493\]\[1\] _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11426__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ mod.u_cpu.rf_ram.memory\[509\]\[0\] _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10097__I _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08281_ _02198_ mod.u_cpu.rf_ram.memory\[460\]\[1\] _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08842__A2 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13179__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07232_ _01539_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ mod.u_cpu.cpu.immdec.imm24_20\[2\] _01467_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12018__S _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08445__I2 mod.u_cpu.rf_ram.memory\[398\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11857__S _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10761__S _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _03972_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07996_ mod.u_cpu.rf_ram.memory\[111\]\[0\] _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09735_ _03918_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10468__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ _03768_ _03848_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08617_ mod.u_cpu.rf_ram.memory\[136\]\[1\] mod.u_cpu.rf_ram.memory\[137\]\[1\] mod.u_cpu.rf_ram.memory\[138\]\[1\]
+ mod.u_cpu.rf_ram.memory\[139\]\[1\] _02022_ _02043_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _03805_ _03810_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ mod.u_cpu.rf_ram.memory\[312\]\[1\] mod.u_cpu.rf_ram.memory\[313\]\[1\] mod.u_cpu.rf_ram.memory\[314\]\[1\]
+ mod.u_cpu.rf_ram.memory\[315\]\[1\] _01802_ _01932_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14747__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11968__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08479_ _01997_ _02782_ _02785_ _02096_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10510_ _04429_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10640__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11490_ _05128_ mod.u_cpu.rf_ram.memory\[285\]\[1\] _05131_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _04419_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14897__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13160_ _06271_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10372_ _04372_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11440__I1 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12111_ _05539_ mod.u_cpu.rf_ram.memory\[68\]\[0\] _05556_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13091_ _06229_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13342__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ _05501_ mod.u_cpu.rf_ram.memory\[60\]\[1\] _05509_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14142__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14277__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] _06954_ _06957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09849__A1 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15522__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12944_ _06118_ _06120_ _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08521__A1 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08808__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12875_ _06072_ _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14614_ _00468_ net3 mod.u_cpu.rf_ram.memory\[380\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _04294_ _03942_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15594_ _01365_ net3 mod.u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14070__A2 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14545_ _00399_ net3 mod.u_cpu.rf_ram.memory\[415\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11757_ _05315_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10708_ _04168_ _04599_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14476_ _00330_ net3 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11688_ _05221_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08543__C _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10645__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13427_ _06513_ _06514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10639_ _04553_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13358_ _06395_ _06380_ _06131_ _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10395__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _05679_ mod.u_cpu.rf_ram.memory\[185\]\[0\] _05690_ _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13289_ _03501_ _03428_ _06386_ _06387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__15052__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09147__S _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15028_ _00882_ net3 mod.u_cpu.rf_ram.memory\[203\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10147__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11476__I _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13884__A2 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08060__I0 mod.u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ mod.u_cpu.rf_ram.memory\[197\]\[0\] _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08760__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14133__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07781_ _01818_ _02082_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09520_ _03741_ _03743_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ _03678_ _03294_ _03677_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08402_ _02654_ _02705_ _02708_ _01979_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12100__I _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10870__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09382_ _03564_ _03617_ _03620_ _03417_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_178_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08333_ _02197_ _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ mod.u_cpu.rf_ram.memory\[536\]\[0\] mod.u_cpu.rf_ram.memory\[537\]\[0\] mod.u_cpu.rf_ram.memory\[538\]\[0\]
+ mod.u_cpu.rf_ram.memory\[539\]\[0\] _02450_ _02451_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10555__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07215_ _01497_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08195_ _02461_ mod.u_cpu.rf_ram.memory\[574\]\[0\] _02502_ _02465_ _02503_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08579__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07146_ _01452_ _01454_ _01448_ _01425_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07864__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08426__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15545__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10933__I0 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07979_ mod.u_cpu.rf_ram.memory\[103\]\[0\] _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09718_ _03902_ _03905_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__B _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _04772_ mod.u_cpu.rf_ram.memory\[363\]\[1\] _04789_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08503__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _03850_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12438__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12660_ _05300_ _05920_ _05931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _04804_ _05214_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12945__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12063__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12591_ _05874_ mod.u_cpu.rf_ram.memory\[156\]\[1\] _05883_ _05885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08806__A2 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14330_ _00184_ net3 mod.u_cpu.rf_ram.memory\[522\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11810__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11542_ _05169_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14261_ _00115_ net3 mod.u_cpu.rf_ram.memory\[557\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07490__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11473_ _02002_ _05121_ _05122_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15075__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08114__S0 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13212_ _06318_ _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10424_ _04262_ _04407_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14192_ mod.u_cpu.rf_ram_if.rgnt _07092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13143_ mod.u_arbiter.i_wb_cpu_rdt\[23\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _06258_ _06262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10355_ _04360_ _04353_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A2 _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10286_ _04314_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13074_ _06218_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13866__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12025_ _05500_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12913__I1 mod.u_cpu.rf_ram.memory\[399\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11877__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14912__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11629__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12677__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13976_ mod.u_arbiter.i_wb_cpu_rdt\[6\] _06938_ _06928_ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _06945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12927_ _06072_ _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15646_ _01417_ net3 mod.u_cpu.rf_ram.memory\[249\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12858_ mod.u_cpu.rf_ram_if.rdata1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10852__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11809_ _05351_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15577_ _01348_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12789_ _06010_ mod.u_cpu.rf_ram.memory\[130\]\[0\] _06015_ _06016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09845__I1 mod.u_cpu.rf_ram.memory\[542\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15418__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14528_ _00382_ net3 mod.u_cpu.rf_ram.memory\[423\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13929__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07481__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14459_ _00313_ net3 mod.u_cpu.rf_ram.memory\[458\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14442__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15568__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07684__I _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08951_ _03252_ _03253_ _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13857__A2 _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07902_ mod.u_cpu.rf_ram.memory\[211\]\[0\] _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11868__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08882_ _02457_ _03188_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10915__I0 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14592__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07833_ _01716_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15553__D _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07764_ mod.u_cpu.rf_ram.memory\[140\]\[0\] mod.u_cpu.rf_ram.memory\[141\]\[0\] mod.u_cpu.rf_ram.memory\[142\]\[0\]
+ mod.u_cpu.rf_ram.memory\[143\]\[0\] _02070_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09503_ _03714_ _03728_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11340__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07695_ _01967_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ mod.u_cpu.cpu.immdec.imm11_7\[4\] _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14034__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12045__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10486__S _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09365_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03595_
+ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_178_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15098__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ _02566_ mod.u_cpu.rf_ram.memory\[468\]\[1\] _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12596__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09296_ _03541_ _03543_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12840__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _02308_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ _02484_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08647__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07129_ _01425_ _01432_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_137_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__I2 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10140_ _04208_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14935__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13848__A2 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10071_ _03797_ _04143_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12005__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12520__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10531__A1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13830_ mod.u_cpu.cpu.immdec.imm30_25\[4\] _06773_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[5\]
+ _06827_ _06339_ _06828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13761_ _03686_ _06764_ _06765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10973_ _03663_ _04223_ _03724_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10134__I1 mod.u_cpu.rf_ram.memory\[498\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15500_ _01271_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14315__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12712_ _05937_ _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13692_ _06656_ _06701_ _06702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14025__A2 _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15431_ _01206_ net3 mod.u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _05919_ _05920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07769__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13784__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15362_ _01137_ net3 mod.u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12574_ _05873_ _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12831__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11634__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14465__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08093__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14313_ _00167_ net3 mod.u_cpu.rf_ram.memory\[531\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10195__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11525_ _05147_ mod.u_cpu.rf_ram.memory\[27\]\[1\] _05156_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15293_ _00053_ net4 mod.u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14244_ _00098_ net3 mod.u_cpu.rf_ram.memory\[565\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11456_ _04195_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08638__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08821__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _03714_ _04380_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14175_ _07081_ mod.u_cpu.rf_ram.memory\[88\]\[1\] _07079_ _07082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11387_ _01964_ _05063_ _05064_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13139__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13126_ _05785_ _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10338_ _04348_ mod.u_cpu.rf_ram.memory\[468\]\[0\] _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13839__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _06199_ mod.u_cpu.rf_ram.memory\[82\]\[1\] _06206_ _06208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10269_ _04132_ _04300_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08715__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _02501_ _05486_ _05489_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08810__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12275__A1 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13959_ _06920_ _05794_ _06930_ _06931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15240__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15629_ _01400_ net3 mod.u_cpu.rf_ram.memory\[279\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14808__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09818__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09150_ _03417_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10589__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08101_ _02316_ mod.u_cpu.rf_ram.memory\[20\]\[0\] _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15390__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09081_ _03301_ _03378_ _03382_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11250__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09894__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14958__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08032_ mod.u_cpu.rf_ram.memory\[84\]\[0\] mod.u_cpu.rf_ram.memory\[85\]\[0\] mod.u_cpu.rf_ram.memory\[86\]\[0\]
+ mod.u_cpu.rf_ram.memory\[87\]\[0\] _01857_ _02054_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_163_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08629__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08731__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07206__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10061__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A2 _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09983_ _04098_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ _02550_ mod.u_cpu.rf_ram.memory\[534\]\[1\] _03240_ _02515_ _03241_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08865_ mod.u_cpu.rf_ram.memory\[551\]\[1\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14338__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07816_ _01687_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08796_ mod.u_cpu.rf_ram.memory\[72\]\[1\] mod.u_cpu.rf_ram.memory\[73\]\[1\] mod.u_cpu.rf_ram.memory\[74\]\[1\]
+ mod.u_cpu.rf_ram.memory\[75\]\[1\] _02211_ _02386_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07747_ mod.u_cpu.rf_ram.memory\[132\]\[0\] mod.u_cpu.rf_ram.memory\[133\]\[0\] mod.u_cpu.rf_ram.memory\[134\]\[0\]
+ mod.u_cpu.rf_ram.memory\[135\]\[0\] _01893_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09131__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07678_ _01949_ _01985_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11864__I1 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14488__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ _03614_ _03649_ _03650_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_125_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07693__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ _03568_ _03591_ _03592_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _03533_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_148_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _04873_ _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12290_ _05678_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10743__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11241_ _04952_ mod.u_cpu.rf_ram.memory\[324\]\[1\] _04962_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07748__A2 _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11172_ _04916_ mod.u_cpu.rf_ram.memory\[335\]\[1\] _04914_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15113__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10123_ _04196_ _03961_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10054_ _04147_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14931_ _00785_ net3 mod.u_cpu.rf_ram.memory\[227\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11552__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14862_ _00716_ net3 mod.u_cpu.rf_ram.memory\[257\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15263__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13813_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _06773_ _06807_ _06811_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[3\]
+ _06813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14793_ _00647_ net3 mod.u_cpu.rf_ram.memory\[291\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09122__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07359__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13744_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _06139_ _06338_ _06741_ _06750_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10956_ _04753_ mod.u_cpu.rf_ram.memory\[368\]\[0\] _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13057__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13675_ _06431_ _06490_ _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10887_ _04721_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15414_ _01189_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13757__A1 _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13757__B2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12626_ _05494_ _05900_ _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12804__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__A2 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__I3 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15345_ _01120_ net3 mod.u_cpu.rf_ram.memory\[389\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12557_ _05862_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10035__A3 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11508_ _05107_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15276_ _00034_ net4 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12980__A2 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12488_ _05818_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11749__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14227_ _00081_ net3 mod.u_cpu.rf_ram.memory\[574\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14182__A1 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12032__I1 mod.u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11439_ _05098_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12732__A2 _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14158_ _07069_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13109_ _06241_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14089_ _03774_ _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15606__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11543__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11484__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ _02129_ mod.u_cpu.rf_ram.memory\[164\]\[1\] _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _01874_ _01905_ _01908_ _01884_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08581_ mod.u_cpu.rf_ram.memory\[287\]\[1\] _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14630__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ mod.u_cpu.rf_ram.memory\[340\]\[0\] mod.u_cpu.rf_ram.memory\[341\]\[0\] mod.u_cpu.rf_ram.memory\[342\]\[0\]
+ mod.u_cpu.rf_ram.memory\[343\]\[0\] _01826_ _01828_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__I1 mod.u_cpu.rf_ram.memory\[233\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ _01569_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07675__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11471__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13204__I _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09202_ _03473_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14780__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07394_ _01701_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07202__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _03363_ _03416_ _03426_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07427__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _03362_ _03363_ _03355_ _03364_ _03366_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__12971__A2 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15136__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08015_ _01665_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09129__I _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10585__I1 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09966_ _04086_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15286__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07872__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _02471_ _03216_ _03223_ _02491_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09897_ _04040_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11394__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08848_ mod.u_cpu.rf_ram.memory\[37\]\[1\] _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13287__I0 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08779_ _01688_ _03078_ _03085_ _02291_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09799__I _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13987__A1 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _03941_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _05338_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11837__I1 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13039__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ _04620_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13739__A1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13460_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _06531_ _06532_ _03569_ _06534_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10672_ _04299_ _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12411_ _02117_ _05758_ _05760_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07418__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13391_ _06435_ _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15130_ _00983_ net3 mod.u_cpu.rf_ram.memory\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07969__A2 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12342_ _05494_ _05703_ _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08091__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10973__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11569__I _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14164__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08371__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15061_ _00915_ net3 mod.u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07268__B _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12273_ _05666_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14503__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14012_ _03458_ _06964_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _06972_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15629__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11224_ _04795_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11155_ _04846_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07782__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10106_ _03835_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11086_ _04858_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14653__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11525__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10037_ _03992_ _04132_ _04134_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_14914_ _00768_ net3 mod.u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11150__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14845_ _00699_ net3 mod.u_cpu.rf_ram.memory\[265\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15009__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13978__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14776_ _00630_ net3 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11988_ _05448_ _05475_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13727_ _06417_ _06733_ _06321_ _06486_ _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07657__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _04719_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12650__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07752__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13658_ _06667_ _06669_ _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15159__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12609_ _05887_ mod.u_cpu.rf_ram.memory\[153\]\[0\] _05897_ _05898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12863__I _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11205__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12402__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13589_ _06615_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10264__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15328_ _01105_ net3 mod.u_cpu.rf_ram.memory\[409\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13895__S _06882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14155__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15259_ _00015_ net4 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__I0 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13902__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__B2 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _03870_ _03966_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07906__B _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _03711_ _03779_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08137__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09334__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08702_ _02665_ _03000_ _03008_ _02852_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09682_ _03876_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _02090_ _02939_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07440__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13643__B _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08564_ _01961_ _02867_ _02870_ _01972_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09637__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08456__C _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07515_ _01506_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08495_ _02041_ mod.u_cpu.rf_ram.memory\[332\]\[1\] _02801_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07446_ mod.u_cpu.rf_ram.memory\[421\]\[0\] _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07377_ _01680_ _01684_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14526__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09116_ _03414_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12944__A2 _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08073__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10955__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _03349_ _03296_ _03350_ _03250_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14676__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09949_ _04071_ mod.u_cpu.rf_ram.memory\[526\]\[1\] _04074_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09325__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12960_ mod.u_arbiter.i_wb_cpu_ack _03399_ _06136_ _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12180__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11911_ _05422_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _06083_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14630_ _00484_ net3 mod.u_cpu.rf_ram.memory\[372\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11842_ _05373_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14561_ _00415_ net3 mod.u_cpu.rf_ram.memory\[407\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07639__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11773_ _05311_ mod.u_cpu.rf_ram.memory\[236\]\[0\] _05326_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15301__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08300__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13512_ _06567_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10724_ _04184_ _04574_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14492_ _00346_ net3 mod.u_cpu.rf_ram.memory\[441\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13188__A2 _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13443_ _06523_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10655_ _04560_ mod.u_cpu.rf_ram.memory\[417\]\[1\] _04562_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07777__I _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15451__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13374_ _06374_ _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10586_ _04517_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09800__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15113_ _00002_ net3 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12325_ _05692_ mod.u_cpu.rf_ram.memory\[179\]\[1\] _05700_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07811__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15044_ _00898_ net3 mod.u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12256_ _05655_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08367__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11207_ _04940_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12187_ _05608_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _04749_ _04887_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09316__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ _04846_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_140 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_151 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_162 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10579__S _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_173 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07878__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14828_ _00682_ net3 mod.u_cpu.rf_ram.memory\[273\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14759_ _00613_ net3 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07300_ _01510_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14549__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08280_ mod.u_cpu.rf_ram.memory\[461\]\[1\] _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12593__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07162_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11985__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14699__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08445__I3 mod.u_cpu.rf_ram.memory\[399\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13351__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11362__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09803_ _03964_ mod.u_cpu.rf_ram.memory\[547\]\[1\] _03970_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07995_ _01862_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09734_ _03917_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09665_ _03863_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07869__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15324__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _02916_ _02918_ _02920_ _02922_ _01658_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09596_ _03809_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12614__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08547_ _02841_ _02843_ _01891_ _02853_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08294__A1 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15474__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _01875_ mod.u_cpu.rf_ram.memory\[366\]\[1\] _02784_ _02030_ _02785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07429_ _01486_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12217__I1 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10440_ _04410_ mod.u_cpu.rf_ram.memory\[452\]\[1\] _04417_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08046__A1 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08597__A2 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ _04363_ mod.u_cpu.rf_ram.memory\[463\]\[1\] _04370_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10952__S _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12110_ _05367_ _05543_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13090_ _06217_ mod.u_cpu.rf_ram.memory\[103\]\[1\] _06227_ _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13878__B1 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13342__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12041_ _05510_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14142__I1 mod.u_cpu.rf_ram.memory\[289\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13992_ _06955_ _06956_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09849__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12943_ _05784_ _03458_ _06119_ _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _03923_ _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11825_ _05361_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14613_ _00467_ net3 mod.u_cpu.rf_ram.memory\[381\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15593_ _01364_ net3 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13802__B1 _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14544_ _00398_ net3 mod.u_cpu.rf_ram.memory\[415\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11756_ _05304_ mod.u_cpu.rf_ram.memory\[238\]\[1\] _05313_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13730__C _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10092__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ _04574_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14475_ _00329_ net3 mod.u_cpu.rf_ram.memory\[450\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14841__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11687_ _05267_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08037__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13426_ _06512_ _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10638_ _04537_ mod.u_cpu.rf_ram.memory\[420\]\[1\] _04551_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13030__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07300__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13357_ _06449_ _06451_ _06452_ _06453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10569_ _04505_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10395__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14991__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12308_ _04873_ _05686_ _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ _06377_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _06386_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15027_ _00881_ net3 mod.u_cpu.rf_ram.memory\[204\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12239_ mod.u_cpu.rf_ram.memory\[109\]\[1\] _05617_ _05641_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15347__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ _02083_ _02087_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12144__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 io_in[8] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xtiny_user_project_90 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12695__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12844__A1 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09450_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r
+ _03265_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14371__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15497__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08401_ _02692_ mod.u_cpu.rf_ram.memory\[438\]\[1\] _02707_ _01981_ _02708_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09381_ _03618_ _03619_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13413__S _06503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10458__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08332_ mod.u_cpu.rf_ram.memory\[503\]\[1\] _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08276__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ _02523_ _02562_ _02570_ _02469_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07214_ _01520_ _01521_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08028__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08194_ _02500_ _02501_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07210__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09776__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07145_ mod.u_cpu.cpu.decode.op26 _01453_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A2 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10933__I1 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08751__A2 _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13088__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ _02129_ mod.u_cpu.rf_ram.memory\[100\]\[0\] _02285_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07880__I _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14714__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12135__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09717_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07813__C _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09648_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14864__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09579_ _03745_ _03786_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10449__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11610_ _05119_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08267__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12063__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12590_ _05884_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__C _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11541_ _05159_ mod.u_cpu.rf_ram.memory\[276\]\[0\] _05168_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11810__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14260_ _00114_ net3 mod.u_cpu.rf_ram.memory\[557\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13012__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _05022_ _05121_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07490__A2 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07120__I mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13211_ _06317_ _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08114__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ _04308_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12961__I _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14191_ _07091_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13142_ _06261_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10354_ _03865_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14244__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09519__A1 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13073_ _06217_ mod.u_cpu.rf_ram.memory\[81\]\[1\] _06215_ _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10285_ _04313_ mod.u_cpu.rf_ram.memory\[477\]\[1\] _04310_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12024_ _05498_ mod.u_cpu.rf_ram.memory\[58\]\[0\] _05499_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14394__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13725__C _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07790__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12126__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12826__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11629__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13975_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] _06943_ _06944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07723__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11018__S _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10688__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12926_ _06106_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15645_ _01416_ net3 mod.u_cpu.rf_ram.memory\[249\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12857_ _01464_ mod.u_cpu.rf_ram.regzero _06059_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11808_ _05350_ mod.u_cpu.rf_ram.memory\[231\]\[1\] _05347_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15576_ _01347_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12788_ _03974_ _06011_ _06015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10065__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14527_ _00381_ net3 mod.u_cpu.rf_ram.memory\[424\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11739_ _05289_ mod.u_cpu.rf_ram.memory\[240\]\[0\] _05302_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13003__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14458_ _00312_ net3 mod.u_cpu.rf_ram.memory\[458\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07481__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13409_ _06501_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14389_ _00243_ net3 mod.u_cpu.rf_ram.memory\[493\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10368__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10612__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11487__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08950_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12365__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14737__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07901_ _02091_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08881_ mod.u_cpu.rf_ram.memory\[573\]\[1\] _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11868__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07832_ _02135_ mod.u_cpu.rf_ram.memory\[166\]\[0\] _02138_ _02139_ _02140_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12117__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08729__C _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07763_ _01746_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14887__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09502_ _03723_ _03727_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08497__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07694_ mod.u_cpu.rf_ram.memory\[287\]\[0\] _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11340__I1 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09433_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13143__S _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12045__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _02225_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09295_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08246_ _02550_ mod.u_cpu.rf_ram.memory\[526\]\[0\] _02553_ _02515_ _02554_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14267__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15512__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__I _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08177_ mod.u_cpu.rf_ram.memory\[559\]\[0\] _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07128_ _01433_ _01434_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08421__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11397__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__I3 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10070_ _04158_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13826__B _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12108__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__I2 mod.u_cpu.rf_ram.memory\[498\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13760_ mod.u_cpu.cpu.immdec.imm31 _03274_ _06764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_29_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10972_ _04778_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08032__S0 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08488__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12711_ _05965_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13691_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _06678_ _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15042__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15430_ _01205_ net3 mod.u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12642_ _05372_ _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__A1 _06325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__B2 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15361_ _01136_ net3 mod.u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12573_ _05709_ _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14312_ _00166_ net3 mod.u_cpu.rf_ram.memory\[531\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11524_ _05157_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15292_ _00051_ net4 mod.u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08660__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15192__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14243_ _00097_ net3 mod.u_cpu.rf_ram.memory\[566\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11455_ _05109_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07785__I _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10406_ _03924_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08412__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14174_ _03928_ _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11386_ _04817_ _05063_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13125_ _06251_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10337_ _04189_ _04327_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11100__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _06207_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10268_ _03721_ _04133_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_12007_ _05488_ _05486_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10199_ _04249_ mod.u_cpu.rf_ram.memory\[48\]\[0\] _04252_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07923__B1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13958_ _03441_ _05793_ _06930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12909_ _06095_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13889_ _06868_ _06836_ _06872_ _06880_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15628_ _01399_ net3 mod.u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13224__A1 _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09240__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15535__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10386__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15559_ _01330_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08100_ _02406_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11786__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09080_ _03378_ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08031_ _02090_ _02338_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09396__B _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07206__A2 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08403__A1 _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08254__I1 mod.u_cpu.rf_ram.memory\[529\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10061__I1 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04096_ mod.u_cpu.rf_ram.memory\[520\]\[0\] _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _02551_ _03239_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11010__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08864_ _02456_ mod.u_cpu.rf_ram.memory\[548\]\[1\] _03170_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07815_ _01670_ _02108_ _02121_ _02122_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _02465_ _03098_ _03101_ _02660_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ _01569_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15065__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12510__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09131__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07677_ mod.u_cpu.rf_ram.memory\[279\]\[0\] _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11680__I _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09416_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03635_
+ _03632_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10029__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09150__I _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _03436_ mod.u_scanchain_local.module_data_in\[55\] _03402_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13766__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09278_ _03525_ _03532_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14902__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _01747_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13518__A2 _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11240_ _04963_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11171_ _04879_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12016__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12329__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10122_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10053_ _03738_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09745__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14930_ _00784_ net3 mod.u_cpu.rf_ram.memory\[227\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15408__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__C _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14861_ _00715_ net3 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13829__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13812_ _06482_ _06772_ _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14792_ _00646_ net3 mod.u_cpu.rf_ram.memory\[291\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14432__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13743_ _06678_ _06456_ _06742_ _06748_ _06749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__15558__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10955_ _04766_ _04759_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13674_ _06304_ _06370_ _06682_ _06661_ _06684_ _06306_ _06685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _04720_ mod.u_cpu.rf_ram.memory\[380\]\[1\] _04717_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15413_ _01188_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13757__A2 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12625_ _05908_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14582__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _05858_ mod.u_cpu.rf_ram.memory\[162\]\[1\] _05860_ _05862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15344_ _01119_ net3 mod.u_cpu.rf_ram.memory\[399\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08633__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__I0 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13509__A2 _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11507_ _05146_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08832__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10291__I1 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15275_ _00033_ net4 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12487_ _05813_ mod.u_cpu.rf_ram.memory\[171\]\[0\] _05817_ _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12980__A3 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11031__S _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14226_ _00080_ net3 mod.u_cpu.rf_ram.memory\[574\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11438_ _05096_ mod.u_cpu.rf_ram.memory\[292\]\[0\] _05097_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14182__A2 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11966__S _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14157_ _06056_ mod.u_cpu.cpu.state.o_cnt_r\[2\] _07069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11369_ _05046_ mod.u_cpu.rf_ram.memory\[304\]\[0\] _05052_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08492__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11940__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13108_ mod.u_cpu.rf_ram.memory\[101\]\[1\] _06221_ _06239_ _06241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14088_ _03836_ _05279_ _07025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13039_ _06184_ mod.u_cpu.rf_ram.memory\[83\]\[1\] _06194_ _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15088__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09235__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12797__S _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _01745_ mod.u_cpu.rf_ram.memory\[358\]\[0\] _01907_ _01882_ _01908_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08580_ _01998_ mod.u_cpu.rf_ram.memory\[284\]\[1\] _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07531_ mod.u_cpu.rf_ram.memory\[324\]\[0\] mod.u_cpu.rf_ram.memory\[325\]\[0\] mod.u_cpu.rf_ram.memory\[326\]\[0\]
+ mod.u_cpu.rf_ram.memory\[327\]\[0\] _01837_ _01838_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07911__C _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__S _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07462_ _01741_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08872__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14925__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09201_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] _03469_
+ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11759__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09416__A3 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09132_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_33_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07427__A2 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09672__I0 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10431__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09063_ _03354_ _03365_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12037__S _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ _02293_ _02312_ _02320_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__A2 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__B1 _06474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11231__I0 mod.u_cpu.rf_ram.memory\[325\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14305__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ _04071_ mod.u_cpu.rf_ram.memory\[523\]\[1\] _04084_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08916_ _02545_ _03219_ _03222_ _02489_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14051__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09896_ _04023_ mod.u_cpu.rf_ram.memory\[534\]\[0\] _04039_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14455__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08847_ mod.u_cpu.rf_ram.memory\[32\]\[1\] mod.u_cpu.rf_ram.memory\[33\]\[1\] mod.u_cpu.rf_ram.memory\[34\]\[1\]
+ mod.u_cpu.rf_ram.memory\[35\]\[1\] _01647_ _01732_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08786__S1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13890__I _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _02325_ _03081_ _03084_ _01717_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13287__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ _01471_ _01913_ _02036_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13987__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11998__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10740_ _03737_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08863__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07666__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13739__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _04574_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12410_ _05759_ _05758_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13390_ _05784_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _06484_ _06485_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12411__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12341_ _05695_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10273__I1 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__A2 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10973__A2 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15060_ _00914_ net3 mod.u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14164__A2 _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12272_ _03755_ _05371_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14011_ _06970_ _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10025__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11222__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11223_ _04950_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13911__A2 _06890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15230__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__I1 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _04904_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04183_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11085_ _04841_ mod.u_cpu.rf_ram.memory\[34\]\[1\] _04856_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11525__I1 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10036_ _04133_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14913_ _00767_ net3 mod.u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15380__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14844_ _00698_ net3 mod.u_cpu.rf_ram.memory\[265\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14948__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13978__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14775_ _00629_ net3 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11987_ _03834_ _04068_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13726_ _06438_ _06711_ _06733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10938_ _04755_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08854__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13657_ _06361_ _06668_ _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10869_ _04708_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12789__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _05896_ _05882_ _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08606__A1 _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12402__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13588_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] mod.u_arbiter.i_wb_cpu_dbus_adr\[27\]
+ _06614_ _06615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10413__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15327_ _01104_ net3 mod.u_cpu.rf_ram.memory\[409\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10664__I _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12539_ mod.u_cpu.rf_ram.memory\[165\]\[1\] _05765_ _05849_ _05851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14328__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15258_ _00014_ net4 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12166__A1 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11213__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14209_ _02023_ _07100_ _07101_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13902__A2 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09031__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15189_ _01042_ net3 mod.u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14478__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09750_ _03930_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12713__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08701_ _02063_ _03004_ _03007_ _01669_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09681_ _03862_ mod.u_cpu.rf_ram.memory\[560\]\[1\] _03874_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07345__A1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08632_ mod.u_cpu.rf_ram.memory\[184\]\[1\] mod.u_cpu.rf_ram.memory\[185\]\[1\] mod.u_cpu.rf_ram.memory\[186\]\[1\]
+ mod.u_cpu.rf_ram.memory\[187\]\[1\] _02092_ _02098_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07440__S1 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08563_ _01697_ mod.u_cpu.rf_ram.memory\[310\]\[1\] _02869_ _01970_ _02870_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10839__I _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14091__A1 _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07514_ mod.u_cpu.rf_ram.memory\[332\]\[0\] mod.u_cpu.rf_ram.memory\[333\]\[0\] mod.u_cpu.rf_ram.memory\[334\]\[0\]
+ mod.u_cpu.rf_ram.memory\[335\]\[0\] _01819_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _01729_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14218__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15103__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ mod.u_cpu.rf_ram.memory\[392\]\[0\] mod.u_cpu.rf_ram.memory\[393\]\[0\] mod.u_cpu.rf_ram.memory\[394\]\[0\]
+ mod.u_cpu.rf_ram.memory\[395\]\[0\] _01682_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_176_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09115_ _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08073__A2 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15253__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10955__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _03349_ _03316_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08044__I _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08979__I mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07883__I _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11904__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09948_ _04075_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13657__A1 _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09879_ _04028_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11910_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10191__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A2 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12890_ _06070_ mod.u_cpu.rf_ram.memory\[89\]\[1\] _06081_ _06083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11841_ _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08219__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14560_ _00414_ net3 mod.u_cpu.rf_ram.memory\[407\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11772_ _05325_ _05301_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10723_ _04609_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13511_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _06557_ _06558_ _06566_ _06567_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_14491_ _00345_ net3 mod.u_cpu.rf_ram.memory\[442\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13188__A3 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10654_ _04563_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13442_ _03524_ _06519_ _06520_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _06523_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12396__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13373_ _06468_ _06403_ _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11443__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _04506_ mod.u_cpu.rf_ram.memory\[428\]\[0\] _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09261__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15112_ _00966_ net3 mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12324_ _05701_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12148__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14620__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15043_ _00897_ net3 mod.u_cpu.rf_ram.memory\[197\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12255_ _05645_ mod.u_cpu.rf_ram.memory\[194\]\[0\] _05654_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09013__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ _04938_ mod.u_cpu.rf_ram.memory\[32\]\[0\] _04939_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12186_ _05605_ mod.u_cpu.rf_ram.memory\[203\]\[0\] _05607_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07575__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _04893_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14770__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11068_ _04300_ _04701_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_130 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13236__S _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_141 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10019_ _04117_ mod.u_cpu.rf_ram.memory\[514\]\[0\] _04122_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_152 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_163 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10182__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_174 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__A2 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09513__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15126__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14827_ _00681_ net3 mod.u_cpu.rf_ram.memory\[274\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07461__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13035__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08827__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14758_ _00612_ net3 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13820__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13820__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13709_ _06380_ _06448_ _06717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12874__I _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14689_ _00543_ net3 mod.u_cpu.rf_ram.memory\[343\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15276__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ _01537_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _01463_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _01467_ mod.u_cpu.cpu.immdec.imm24_20\[3\]
+ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_146_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11985__I1 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08438__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13887__B2 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09802_ _03971_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07994_ _02134_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07208__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09733_ _03711_ _03745_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07318__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09664_ _03862_ mod.u_cpu.rf_ram.memory\[562\]\[1\] _03860_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08610__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08467__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08615_ _02057_ _02921_ _01632_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09595_ _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13111__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08546_ _02196_ _02844_ _02851_ _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08039__I _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08818__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15619__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12614__A2 _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10625__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11673__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _02027_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08294__A2 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _01446_ _01721_ _01735_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14643__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07359_ mod.u_cpu.rf_ram.memory\[384\]\[0\] mod.u_cpu.rf_ram.memory\[385\]\[0\] mod.u_cpu.rf_ram.memory\[386\]\[0\]
+ mod.u_cpu.rf_ram.memory\[387\]\[0\] _01664_ _01666_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _01546_ _04370_ _04371_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09029_ _03302_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13878__A1 _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14793__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12040_ _05498_ mod.u_cpu.rf_ram.memory\[60\]\[0\] _05509_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12925__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15149__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13991_ _03449_ _06952_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _06956_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07309__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__B _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12942_ _03500_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _06119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10864__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12873_ _06071_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15299__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14612_ _00466_ net3 mod.u_cpu.rf_ram.memory\[381\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11824_ _05350_ mod.u_cpu.rf_ram.memory\[22\]\[1\] _05359_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08809__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09857__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13802__A1 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15592_ _01363_ net3 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13802__B2 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14543_ _00397_ net3 mod.u_cpu.rf_ram.memory\[416\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11664__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11755_ _05314_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07788__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10706_ _04522_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14474_ _00328_ net3 mod.u_cpu.rf_ram.memory\[450\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11686_ _05250_ mod.u_cpu.rf_ram.memory\[255\]\[1\] _05264_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12369__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13425_ net5 _03677_ _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10637_ _04552_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08037__A2 _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13030__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13356_ _06426_ _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10568_ _04498_ mod.u_cpu.rf_ram.memory\[431\]\[1\] _04503_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12307_ _05689_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13869__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13287_ mod.u_arbiter.i_wb_cpu_rdt\[3\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _06377_ _06385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10499_ _04450_ mod.u_cpu.rf_ram.memory\[443\]\[1\] _04458_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15026_ _00880_ net3 mod.u_cpu.rf_ram.memory\[204\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12238_ _02299_ _05641_ _05643_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07456__C _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12169_ _02176_ _05595_ _05596_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_80 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput5 io_in[9] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_91 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14516__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12844__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ _01709_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09380_ _03616_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13921__C _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _01537_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__I1 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14666__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11655__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08276__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08262_ _02525_ _02565_ _02569_ _02539_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ mod.u_cpu.rf_ram.memory\[455\]\[0\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08193_ mod.u_cpu.rf_ram.memory\[575\]\[0\] _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ mod.u_cpu.cpu.decode.co_ebreak _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07787__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07539__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12532__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__A2 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13384__B _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ _02130_ _02284_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11683__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15441__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09647_ _03788_ _03848_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09839__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09578_ _03794_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08529_ _02148_ _02798_ _02835_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08267__A2 mod.u_cpu.rf_ram.memory\[540\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15591__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11540_ _04749_ _05149_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11271__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07401__I _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11471_ _04700_ _05120_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13012__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13210_ _06309_ _06316_ _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10422_ _04406_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12071__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14190_ _07081_ mod.u_cpu.rf_ram.memory\[244\]\[1\] _07089_ _07091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10353_ _04359_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13141_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _06258_ _06261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13072_ _06104_ _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10284_ _04266_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11326__A2 _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12023_ _05452_ _03810_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13720__B1 _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14539__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08742__A3 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13974_ _06942_ _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10137__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12925_ _06105_ mod.u_cpu.rf_ram.memory\[379\]\[1\] _06102_ _06106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14689__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09998__I _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10002__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15644_ _01415_ net3 mod.u_cpu.rf_ram.memory\[259\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12856_ mod.u_cpu.rf_ram.rdata\[1\] _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11637__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11807_ _05328_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15575_ _01346_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09455__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08889__S0 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12787_ _06014_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10065__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14526_ _00380_ net3 mod.u_cpu.rf_ram.memory\[424\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _05300_ _05301_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14457_ _00311_ net3 mod.u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10873__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13003__A2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _05254_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13408_ _06351_ mod.u_cpu.rf_ram.memory\[91\]\[0\] _06500_ _06501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14388_ _00242_ net3 mod.u_cpu.rf_ram.memory\[493\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__S0 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15314__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13339_ _06434_ _06435_ _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09238__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__I _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12514__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07900_ _02196_ _02201_ _02206_ _02207_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_15009_ _00863_ net3 mod.u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08880_ mod.u_cpu.rf_ram.memory\[568\]\[1\] mod.u_cpu.rf_ram.memory\[569\]\[1\] mod.u_cpu.rf_ram.memory\[570\]\[1\]
+ mod.u_cpu.rf_ram.memory\[571\]\[1\] _02494_ _02451_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08813__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08194__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15464__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07831_ _01746_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12599__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _01806_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_49_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09501_ _03726_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10828__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14019__A1 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13932__B _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07693_ _01998_ mod.u_cpu.rf_ram.memory\[284\]\[0\] _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08497__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11008__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09432_ _03662_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_52_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09363_ _03489_ _03603_ _03604_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08249__A2 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09446__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13223__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08314_ mod.u_cpu.rf_ram.memory\[469\]\[1\] _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09294_ _03488_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07221__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08245_ _02551_ _02552_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08761__B _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08176_ _01745_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _01435_ _01420_ _01423_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_146_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13950__B1 _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14831__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07932__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12302__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12808__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08327__I3 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _04772_ mod.u_cpu.rf_ram.memory\[366\]\[1\] _04776_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08032__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08732__I0 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12710_ _05963_ mod.u_cpu.rf_ram.memory\[7\]\[0\] _05964_ _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11492__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13690_ _06693_ _06463_ _06699_ _06409_ _06700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__14981__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08655__C _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11619__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12641_ _05886_ _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09437__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11244__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15360_ _01135_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12572_ _05872_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13784__A3 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07999__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14311_ _00165_ net3 mod.u_cpu.rf_ram.memory\[532\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15337__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11523_ _05144_ mod.u_cpu.rf_ram.memory\[27\]\[0\] _05156_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15291_ _00050_ net4 mod.u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14242_ _00096_ net3 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14194__B1 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11454_ _05108_ mod.u_cpu.rf_ram.memory\[290\]\[1\] _05103_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12744__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _04395_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14173_ _07080_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11385_ _04377_ _05062_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08412__A2 _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14361__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15487__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13124_ _06237_ mod.u_cpu.rf_ram.memory\[359\]\[1\] _06248_ _06251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10336_ _04347_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12413__S _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13055_ _06205_ mod.u_cpu.rf_ram.memory\[82\]\[0\] _06206_ _06207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10267_ _03751_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13736__C _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12006_ _05487_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10198_ _04251_ _03873_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07923__B2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13957_ _06927_ _06929_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08846__B _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07526__I1 _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12908_ _06086_ mod.u_cpu.rf_ram.memory\[97\]\[1\] _06093_ _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13888_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06640_ _06877_ _06879_ _06835_ _06880_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15627_ _01398_ net3 mod.u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12839_ _05888_ _06048_ _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15558_ _01329_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12283__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08100__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11786__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14509_ _00363_ net3 mod.u_cpu.rf_ram.memory\[433\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14075__S _07015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15489_ _01260_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08030_ mod.u_cpu.rf_ram.memory\[80\]\[0\] mod.u_cpu.rf_ram.memory\[81\]\[0\] mod.u_cpu.rf_ram.memory\[82\]\[0\]
+ mod.u_cpu.rf_ram.memory\[83\]\[0\] _02249_ _02098_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14704__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08403__A2 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10597__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09981_ _03933_ _04087_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14854__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08932_ mod.u_cpu.rf_ram.memory\[535\]\[1\] _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13696__C1 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09903__A2 _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _02472_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07914__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ _01719_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ _02202_ _03099_ _03100_ _02086_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11849__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ _01444_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07676_ _01962_ mod.u_cpu.rf_ram.memory\[276\]\[0\] _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09431__I mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07773__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14234__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09415_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03638_ _03648_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10577__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09419__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09346_ _03588_ _03590_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12792__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09277_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] _03532_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_165_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14384__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08228_ _02534_ _02535_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12726__A1 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _02120_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11201__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11170_ _04915_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10052_ _04146_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07905__A1 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14860_ _00714_ net3 mod.u_cpu.rf_ram.memory\[258\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13829__I1 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13811_ _06337_ _06811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14791_ _00645_ net3 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13742_ _06459_ _06712_ _06747_ _06423_ _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10954_ _03871_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08330__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__S0 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13673_ _06683_ _06293_ _06282_ _06294_ _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10885_ _04719_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15412_ _01187_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14727__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12624_ _05907_ mod.u_cpu.rf_ram.memory\[151\]\[1\] _05905_ _05908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07516__S0 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12965__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11768__A2 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15343_ _01118_ net3 mod.u_cpu.rf_ram.memory\[399\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12555_ _05861_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11506_ _05144_ mod.u_cpu.rf_ram.memory\[282\]\[0\] _05145_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15274_ _00032_ net4 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13509__A3 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12486_ _05606_ _05767_ _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14225_ _00001_ net3 mod.u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14877__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11437_ _04821_ _05089_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10579__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08397__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13390__A1 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14156_ _07067_ _03284_ _07068_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11368_ _04766_ _05038_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08492__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11940__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13107_ _02284_ _06239_ _06240_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10319_ _04311_ _04336_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14087_ _07024_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11299_ _04978_ mod.u_cpu.rf_ram.memory\[315\]\[0\] _05004_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09197__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14190__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13038_ _06195_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10751__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14257__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14989_ _00843_ net3 mod.u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15502__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07530_ _01503_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08321__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07461_ _01742_ _01748_ _01767_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09200_ _03472_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07392_ _01497_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12956__A1 _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _03424_ _03387_ _03427_ _03421_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09416__A4 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08624__A2 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11222__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09062_ _03356_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10431__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08013_ _01719_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08388__A1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__A1 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11231__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ _04085_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15032__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10990__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08915_ _02550_ mod.u_cpu.rf_ram.memory\[526\]\[1\] _03221_ _02515_ _03222_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09895_ _03829_ _04038_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09888__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08846_ _02365_ _03152_ _02377_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11695__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08560__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15182__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08777_ _02329_ mod.u_cpu.rf_ram.memory\[118\]\[1\] _03083_ _01916_ _03084_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11447__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12495__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07728_ _01738_ _01976_ _02035_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09161__I mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08312__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11998__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07659_ _01758_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10100__I _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10670_ _04568_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12947__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09329_ _03554_ mod.u_scanchain_local.module_data_in\[52\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08615__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12340_ _05712_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10973__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12271_ _05665_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14010_ _06909_ _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11222_ _04938_ mod.u_cpu.rf_ram.memory\[326\]\[0\] _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10770__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11153_ _04896_ mod.u_cpu.rf_ram.memory\[338\]\[1\] _04902_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09179__I0 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ _04178_ mod.u_cpu.rf_ram.memory\[502\]\[1\] _04181_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14172__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11084_ _04857_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13675__A2 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15525__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _03715_ _03717_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14912_ _00766_ net3 mod.u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12722__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14843_ _00697_ net3 mod.u_cpu.rf_ram.memory\[266\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14774_ _00628_ net3 mod.u_cpu.rf_ram.memory\[300\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11986_ _05474_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13725_ _06729_ _06730_ _06731_ _06314_ _06713_ _06732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10937_ _04753_ mod.u_cpu.rf_ram.memory\[371\]\[0\] _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13656_ _06312_ _06392_ _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10868_ _04702_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08843__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12607_ _04024_ _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13587_ _03692_ _06614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08606__A2 _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13321__I _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _04660_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15326_ _01103_ net3 mod.u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12538_ _02131_ _05849_ _05850_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07459__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15257_ _00013_ net4 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12469_ _05805_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15055__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12166__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14208_ _03775_ _07100_ _07101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15188_ _01041_ net3 mod.u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11776__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14139_ _03980_ _04996_ _07058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13115__A1 _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09246__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07593__A2 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08790__A1 _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08700_ _01573_ mod.u_cpu.rf_ram.memory\[198\]\[1\] _03006_ _02212_ _03007_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09680_ _03875_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08542__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08631_ _01818_ _02935_ _02937_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12477__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08562_ _01967_ _02868_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13940__B _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10101__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ mod.u_cpu.rf_ram.memory\[333\]\[1\] _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10652__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07444_ _01645_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10855__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07375_ _01665_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09114_ _03405_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08325__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _03253_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14422__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15548__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__I mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13106__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08781__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _04073_ mod.u_cpu.rf_ram.memory\[526\]\[0\] _04074_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13657__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09878_ _04023_ mod.u_cpu.rf_ram.memory\[537\]\[0\] _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13834__C _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14572__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08533__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ _02411_ _03135_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07832__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12468__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11840_ _03993_ _05371_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11771_ _03903_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13510_ _06564_ _06565_ _06566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _04608_ mod.u_cpu.rf_ram.memory\[406\]\[1\] _04606_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14490_ _00344_ net3 mod.u_cpu.rf_ram.memory\[442\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11840__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13441_ _06522_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10653_ _04557_ mod.u_cpu.rf_ram.memory\[417\]\[0\] _04562_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15078__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12396__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13372_ _06292_ _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08235__I _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10584_ _04233_ _04507_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15111_ _00965_ net3 mod.u_cpu.rf_ram.memory\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07272__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12323_ _05696_ mod.u_cpu.rf_ram.memory\[179\]\[0\] _05700_ _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15042_ _00896_ net3 mod.u_cpu.rf_ram.memory\[197\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12254_ _05408_ _05650_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09013__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11205_ _04808_ _03986_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12185_ _05606_ _05568_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07575__A2 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14145__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14915__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11136_ _04880_ mod.u_cpu.rf_ram.memory\[341\]\[1\] _04891_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11659__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11067_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xtiny_user_project_120 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_131 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08524__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_142 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _03975_ _04118_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_153 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_164 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_175 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14826_ _00680_ net3 mod.u_cpu.rf_ram.memory\[274\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12220__I _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14757_ _00611_ net3 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11969_ _05448_ _05462_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13820__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__B _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13708_ _06318_ _06364_ _06713_ _06715_ _06365_ _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14688_ _00542_ net3 mod.u_cpu.rf_ram.memory\[343\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13639_ mod.u_cpu.cpu.immdec.imm19_12_20\[0\] _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10675__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07160_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08145__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11434__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14445__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15309_ _00070_ net4 mod.u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13336__A1 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08438__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13887__A2 _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11898__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10945__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14595__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ _03958_ mod.u_cpu.rf_ram.memory\[547\]\[0\] _03970_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09905__S _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14136__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07993_ _02297_ mod.u_cpu.rf_ram.memory\[108\]\[0\] _02300_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09732_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12698__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12331__S _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08515__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07949__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09663_ _03763_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08610__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08614_ mod.u_cpu.rf_ram.memory\[148\]\[1\] mod.u_cpu.rf_ram.memory\[149\]\[1\] mod.u_cpu.rf_ram.memory\[150\]\[1\]
+ mod.u_cpu.rf_ram.memory\[151\]\[1\] _02059_ _01723_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09594_ _03725_ _03807_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08545_ _01886_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09866__I1 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15220__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08476_ mod.u_cpu.rf_ram.memory\[367\]\[1\] _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _01493_ _01724_ _01734_ _01534_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08055__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07358_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10389__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09243__A2 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15370__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08451__B1 _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ mod.u_cpu.rf_ram.memory\[503\]\[0\] _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07894__I _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11410__S _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14938__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09028_ _03307_ _03330_ _03251_ _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13878__A2 _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08754__A1 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13845__B _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13990_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] _06954_ _06955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12941_ _06117_ _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13136__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14318__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10864__A2 _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12872_ _06070_ mod.u_cpu.rf_ram.memory\[409\]\[1\] _06068_ _06071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14611_ _00465_ net3 mod.u_cpu.rf_ram.memory\[382\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _05360_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15591_ _01362_ net3 mod.u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14542_ _00396_ net3 mod.u_cpu.rf_ram.memory\[416\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11754_ _05311_ mod.u_cpu.rf_ram.memory\[238\]\[0\] _05313_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09482__A2 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14468__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _04597_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10495__I _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14473_ _00327_ net3 mod.u_cpu.rf_ram.memory\[451\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _02273_ _05264_ _05266_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08117__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12369__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13424_ _06510_ _06511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _04523_ mod.u_cpu.rf_ram.memory\[420\]\[0\] _04551_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13355_ _06450_ _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10567_ _01780_ _04503_ _04504_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12416__S _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _05677_ mod.u_cpu.rf_ram.memory\[186\]\[1\] _05687_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13286_ _06291_ _06293_ _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10498_ _04459_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13869__A2 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15025_ _00879_ net3 mod.u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12916__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12237_ _05642_ _05641_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__I0 _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14118__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12168_ _05322_ _05595_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10552__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11119_ _04881_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07753__B _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12099_ _05548_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08348__I1 mod.u_cpu.rf_ram.memory\[495\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_70 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_81 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_92 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11352__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15243__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14809_ _00663_ net3 mod.u_cpu.rf_ram.memory\[283\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02559_ mod.u_cpu.rf_ram.memory\[500\]\[1\] _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A3 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08261_ _02533_ mod.u_cpu.rf_ram.memory\[534\]\[0\] _02568_ _02537_ _02569_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15393__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08192_ _02216_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07236__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _01431_ _01423_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07331__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07647__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10791__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12125__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__S _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07539__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11591__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13157__S _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07976_ mod.u_cpu.rf_ram.memory\[101\]\[0\] _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09434__I mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09715_ _03870_ _03883_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11343__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _03704_ _03819_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09577_ _03764_ mod.u_cpu.rf_ram.memory\[571\]\[1\] _03792_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13096__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14610__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13796__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08528_ _01977_ _02817_ _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09464__A2 _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08459_ mod.u_cpu.rf_ram.memory\[376\]\[1\] mod.u_cpu.rf_ram.memory\[377\]\[1\] mod.u_cpu.rf_ram.memory\[378\]\[1\]
+ mod.u_cpu.rf_ram.memory\[379\]\[1\] _01957_ _01958_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11271__A2 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11204__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14760__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11470_ _05119_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10421_ _04387_ mod.u_cpu.rf_ram.memory\[455\]\[1\] _04404_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07227__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__I2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13140_ _06260_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10352_ _04345_ mod.u_cpu.rf_ram.memory\[466\]\[1\] _04357_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15116__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13071_ _06216_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10283_ _01557_ _04310_ _04312_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10909__I0 _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13720__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12022_ _05412_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11874__I _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15266__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13973_ _06914_ _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12924_ _06104_ _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14290__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12039__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08750__I1 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15643_ _01414_ net3 mod.u_cpu.rf_ram.memory\[259\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12855_ _06058_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13787__A1 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11806_ _02237_ _05347_ _05349_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15574_ _01345_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12786_ _05998_ mod.u_cpu.rf_ram.memory\[131\]\[1\] _06012_ _06014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08889__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14525_ _00379_ net3 mod.u_cpu.rf_ram.memory\[425\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11737_ _05254_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09012__C _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14456_ _00310_ net3 mod.u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11668_ _05253_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14200__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07218__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13407_ _03790_ _06344_ _06500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10619_ _03773_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14387_ _00241_ net3 mod.u_cpu.rf_ram.memory\[494\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11599_ _05199_ mod.u_cpu.rf_ram.memory\[266\]\[0\] _05206_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07313__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13338_ _06379_ _06435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08423__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11985__S _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13269_ _06298_ _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13711__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12514__A2 _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15609__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15008_ _00862_ net3 mod.u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08813__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11784__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11573__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07830_ _02136_ _02137_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08298__C _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _02046_ _02068_ _02051_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14633__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09143__A1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09500_ _03725_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _01711_ _01999_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09431_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13778__A1 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09362_ _03563_ mod.u_scanchain_local.module_data_in\[58\] _03517_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__14783__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ mod.u_cpu.rf_ram.memory\[464\]\[1\] mod.u_cpu.rf_ram.memory\[465\]\[1\] mod.u_cpu.rf_ram.memory\[466\]\[1\]
+ mod.u_cpu.rf_ram.memory\[467\]\[1\] _02593_ _02454_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12450__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _03528_ _03544_ _03545_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08244_ mod.u_cpu.rf_ram.memory\[527\]\[0\] _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15139__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _02175_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13950__A1 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ mod.u_cpu.cpu.decode.op21 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15289__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08709__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09382__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07959_ _01614_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__A1 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08001__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _04777_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09629_ _03702_ _03820_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07696__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13769__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12640_ _05917_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07791__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12816__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07412__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07448__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11244__A2 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12571_ _05869_ mod.u_cpu.rf_ram.memory\[15\]\[0\] _05871_ _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14310_ _00164_ net3 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07999__A2 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11522_ _05110_ _03791_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15290_ _00049_ net4 mod.u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14241_ _00095_ net3 mod.u_cpu.rf_ram.memory\[567\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11453_ _05107_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10773__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14506__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10404_ _04387_ mod.u_cpu.rf_ram.memory\[458\]\[1\] _04393_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12744__A2 _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08243__I _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14172_ _07057_ mod.u_cpu.rf_ram.memory\[88\]\[0\] _07079_ _07080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11384_ _03892_ _04779_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10755__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13123_ _01906_ _06248_ _06250_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10335_ _04247_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07620__A1 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13054_ _03858_ _06193_ _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10266_ _04248_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10507__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14656__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12005_ _03773_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09373__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10197_ _04250_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11180__A1 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13956_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _06906_ _06928_ _03438_ _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12907_ _06094_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13887_ _06823_ _06850_ _06878_ _06423_ _06409_ _06879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_46_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11045__S _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15626_ _01397_ net3 mod.u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12838_ _05720_ _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12432__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12769_ _06002_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15557_ _01328_ net3 mod.u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07534__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14508_ _00362_ net3 mod.u_cpu.rf_ram.memory\[433\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15488_ _01259_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14439_ _00293_ net3 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12035__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09987__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08153__I _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15431__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__S0 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13994__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11794__I0 mod.u_cpu.rf_ram.memory\[233\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04050_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09739__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ _02546_ mod.u_cpu.rf_ram.memory\[532\]\[1\] _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13696__B1 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15581__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13696__C2 _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ mod.u_cpu.rf_ram.memory\[549\]\[1\] _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _02110_ _02114_ _02119_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08793_ _02161_ mod.u_cpu.rf_ram.memory\[76\]\[1\] _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07744_ _02046_ _02050_ _02051_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _01934_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10858__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09414_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07773__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07232__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _03542_ _03538_ _03589_ _03585_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10285__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14529__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09276_ _03528_ _03530_ _03531_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ mod.u_cpu.rf_ram.memory\[519\]\[0\] _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12726__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08158_ _02461_ mod.u_cpu.rf_ram.memory\[550\]\[0\] _02464_ _02465_ _02466_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14679__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ mod.u_cpu.rf_ram_if.rtrig0 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07602__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08089_ _02302_ mod.u_cpu.rf_ram.memory\[28\]\[0\] _02396_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _03722_ _03726_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__A2 mod.u_cpu.rf_ram.memory\[550\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10051_ _04140_ mod.u_cpu.rf_ram.memory\[510\]\[1\] _04144_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11162__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A1 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14100__A1 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13810_ _06476_ _06806_ _06809_ _06810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14790_ _00644_ net3 mod.u_cpu.rf_ram.memory\[292\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13741_ _06745_ _06746_ _06462_ _06747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10953_ _04765_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15304__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08330__A2 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07764__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13672_ _06291_ _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08238__I _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10884_ _04496_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15411_ _01186_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12623_ _05873_ _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07516__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08713__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15342_ _01117_ net3 mod.u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12554_ _05855_ mod.u_cpu.rf_ram.memory\[162\]\[0\] _05860_ _05861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15454__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08094__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11505_ _04868_ _05125_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15273_ _00031_ net4 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12485_ _05816_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09969__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14224_ _00000_ net3 mod.u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11436_ _05045_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09043__B1 _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10579__I1 mod.u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09594__A1 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14155_ _06057_ _06111_ _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11367_ _05051_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13106_ _05948_ _06239_ _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10318_ _04172_ _04335_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14086_ _06904_ mod.u_cpu.rf_ram.memory\[113\]\[1\] _07022_ _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11298_ _04457_ _04990_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13319__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13037_ _06186_ mod.u_cpu.rf_ram.memory\[83\]\[0\] _06194_ _06195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10249_ _04276_ mod.u_cpu.rf_ram.memory\[481\]\[0\] _04286_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14988_ _00842_ net3 mod.u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13939_ _06913_ _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08321__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07460_ _01586_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13989__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15609_ _01380_ net3 mod.u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07391_ mod.u_cpu.rf_ram.memory\[408\]\[0\] mod.u_cpu.rf_ram.memory\[409\]\[0\] mod.u_cpu.rf_ram.memory\[410\]\[0\]
+ mod.u_cpu.rf_ram.memory\[411\]\[0\] _01697_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14086__S _07022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09130_ _03425_ _03426_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12956__A2 _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ mod.u_cpu.cpu.csr_imm _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_175_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13205__I0 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14821__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10019__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08012_ _02283_ _02315_ _02319_ _02308_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13905__A1 _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13381__A2 _06461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12334__S _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14971__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04073_ mod.u_cpu.rf_ram.memory\[523\]\[0\] _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08914_ _02551_ _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09894_ _04002_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11144__A1 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09888__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ mod.u_cpu.rf_ram.memory\[40\]\[1\] mod.u_cpu.rf_ram.memory\[41\]\[1\] mod.u_cpu.rf_ram.memory\[42\]\[1\]
+ mod.u_cpu.rf_ram.memory\[43\]\[1\] _02349_ _02393_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11695__A2 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12892__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15327__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13165__S _06274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__A2 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _01863_ _03082_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07727_ _01977_ _02009_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12644__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14351__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15477__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07658_ _01962_ mod.u_cpu.rf_ram.memory\[300\]\[0\] _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07589_ mod.u_cpu.rf_ram.memory\[367\]\[0\] _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10258__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12947__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _03574_ _03575_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_159_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14149__A1 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _03517_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__S _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12270_ _05660_ mod.u_cpu.rf_ram.memory\[192\]\[1\] _05663_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11221_ _04812_ _04945_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A3 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11152_ _04903_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10103_ _04182_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11083_ _04843_ mod.u_cpu.rf_ram.memory\[34\]\[0\] _04856_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10034_ _03662_ _03665_ _03753_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_14911_ _00765_ net3 mod.u_cpu.rf_ram.memory\[230\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10733__I1 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08551__A2 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14842_ _00696_ net3 mod.u_cpu.rf_ram.memory\[266\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11985_ _05464_ mod.u_cpu.rf_ram.memory\[216\]\[1\] _05472_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14773_ _00627_ net3 mod.u_cpu.rf_ram.memory\[301\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10497__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13724_ _06382_ _06493_ _06731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10936_ _04352_ _04733_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13655_ _06304_ _06666_ _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12419__S _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10867_ _04707_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14844__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12606_ _05895_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13586_ _06613_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13060__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10949__A1 _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10798_ mod.u_cpu.rf_ram.memory\[393\]\[0\] _04658_ _04659_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12537_ _05642_ _05849_ _05850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15325_ mod.u_cpu.cpu.o_wdata0 net3 mod.u_cpu.rf_ram_if.wdata0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14994__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07290__A2 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15256_ _00012_ net4 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12468_ _05753_ mod.u_cpu.rf_ram.memory\[419\]\[0\] _05804_ _05805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11419_ _04539_ _05020_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14207_ _03895_ _05210_ _07100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15187_ _01040_ net3 mod.u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12399_ _05745_ mod.u_cpu.rf_ram.memory\[479\]\[1\] _05750_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11374__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10421__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09527__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14138_ _06577_ _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14224__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13115__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14069_ mod.u_arbiter.i_wb_cpu_rdt\[31\] _06940_ _07013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08542__A2 _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ _02097_ _02936_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14374__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ mod.u_cpu.rf_ram.memory\[311\]\[1\] _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12626__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13823__B1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07512_ _01523_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08492_ mod.u_cpu.rf_ram.memory\[328\]\[1\] mod.u_cpu.rf_ram.memory\[329\]\[1\] mod.u_cpu.rf_ram.memory\[330\]\[1\]
+ mod.u_cpu.rf_ram.memory\[331\]\[1\] _01920_ _02666_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07443_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12329__S _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07374_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07510__I _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09113_ mod.u_arbiter.i_wb_cpu_ack _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07805__A1 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12128__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10660__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09044_ _03257_ _03296_ _03319_ _03347_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09946_ _03886_ _04062_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14717__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07416__S0 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12865__A1 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ _03996_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08533__A2 _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08384__I2 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08828_ mod.u_cpu.rf_ram.memory\[23\]\[1\] _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _02352_ _03062_ _03065_ _02361_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12468__I1 mod.u_cpu.rf_ram.memory\[419\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14867__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09089__A3 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10479__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11770_ _05324_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10721_ _04578_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13440_ _03520_ _06519_ _06520_ _03524_ _06522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10652_ _04285_ _04437_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07420__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08144__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13371_ _06463_ _06448_ _06465_ _06466_ _06467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10583_ _04515_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15110_ _00964_ net3 mod.u_cpu.rf_ram.memory\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12322_ _05037_ _05686_ _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14247__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15041_ _00895_ net3 mod.u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12253_ _05653_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11204_ _04882_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08251__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12184_ _03909_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11135_ _04892_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14397__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11108__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12156__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13648__A3 _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15642__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11066_ _03990_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_110 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11659__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_121 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_132 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10017_ _04121_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08524__A2 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_143 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_154 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_165 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_176 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12608__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14825_ _00679_ net3 mod.u_cpu.rf_ram.memory\[275\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11117__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08127__I2 mod.u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14756_ _00610_ net3 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11968_ _04025_ _05433_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__I1 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13707_ _06683_ _06667_ _06714_ _06493_ _06406_ _06715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__13408__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ _04728_ mod.u_cpu.rf_ram.memory\[374\]\[0\] _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14687_ _00541_ net3 mod.u_cpu.rf_ram.memory\[344\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11899_ _05413_ mod.u_cpu.rf_ram.memory\[225\]\[0\] _05414_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15022__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13638_ _06641_ _06648_ _06650_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07330__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13569_ _03692_ _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15308_ _00069_ net4 mod.u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08460__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15172__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15239_ _01092_ net3 mod.u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09257__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08161__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _03948_ _03969_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07992_ _02298_ _02299_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09731_ _03738_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07933__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12847__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13895__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08515__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _03861_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07949__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ _02053_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09593_ _03718_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13647__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11027__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08544_ _02295_ _02847_ _02850_ _01492_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08475_ _02022_ mod.u_cpu.rf_ram.memory\[364\]\[1\] _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07426_ _01703_ _01727_ _01733_ _01529_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15515__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07357_ _01499_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08451__A1 _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ _01556_ mod.u_cpu.rf_ram.memory\[500\]\[0\] _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _03254_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12386__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08203__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__S0 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13618__S _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _04061_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12689__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09703__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12940_ mod.u_arbiter.i_wb_cpu_rdt\[14\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _06116_ _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12871_ _06018_ _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15045__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14610_ _00464_ net3 mod.u_cpu.rf_ram.memory\[382\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _05342_ mod.u_cpu.rf_ram.memory\[22\]\[0\] _05359_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15590_ _01361_ net3 mod.u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14541_ _00395_ net3 mod.u_cpu.rf_ram.memory\[417\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _05312_ _05301_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _04593_ mod.u_cpu.rf_ram.memory\[40\]\[1\] _04595_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14472_ _00326_ net3 mod.u_cpu.rf_ram.memory\[451\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08690__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11684_ _05265_ _05264_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08117__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15195__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _04272_ _04534_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13423_ _06509_ _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13354_ _06434_ _06435_ _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10566_ _04439_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12305_ _05688_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13285_ _06367_ _06382_ _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10497_ _04453_ mod.u_cpu.rf_ram.memory\[443\]\[0\] _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11329__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12377__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12236_ _03944_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15024_ _00878_ net3 mod.u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12167_ _05593_ _05594_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13755__C _06759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11118_ _04880_ mod.u_cpu.rf_ram.memory\[344\]\[1\] _04877_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12098_ _05539_ mod.u_cpu.rf_ram.memory\[67\]\[0\] _05547_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_60 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_71 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11049_ _04827_ mod.u_cpu.rf_ram.memory\[354\]\[0\] _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_82 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_93 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14808_ _00662_ net3 mod.u_cpu.rf_ram.memory\[283\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08584__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14412__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15538__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14739_ _00593_ net3 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08276__A4 _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _02566_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08681__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07211_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _02456_ mod.u_cpu.rf_ram.memory\[572\]\[0\] _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07995__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _01432_ _01440_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14562__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08433__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11591__I1 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__C _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _02212_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09714_ _03766_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15068__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11343__I1 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ _03739_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07172__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11980__I _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _03793_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08527_ _02822_ _02824_ _02040_ _02833_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_169_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13796__A2 _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ _02759_ _02760_ _02763_ _02764_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__14905__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ mod.u_cpu.rf_ram.memory\[423\]\[1\] _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11559__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13700__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10420_ _01521_ _04404_ _04405_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07227__A2 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__I3 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ _04358_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12316__I _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13070_ _06205_ mod.u_cpu.rf_ram.memory\[81\]\[0\] _06215_ _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10282_ _04311_ _04310_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12021_ _05497_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13720__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11731__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__I _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__C _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13972_ _03446_ _06911_ _06919_ _05798_ _06941_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14435__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12923_ _06017_ _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07163__A1 mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11890__I _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15642_ _01413_ net3 mod.u_cpu.rf_ram.memory\[269\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12039__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12854_ _06057_ mod.u_cpu.rf_ram_if.rreq_r _06058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_92_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11098__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _05348_ _05347_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15573_ _01344_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12785_ _06013_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11798__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14524_ _00378_ net3 mod.u_cpu.rf_ram.memory\[425\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14585__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11736_ _03871_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10470__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14455_ _00309_ net3 mod.u_cpu.rf_ram.memory\[460\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _04226_ _05252_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13406_ _04223_ _06358_ _06498_ _06499_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08415__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _04539_ _04447_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14386_ _00240_ net3 mod.u_cpu.rf_ram.memory\[494\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11598_ _04792_ _05191_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10549_ _04492_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13337_ _06125_ _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12226__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13268_ _06318_ _06364_ _06365_ _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15007_ _00861_ net3 mod.u_cpu.rf_ram.memory\[210\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11022__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12219_ _03726_ _04226_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13199_ _06305_ _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15210__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09391__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07760_ mod.u_cpu.rf_ram.memory\[152\]\[0\] mod.u_cpu.rf_ram.memory\[153\]\[0\] mod.u_cpu.rf_ram.memory\[154\]\[0\]
+ mod.u_cpu.rf_ram.memory\[155\]\[0\] _02066_ _02067_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09143__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08577__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ mod.u_cpu.rf_ram.memory\[285\]\[0\] _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15360__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11506__S _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _03659_ _03402_ _03493_ _03660_ _03661_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14928__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11089__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09361_ _03602_ _03599_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13778__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _02592_ _02610_ _02618_ _01678_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08654__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09292_ _03535_ mod.u_scanchain_local.module_data_in\[47\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _01863_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12589__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08174_ _02478_ mod.u_cpu.rf_ram.memory\[556\]\[0\] _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ mod.u_cpu.cpu.genblk3.csr.o_new_irq _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08501__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14308__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09206__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13168__S _06274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11713__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08489__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14458__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07958_ _02058_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07889_ _01519_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09628_ _03766_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07696__A2 mod.u_cpu.rf_ram.memory\[286\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09559_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11215__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12570_ _05870_ _04913_ _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08645__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__A2 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11521_ _05155_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11151__S _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14240_ _00094_ net3 mod.u_cpu.rf_ram.memory\[567\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11452_ _05106_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14194__A2 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10403_ _04394_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10204__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14171_ _03804_ _05397_ _07079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09070__A1 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11383_ _05061_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15233__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10334_ _04346_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13122_ _06249_ _06248_ _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__A2 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11885__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13053_ _06204_ _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10265_ _04297_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12004_ _03834_ _04984_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10196_ _03808_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15383__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07384__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11180__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12504__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09125__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13955_ _06910_ _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__I3 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12906_ _06088_ mod.u_cpu.rf_ram.memory\[97\]\[0\] _06093_ _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13886_ _06382_ _06285_ _06871_ _06441_ _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09090__I _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15625_ _01396_ net3 mod.u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12837_ _06047_ _05788_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15556_ _01327_ net3 mod.u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12432__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12768_ _05998_ mod.u_cpu.rf_ram.memory\[134\]\[1\] _06000_ _06002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14507_ _00361_ net3 mod.u_cpu.rf_ram.memory\[434\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11719_ _05221_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15487_ _01258_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12699_ _05957_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14438_ _00292_ net3 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07478__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09987__I1 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13932__A2 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14369_ _00223_ net3 mod.u_cpu.rf_ram.memory\[503\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11794__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14600__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08930_ _02509_ _03236_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13696__B2 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ mod.u_cpu.rf_ram.memory\[544\]\[1\] mod.u_cpu.rf_ram.memory\[545\]\[1\] mod.u_cpu.rf_ram.memory\[546\]\[1\]
+ mod.u_cpu.rf_ram.memory\[547\]\[1\] _02450_ _02451_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__S1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07812_ _01716_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13448__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ mod.u_cpu.rf_ram.memory\[77\]\[1\] _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14750__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13448__B2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07743_ _01661_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07127__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07674_ mod.u_cpu.rf_ram.memory\[277\]\[0\] _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15106__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09413_ _03623_ _03646_ _03647_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09344_ _03570_ _03559_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_179_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10434__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11482__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09275_ _03516_ mod.u_scanchain_local.module_data_in\[44\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15256__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _02216_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08157_ _01747_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09978__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13923__A2 _06899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _02369_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07602__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14280__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13687__A1 _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10050_ _04145_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07756__I3 mod.u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14100__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13740_ _06470_ _06425_ _06458_ _06746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08866__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ _04756_ mod.u_cpu.rf_ram.memory\[36\]\[1\] _04763_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13671_ _06670_ _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10883_ _04718_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15410_ _01185_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12622_ _05906_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08618__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08682__C _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15341_ _01116_ net3 mod.u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12553_ _05408_ _05757_ _05860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08713__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08094__A2 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10976__A2 _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11504_ _05143_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15272_ _00029_ net4 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12484_ _05807_ mod.u_cpu.rf_ram.memory\[449\]\[1\] _05814_ _05816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14623__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14223_ _00079_ net3 mod.u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09043__A1 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11435_ _05095_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12705__S _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09594__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11366_ _05050_ mod.u_cpu.rf_ram.memory\[305\]\[1\] _05048_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14154_ _06063_ _07067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ _04308_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13105_ _04107_ _05640_ _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13678__A1 _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14085_ _07023_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11297_ _05003_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14773__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09085__I _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09346__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _04285_ _04137_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13036_ _05732_ _06193_ _06194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10179_ _04237_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15129__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08857__C _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14987_ _00841_ net3 mod.u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11056__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13150__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13938_ _05800_ _06909_ _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08857__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13869_ _06694_ _06438_ _06664_ _06283_ _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15279__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15608_ _01379_ net3 mod.u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08609__A1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07390_ _01500_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11464__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15539_ _01310_ net3 mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09282__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _01429_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08164__I _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__I1 mod.u_cpu.rf_ram.memory\[569\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08011_ _02316_ mod.u_cpu.rf_ram.memory\[126\]\[0\] _02318_ _02306_ _02319_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13905__A2 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07596__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09962_ _03911_ _04062_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12716__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08913_ mod.u_cpu.rf_ram.memory\[527\]\[1\] _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09893_ _04037_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07348__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11144__A2 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _02578_ _03147_ _03150_ _02660_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12892__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10869__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08775_ mod.u_cpu.rf_ram.memory\[119\]\[1\] _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13141__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07726_ _01740_ _02019_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09896__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13841__A1 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07243__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ _01963_ _01964_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07588_ _01893_ mod.u_cpu.rf_ram.memory\[364\]\[0\] _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14646__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _03569_ _03560_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _03407_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _02476_ _02512_ _02516_ _02489_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09189_ _03466_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08459__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11220_ _04948_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14796__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A4 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _04901_ mod.u_cpu.rf_ram.memory\[338\]\[0\] _04902_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__B _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10102_ _04162_ mod.u_cpu.rf_ram.memory\[502\]\[0\] _04181_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11082_ _04808_ _03975_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10033_ _04131_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14910_ _00764_ net3 mod.u_cpu.rf_ram.memory\[230\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08677__C _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14841_ _00695_ net3 mod.u_cpu.rf_ram.memory\[267\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13132__I0 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14772_ _00626_ net3 mod.u_cpu.rf_ram.memory\[301\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15421__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13832__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11984_ _05473_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07153__I _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13723_ _06362_ _06668_ _06293_ _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10646__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ _04694_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13654_ _06298_ _06299_ _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10866_ _04698_ mod.u_cpu.rf_ram.memory\[383\]\[1\] _04705_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12605_ _05891_ mod.u_cpu.rf_ram.memory\[154\]\[1\] _05893_ _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15571__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A2 mod.u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13585_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] mod.u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _06609_ _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10797_ _04527_ _04644_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10949__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15324_ _01102_ net3 mod.u_cpu.rf_ram_if.rdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11071__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12536_ _05226_ _05438_ _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15255_ _00011_ net4 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12467_ _05649_ _04437_ _05804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13899__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14206_ _06047_ _07073_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11418_ _05084_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09811__I0 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15186_ _01039_ net3 mod.u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12398_ _01562_ _05750_ _05751_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14137_ _07056_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11349_ _05037_ _05038_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08870__S0 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13774__B _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14068_ _03309_ _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13019_ _06107_ mod.u_cpu.rf_ram.memory\[10\]\[0\] _06182_ _06183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14519__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07491__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08159__I _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ _01998_ mod.u_cpu.rf_ram.memory\[308\]\[1\] _02866_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09878__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12626__A2 _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07511_ _01506_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14669__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08491_ _01848_ _02777_ _02797_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__A1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07998__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ _01509_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09112_ _03404_ _03408_ _03411_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13949__B _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09043_ _03325_ _03326_ _01394_ _03332_ _03346_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09558__A2 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07569__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09945_ _04050_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10176__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09876_ _04025_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07416__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15444__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12865__A2 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08827_ _02316_ mod.u_cpu.rf_ram.memory\[20\]\[1\] _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10876__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14067__A1 _07010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08069__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08758_ _02204_ mod.u_cpu.rf_ram.memory\[102\]\[1\] _03064_ _02359_ _03065_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09869__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10479__I1 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11676__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07709_ _01722_ mod.u_cpu.rf_ram.memory\[262\]\[0\] _02016_ _01970_ _02017_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15594__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _02202_ _02994_ _02995_ _02093_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10720_ _04607_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10651_ _04561_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11053__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13370_ _06369_ _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10582_ _04514_ mod.u_cpu.rf_ram.memory\[42\]\[1\] _04512_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12321_ _05699_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15040_ _00894_ net3 mod.u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12252_ _05635_ mod.u_cpu.rf_ram.memory\[195\]\[1\] _05651_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12553__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11203_ _04937_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12183_ _05604_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11134_ _04883_ mod.u_cpu.rf_ram.memory\[341\]\[0\] _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11065_ _04802_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_100 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_135_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_111 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _04115_ mod.u_cpu.rf_ram.memory\[515\]\[1\] _04119_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_122 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_133 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_144 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_155 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__14811__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_166 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_177 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14824_ _00678_ net3 mod.u_cpu.rf_ram.memory\[275\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13805__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08127__I3 mod.u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14755_ _00609_ net3 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11967_ _05461_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13281__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13706_ _06669_ _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10918_ _04741_ _04733_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14961__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13408__I1 mod.u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14686_ _00540_ net3 mod.u_cpu.rf_ram.memory\[344\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07611__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11898_ _04973_ _05401_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13637_ mod.u_cpu.cpu.immdec.imm31 _06649_ _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10849_ _04693_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13568_ _06603_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08835__I1 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15317__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15307_ _00068_ net4 mod.u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12519_ _05838_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08460__A2 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13499_ _06539_ _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09538__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15238_ _01091_ net3 mod.u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13592__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15169_ _01022_ net3 mod.u_cpu.rf_ram.memory\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14341__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15467__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07991_ mod.u_cpu.rf_ram.memory\[109\]\[0\] _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11509__S _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07971__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09730_ _03914_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10158__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _03847_ mod.u_cpu.rf_ram.memory\[562\]\[0\] _03860_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14049__A1 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14491__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07723__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08612_ mod.u_cpu.rf_ram.memory\[132\]\[1\] mod.u_cpu.rf_ram.memory\[133\]\[1\] mod.u_cpu.rf_ram.memory\[134\]\[1\]
+ mod.u_cpu.rf_ram.memory\[135\]\[1\] _01893_ _02054_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09592_ _03374_ _03720_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13647__I1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08543_ _02216_ mod.u_cpu.rf_ram.memory\[294\]\[1\] _02849_ _01504_ _02850_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08474_ _01729_ _02780_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _01728_ mod.u_cpu.rf_ram.memory\[406\]\[0\] _01731_ _01732_ _01733_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09228__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12139__I _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11035__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12083__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07356_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12783__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13980__B1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07287_ _01573_ _01594_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10633__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11830__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _03315_ _03327_ _03328_ _03330_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09400__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07637__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A2 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07962__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14834__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09928_ _04054_ mod.u_cpu.rf_ram.memory\[52\]\[1\] _04059_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A2 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09859_ _03809_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08762__I0 mod.u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10122__I _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12870_ _06069_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14984__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13799__B1 _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _05239_ _03829_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11649__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14540_ _00394_ net3 mod.u_cpu.rf_ram.memory\[417\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11752_ _03884_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10321__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10703_ _04596_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14471_ _00325_ net3 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12049__I _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14212__A1 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11683_ _05132_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11026__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13422_ _03377_ _03668_ net5 _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10634_ _04550_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12074__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08690__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13353_ _06448_ _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10565_ _04369_ _04447_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14364__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12304_ _05679_ mod.u_cpu.rf_ram.memory\[186\]\[0\] _05687_ _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13284_ _06368_ _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10496_ _04457_ _04443_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15023_ _00877_ net3 mod.u_cpu.rf_ram.memory\[205\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13869__A4 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12235_ _05593_ _05640_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10001__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12166_ _04379_ _05319_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11117_ _04879_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12097_ _04965_ _05543_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09093__I _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07606__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_50 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_61 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11048_ _04831_ _04822_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xtiny_user_project_72 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07705__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_83 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_94 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07800__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09821__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14807_ _00661_ net3 mod.u_cpu.rf_ram.memory\[284\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12999_ _06161_ _06164_ _06169_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09042__B _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14738_ _00592_ net3 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08130__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14669_ _00523_ net3 mod.u_cpu.rf_ram.memory\[353\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A2 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09469__S _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07210_ _01515_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08190_ _02457_ _02497_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14707__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07141_ _01449_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12765__A1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14174__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14857__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13190__A1 _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ mod.u_cpu.rf_ram.memory\[96\]\[0\] mod.u_cpu.rf_ram.memory\[97\]\[0\] mod.u_cpu.rf_ram.memory\[98\]\[0\]
+ mod.u_cpu.rf_ram.memory\[99\]\[0\] _02125_ _02127_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09713_ _03901_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11879__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11038__I _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ _03846_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09731__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14237__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09575_ _03740_ mod.u_cpu.rf_ram.memory\[571\]\[0\] _03792_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11256__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08526_ _01872_ _02825_ _02832_ _01887_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08347__I _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08457_ _01660_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14387__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ _01527_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08388_ _02692_ mod.u_cpu.rf_ram.memory\[420\]\[1\] _02694_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15632__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10350_ _04348_ mod.u_cpu.rf_ram.memory\[466\]\[0\] _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09009_ _01430_ _03313_ _03260_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__13556__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10281_ _04043_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12020_ _05484_ mod.u_cpu.rf_ram.memory\[214\]\[1\] _05495_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11031__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15012__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13971_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06940_ _06941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12922_ _06103_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08685__C _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15641_ _01412_ net3 mod.u_cpu.rf_ram.memory\[269\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15162__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12853_ _06056_ _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13163__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11804_ _05132_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15572_ _01343_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12295__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12784_ _06010_ mod.u_cpu.rf_ram.memory\[131\]\[0\] _06012_ _06013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14523_ _00377_ net3 mod.u_cpu.rf_ram.memory\[426\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11798__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11735_ _05299_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08663__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11612__S _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14454_ _00308_ net3 mod.u_cpu.rf_ram.memory\[460\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12047__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11666_ _03665_ _04224_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13405_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06413_ _06357_ _06499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _03940_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14385_ _00239_ net3 mod.u_cpu.rf_ram.memory\[495\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11597_ _05205_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ _06423_ _06430_ _06432_ _06433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10548_ _04486_ mod.u_cpu.rf_ram.memory\[434\]\[0\] _04491_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11970__A2 _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13267_ _06329_ _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10479_ _04430_ mod.u_cpu.rf_ram.memory\[446\]\[1\] _04444_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13172__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15006_ _00860_ net3 mod.u_cpu.rf_ram.memory\[210\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12218_ _05628_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11022__I1 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13198_ _06301_ _06304_ _06305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _02181_ _05580_ _05582_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15505__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10533__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07690_ _01752_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09551__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08351__A1 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11238__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12286__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__I0 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07537__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ _02611_ _02614_ _02617_ _01742_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12986__A1 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _03541_ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_61_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ _02156_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12738__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08173_ _02479_ _02480_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11321__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07124_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15035__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12910__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08590__A1 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15185__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07957_ _02170_ _02257_ _02264_ _02168_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _01851_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08342__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07145__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09627_ _03833_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09558_ _03700_ _03743_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08509_ _02665_ _02808_ _02815_ _02677_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09489_ _01460_ _03374_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_70_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11520_ _05147_ mod.u_cpu.rf_ram.memory\[280\]\[1\] _05153_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11451_ _05105_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12327__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _04365_ mod.u_cpu.rf_ram.memory\[458\]\[0\] _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10204__A2 _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14170_ _06047_ _07078_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13867__B _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11382_ _05050_ mod.u_cpu.rf_ram.memory\[302\]\[1\] _05059_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13121_ _03774_ _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10333_ _04345_ mod.u_cpu.rf_ram.memory\[46\]\[1\] _04342_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09358__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13052_ _03923_ _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11004__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12201__I0 mod.u_cpu.rf_ram.memory\[201\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ _04288_ mod.u_cpu.rf_ram.memory\[47\]\[1\] _04295_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14402__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15528__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ _05485_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10195_ _04248_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10763__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11468__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13954_ _03441_ _06917_ _06918_ _06926_ _06927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10515__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14552__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08333__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07767__S0 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12905_ _05657_ _06092_ _06093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13885_ _06735_ _06672_ _06875_ _06876_ _06877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15624_ _01395_ net3 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12268__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12836_ _06046_ _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12968__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15555_ _01326_ net3 mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12767_ _06001_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14506_ _00360_ net3 mod.u_cpu.rf_ram.memory\[434\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11718_ _05288_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15486_ _01257_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12698_ _05934_ mod.u_cpu.rf_ram.memory\[140\]\[0\] _05956_ _05957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14437_ _00291_ net3 mod.u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11649_ _05222_ mod.u_cpu.rf_ram.memory\[24\]\[0\] _05240_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11141__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15058__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13393__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14368_ _00222_ net3 mod.u_cpu.rf_ram.memory\[503\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08939__A3 _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12440__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13319_ _06415_ _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10980__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14299_ _00153_ net3 mod.u_cpu.rf_ram.memory\[538\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13696__A2 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ _01468_ _03051_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_111_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07811_ _02115_ mod.u_cpu.rf_ram.memory\[174\]\[0\] _02118_ _01771_ _02119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08791_ mod.u_cpu.rf_ram.memory\[78\]\[1\] mod.u_cpu.rf_ram.memory\[79\]\[1\] _01517_
+ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07742_ mod.u_cpu.rf_ram.memory\[144\]\[0\] mod.u_cpu.rf_ram.memory\[145\]\[0\] mod.u_cpu.rf_ram.memory\[146\]\[0\]
+ mod.u_cpu.rf_ram.memory\[147\]\[0\] _02048_ _02049_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09281__I _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07127__A2 _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10131__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ _01750_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09412_ _03439_ mod.u_scanchain_local.module_data_in\[65\] _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12959__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09343_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__A2 _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09274_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _03529_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ _02532_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13384__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08156_ _02462_ _02463_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14425__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ mod.u_cpu.rf_ram.memory\[29\]\[0\] _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13687__A2 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14575__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10745__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08563__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10370__A1 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ _03267_ _03278_ _03293_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__12498__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08315__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _04764_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10130__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13670_ _06651_ _06657_ _06681_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10882_ _04695_ mod.u_cpu.rf_ram.memory\[380\]\[0\] _04717_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12621_ _05904_ mod.u_cpu.rf_ram.memory\[151\]\[0\] _05905_ _05906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09815__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08618__A2 _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13611__A2 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15340_ _01115_ net3 mod.u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12552_ _05859_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15200__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11503_ _04959_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15271_ _00028_ net4 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12057__I _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12483_ _05815_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14222_ _00078_ net3 mod.u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11434_ mod.u_cpu.rf_ram.memory\[293\]\[1\] _05065_ _05093_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11896__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15350__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14153_ _07066_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11365_ _05031_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10984__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14175__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14918__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13104_ _06238_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10316_ _04334_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__I _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14084_ _07021_ mod.u_cpu.rf_ram.memory\[113\]\[0\] _07022_ _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11296_ _04999_ mod.u_cpu.rf_ram.memory\[316\]\[1\] _05001_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10305__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13035_ _05396_ _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10247_ _04125_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11689__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10736__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10178_ _04215_ mod.u_cpu.rf_ram.memory\[492\]\[1\] _04235_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12489__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08306__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14986_ _00840_ net3 mod.u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13937_ _05792_ _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08857__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13850__A2 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13868_ _06365_ _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15607_ _01378_ net3 mod.u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12819_ _03751_ _05721_ _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13799_ _06339_ _06790_ _06796_ _06799_ _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08609__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15538_ _01309_ net3 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14448__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15469_ _01243_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08010_ _02303_ _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12413__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14598__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _04083_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _02546_ mod.u_cpu.rf_ram.memory\[524\]\[1\] _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10215__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09892_ _04036_ mod.u_cpu.rf_ram.memory\[535\]\[1\] _04034_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__A2 _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _02191_ _03148_ _03149_ _02093_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08774_ _02477_ mod.u_cpu.rf_ram.memory\[116\]\[1\] _03080_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07524__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07725_ _01992_ _02021_ _02032_ _02007_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09896__I1 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13841__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15223__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ mod.u_cpu.rf_ram.memory\[301\]\[0\] _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10885__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07587_ _01759_ _01894_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10407__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09326_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11604__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15373__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _03495_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ _02483_ mod.u_cpu.rf_ram.memory\[566\]\[0\] _02514_ _02515_ _02516_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09188_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] _03464_
+ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08459__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ _01471_ _02382_ _02446_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08084__I0 _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07587__A2 _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ _04758_ _04887_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _04180_ _04164_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11081_ _04855_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08536__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10032_ _04115_ mod.u_cpu.rf_ram.memory\[512\]\[1\] _04129_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13436__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14840_ _00694_ net3 mod.u_cpu.rf_ram.memory\[267\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07434__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13132__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14771_ _00625_ net3 mod.u_cpu.rf_ram.memory\[302\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11983_ _05470_ mod.u_cpu.rf_ram.memory\[216\]\[0\] _05472_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13832__A2 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13722_ _06463_ _06662_ _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08395__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10934_ _04752_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11843__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13653_ _06447_ _06660_ _06663_ _06664_ _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10865_ _01865_ _04705_ _04706_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13596__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12604_ _05894_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13584_ _06612_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09264__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10796_ _03924_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_169_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15323_ _01101_ net3 mod.u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07275__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12535_ _05848_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11071__A2 _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12716__S _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15254_ _00010_ net4 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14740__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12466_ _05789_ _05803_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13899__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14205_ _07076_ _07099_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11417_ _05069_ mod.u_cpu.rf_ram.memory\[296\]\[1\] _05082_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15185_ _01038_ net3 mod.u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12397_ _05581_ _05750_ _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14136_ _07055_ mod.u_cpu.rf_ram.memory\[115\]\[1\] _07053_ _07056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11348_ _04989_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08870__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13547__S _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14890__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14067_ _07010_ _07011_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13774__C _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10709__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11279_ _04852_ _04990_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08527__A1 _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08868__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13520__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13018_ _06181_ _03919_ _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11382__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__I _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15246__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14969_ _00823_ net3 mod.u_cpu.rf_ram.memory\[575\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07510_ _01657_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08490_ _02664_ _02787_ _02796_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12882__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11834__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07502__A2 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14270__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07441_ _01498_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15396__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13081__I _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08175__I _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12634__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _03410_ mod.timer_irq _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _01432_ _03333_ _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07947__C _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12011__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07519__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08861__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04072_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09734__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09566__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08778__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13511__B2 _06566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _04024_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08826_ _02406_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10876__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08757_ _02220_ _03063_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14613__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13192__S _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07708_ _01967_ _02015_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _02179_ mod.u_cpu.rf_ram.memory\[204\]\[1\] _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _01934_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11504__I _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _04560_ mod.u_cpu.rf_ram.memory\[418\]\[1\] _04558_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14763__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07257__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09309_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _03559_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10581_ _04497_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15313__CLKN net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _05692_ mod.u_cpu.rf_ram.memory\[189\]\[1\] _05697_ _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07857__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15119__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _05652_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10056__S _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13050__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11202_ _04936_ mod.u_cpu.rf_ram.memory\[330\]\[1\] _04934_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08757__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13750__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12553__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12182_ _05309_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ _04014_ _04887_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15269__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08509__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07980__A2 _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _04842_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_101 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10015_ _04120_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_112 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_123 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_134 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_145 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_156 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14293__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_167 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14823_ _00677_ net3 mod.u_cpu.rf_ram.memory\[276\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_178 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13805__A2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11816__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11966_ _05450_ mod.u_cpu.rf_ram.memory\[539\]\[1\] _05459_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14754_ _00608_ net3 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13705_ _06317_ _06644_ _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07496__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ _03827_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14685_ _00539_ net3 mod.u_cpu.rf_ram.memory\[345\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11897_ _05412_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09312__C _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13636_ _06412_ _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _04682_ mod.u_cpu.rf_ram.memory\[385\]\[1\] _04691_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13567_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] mod.u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _06599_ _06603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10779_ _04647_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _05837_ mod.u_cpu.rf_ram.memory\[167\]\[1\] _05835_ _05838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15306_ _00067_ net4 mod.u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13498_ _06537_ _06557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12449_ _05786_ _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15237_ _01090_ net3 mod.u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08748__A1 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07339__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__S _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13592__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15168_ _01021_ net3 mod.u_cpu.rf_ram.memory\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__B _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14119_ _07045_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07990_ _01744_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15099_ _00953_ net3 mod.u_cpu.rf_ram.memory\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14636__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _03855_ _03859_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14049__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08611_ _02074_ _02917_ _01662_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__A2 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09591_ _03804_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11525__S _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08542_ _02091_ _02848_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14786__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07487__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08473_ mod.u_cpu.rf_ram.memory\[365\]\[1\] _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11324__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07424_ _01614_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07239__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07355_ _01538_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12083__I1 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13980__A1 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12783__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ mod.u_cpu.rf_ram.memory\[501\]\[0\] _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09025_ _01428_ _03328_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08739__A1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15411__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09400__A2 _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08789__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10604__S _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07962__A2 _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ _04060_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15561__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _04012_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13099__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ _01483_ _03088_ _03115_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _03960_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13799__A1 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11820_ _05358_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07712__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07478__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11751_ _05310_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _04584_ mod.u_cpu.rf_ram.memory\[40\]\[0\] _04595_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14470_ _00324_ net3 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11682_ _04700_ _05263_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14212__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13421_ _06508_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10633_ mod.u_cpu.rf_ram.memory\[421\]\[1\] _04532_ _04548_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11026__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12223__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14509__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__I _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13352_ _06316_ _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13971__A1 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10564_ _04502_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12303_ _05452_ _05686_ _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13283_ _06380_ _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10495_ _03790_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15091__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15022_ _00876_ net3 mod.u_cpu.rf_ram.memory\[205\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12234_ _03727_ _04227_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__13574__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14659__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12165_ _03894_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11116_ _04795_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12096_ _05546_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_40 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_51 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11047_ _03973_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xtiny_user_project_62 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_73 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08902__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_84 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_95 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11345__S _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14806_ _00660_ net3 mod.u_cpu.rf_ram.memory\[284\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12998_ _06164_ _06168_ _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07469__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12462__A1 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14737_ _00591_ net3 mod.u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11949_ _05405_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08130__A2 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14668_ _00522_ net3 mod.u_cpu.rf_ram.memory\[353\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12214__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13619_ _06635_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14599_ _00453_ net3 mod.u_cpu.rf_ram.memory\[388\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09549__I _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08969__A1 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15434__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07140_ _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12765__A2 _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13714__A1 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15584__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _02079_ _02147_ _01481_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09712_ mod.u_cpu.rf_ram.memory\[557\]\[1\] _03735_ _03897_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09643_ _03832_ mod.u_cpu.rf_ram.memory\[564\]\[1\] _03844_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _03758_ _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12828__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _01874_ _02828_ _02831_ _01884_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12453__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11256__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__A2 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08752__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08456_ _02711_ _02761_ _02762_ _01698_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_195_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07407_ _01709_ mod.u_cpu.rf_ram.memory\[414\]\[0\] _01713_ _01714_ _01715_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _02532_ _02693_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13253__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07338_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07632__A1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14801__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _01516_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13705__A1 _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ mod.u_cpu.cpu.alu.cmp_r _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_152_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13556__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10280_ _04307_ _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11567__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12613__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09194__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14951__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11319__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09137__A1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11229__I _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13970_ _03412_ _03614_ _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09932__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__I2 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12921_ _06088_ mod.u_cpu.rf_ram.memory\[379\]\[0\] _06102_ _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12692__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15307__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11165__S _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15640_ _01411_ net3 mod.u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12852_ _03398_ _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07442__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _04539_ _05279_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15571_ _01342_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12783_ _05649_ _06011_ _06012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14331__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14522_ _00376_ net3 mod.u_cpu.rf_ram.memory\[426\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11734_ _05287_ mod.u_cpu.rf_ram.memory\[241\]\[1\] _05297_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15457__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14453_ _00307_ net3 mod.u_cpu.rf_ram.memory\[461\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13244__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11665_ _05251_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13404_ _06483_ _06492_ _06497_ _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10616_ _04538_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14384_ _00238_ net3 mod.u_cpu.rf_ram.memory\[495\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _05194_ mod.u_cpu.rf_ram.memory\[267\]\[1\] _05203_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14481__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13335_ _06431_ _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _04201_ _04487_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12724__S _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13266_ _06361_ _06364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ _04445_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12217_ _05609_ mod.u_cpu.rf_ram.memory\[198\]\[1\] _05626_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15005_ _00859_ net3 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13197_ _06302_ _06303_ _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10230__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12148_ _05581_ _05580_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10930__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12079_ _03841_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09923__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08876__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11238__A2 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13290__S _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08310_ _02198_ mod.u_cpu.rf_ram.memory\[478\]\[1\] _02616_ _01751_ _02617_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07537__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12986__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ _03542_ _03538_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_178_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09851__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _02546_ mod.u_cpu.rf_ram.memory\[524\]\[0\] _02548_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14824__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10049__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12738__A2 _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08183__I _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08172_ mod.u_cpu.rf_ram.memory\[557\]\[0\] _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09603__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07123_ mod.u_cpu.cpu.decode.co_ebreak _01427_ _01424_ _01431_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07614__A1 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12634__S _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14974__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11549__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07955__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13529__I _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12210__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09943__S _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12910__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07956_ _02174_ _02260_ _02263_ _01766_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09742__I _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ _02188_ _02189_ _02194_ _01833_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__12674__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13264__I _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08342__A2 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14354__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09626_ _03832_ mod.u_cpu.rf_ram.memory\[566\]\[1\] _03830_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08358__I _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13218__A3 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _03777_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12809__S _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08508_ _02668_ _02811_ _02814_ _01687_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09488_ _03713_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_93_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _01770_ _02745_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10329__S _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11450_ _03732_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10401_ _04242_ _04373_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08026__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07605__A1 _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11381_ _05060_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09917__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13120_ _03941_ _04708_ _06248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10332_ _04344_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09358__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13051_ _06203_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08405__I0 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ _02439_ _04295_ _04296_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12201__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10212__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12002_ _05484_ mod.u_cpu.rf_ram.memory\[215\]\[1\] _05481_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07437__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10194_ _04247_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07464__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10763__I1 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13953_ _06920_ _05793_ _06925_ _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10515__I1 mod.u_cpu.rf_ram.memory\[440\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07767__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12904_ _05720_ _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13884_ _06492_ _06311_ _06876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15623_ _01394_ net3 mod.u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14847__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12835_ net5 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15554_ _01325_ net3 mod.u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12766_ _05992_ mod.u_cpu.rf_ram.memory\[134\]\[0\] _06000_ _06001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14505_ _00359_ net3 mod.u_cpu.rf_ram.memory\[435\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _05287_ mod.u_cpu.rf_ram.memory\[248\]\[1\] _05285_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__S _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12697_ _03904_ _05940_ _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15485_ _01256_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11422__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09099__I _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14436_ _00290_ net3 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14997__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11648_ _05239_ _03805_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__A1 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13393__A2 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14367_ _00221_ net3 mod.u_cpu.rf_ram.memory\[504\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11579_ _05177_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08939__A4 _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13318_ _06138_ _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14298_ _00152_ net3 mod.u_cpu.rf_ram.memory\[538\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14227__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13249_ _06276_ mod.u_cpu.rf_ram.memory\[92\]\[1\] _06348_ _06350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _02116_ _02117_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14377__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10702__S _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ _03090_ _03092_ _03094_ _03096_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09562__I _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15622__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07741_ _02042_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11703__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ mod.u_cpu.rf_ram.memory\[272\]\[0\] mod.u_cpu.rf_ram.memory\[273\]\[0\] mod.u_cpu.rf_ram.memory\[274\]\[0\]
+ mod.u_cpu.rf_ram.memory\[275\]\[0\] _01957_ _01958_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10131__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] _03561_ _03644_ _03645_ _03646_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12408__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09342_ _03568_ _03584_ _03586_ _03587_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_179_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12959__A2 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08088__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09273_ _03524_ _03525_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11631__A2 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13908__A1 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08224_ _01635_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15002__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13908__B2 _06889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ mod.u_cpu.rf_ram.memory\[551\]\[0\] _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08260__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ mod.u_cpu.rf_ram.memory\[24\]\[0\] mod.u_cpu.rf_ram.memory\[25\]\[0\] mod.u_cpu.rf_ram.memory\[26\]\[0\]
+ mod.u_cpu.rf_ram.memory\[27\]\[0\] _02349_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_161_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15152__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08797__B _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08563__A2 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09760__A1 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _03279_ _03292_ _03256_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09472__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10370__A2 _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07939_ _02245_ _02246_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10950_ _04753_ mod.u_cpu.rf_ram.memory\[36\]\[0\] _04763_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09609_ _03707_ _03748_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10881_ _04315_ _04709_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12620_ _03879_ _05900_ _05905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09815__A2 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12551_ _05858_ mod.u_cpu.rf_ram.memory\[163\]\[1\] _05856_ _05859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__I _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08037__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11502_ _05142_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15270_ _00027_ net4 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12482_ _05813_ mod.u_cpu.rf_ram.memory\[449\]\[0\] _05814_ _05815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A1 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14221_ _07108_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11433_ _01946_ _05093_ _05094_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11386__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14152_ _07055_ mod.u_cpu.rf_ram.memory\[247\]\[1\] _07064_ _07066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11364_ _05049_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10984__I1 mod.u_cpu.rf_ram.memory\[364\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10315_ _04330_ mod.u_cpu.rf_ram.memory\[472\]\[1\] _04332_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13103_ _06237_ mod.u_cpu.rf_ram.memory\[102\]\[1\] _06234_ _06238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14083_ _03865_ _07014_ _07022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11295_ _05002_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11138__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09583__S _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13034_ _06192_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15645__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _04284_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08003__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11689__A2 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08554__A2 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07988__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10522__S _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ _04236_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14985_ _00839_ net3 mod.u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09503__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13936_ _06910_ _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11310__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13867_ _06823_ _06449_ _06791_ _06131_ _06860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15025__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15606_ _01377_ net3 mod.u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12818_ _05962_ _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13798_ _06401_ _06798_ _06409_ _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07630__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15537_ _01308_ net3 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12248__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12749_ _05843_ _05989_ _05990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09758__S _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__A2 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A1 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15468_ _01242_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15175__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14419_ _00273_ net3 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13366__A2 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15399_ _01174_ net3 mod.u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09960_ _04071_ mod.u_cpu.rf_ram.memory\[524\]\[1\] _04081_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _02509_ _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09891_ _04017_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__A3 _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _02272_ mod.u_cpu.rf_ram.memory\[44\]\[1\] _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08773_ _01682_ _03079_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08928__S0 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07724_ _01997_ _02025_ _02031_ _02005_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07655_ _01644_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13542__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13054__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07586_ mod.u_cpu.rf_ram.memory\[365\]\[0\] _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07540__I _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09325_ _03568_ _03572_ _03573_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12801__A1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15518__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11604__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11062__I _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09256_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _03514_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14003__B1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08207_ _02306_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09187_ _03465_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13601__I0 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11368__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14542__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08138_ _01475_ _02419_ _02445_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08233__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09430__B1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09981__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08069_ _01551_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10406__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ _03828_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11080_ _04841_ mod.u_cpu.rf_ram.memory\[350\]\[1\] _04853_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12868__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14692__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _04130_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08536__A2 _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11540__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11237__I _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__S0 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10141__I _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15048__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14770_ _00624_ net3 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11982_ _05283_ _05471_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09930__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08395__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13721_ _06717_ _06727_ _06475_ _06728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10933_ _04739_ mod.u_cpu.rf_ram.memory\[372\]\[1\] _04750_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13652_ _06129_ _06664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10864_ _04611_ _04705_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14093__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07450__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15198__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12603_ _05887_ mod.u_cpu.rf_ram.memory\[154\]\[0\] _05893_ _05894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13596__A2 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13583_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] mod.u_arbiter.i_wb_cpu_dbus_adr\[25\]
+ _06609_ _06612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10795_ _04657_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08990__B _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15322_ _01100_ net3 mod.u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07275__A2 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12534_ mod.u_cpu.rf_ram.memory\[429\]\[1\] _05765_ _05846_ _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13401__B _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15253_ _00009_ net4 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12465_ _01433_ _03284_ _03377_ _05802_ _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_172_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14204_ _06153_ _07098_ _07099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11416_ _05083_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12396_ _04700_ _04335_ _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15184_ _01037_ net3 mod.u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08614__I3 mod.u_cpu.rf_ram.memory\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14135_ _06903_ _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11347_ _03849_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14066_ mod.u_arbiter.i_wb_cpu_rdt\[30\] _06937_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _04989_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10709__I1 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13627__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A2 _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10229_ _04272_ _04263_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13520__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13017_ _04982_ _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13808__B1 _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14968_ _00822_ net3 mod.u_cpu.rf_ram.memory\[575\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12331__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14415__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13919_ _03403_ _06649_ _06896_ _06897_ _06898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10986__I _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11834__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13362__I _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14899_ _00753_ net3 mod.u_cpu.rf_ram.memory\[235\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__S _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ mod.u_cpu.rf_ram.memory\[416\]\[0\] mod.u_cpu.rf_ram.memory\[417\]\[0\] mod.u_cpu.rf_ram.memory\[418\]\[0\]
+ mod.u_cpu.rf_ram.memory\[419\]\[0\] _01745_ _01747_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13036__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14084__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _01660_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11811__S _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11598__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09255__A3 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09110_ _03409_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14565__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ _03336_ _03341_ _03344_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie _03345_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_176_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11610__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12011__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__C _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04071_ mod.u_cpu.rf_ram.memory\[527\]\[1\] _04069_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _03768_ _03786_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11522__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07535__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08825_ mod.u_cpu.rf_ram.memory\[21\]\[1\] _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08756_ mod.u_cpu.rf_ram.memory\[103\]\[1\] _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08794__C _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07707_ mod.u_cpu.rf_ram.memory\[263\]\[0\] _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08687_ mod.u_cpu.rf_ram.memory\[205\]\[1\] _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15340__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13272__I _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14908__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07638_ mod.u_cpu.rf_ram.memory\[293\]\[0\] _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14075__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _01759_ _01876_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10636__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09308_ _03552_ _03547_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03543_ _03558_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_10580_ _04513_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15490__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10261__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09239_ _03499_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12389__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12250_ _05645_ mod.u_cpu.rf_ram.memory\[195\]\[0\] _05651_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10013__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ _04879_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08757__A2 _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13750__A2 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12181_ _05603_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _04890_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13447__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08509__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11063_ _04841_ mod.u_cpu.rf_ram.memory\[352\]\[1\] _04839_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07445__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _04117_ mod.u_cpu.rf_ram.memory\[515\]\[0\] _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_102 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__13891__B _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_113 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__14438__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_124 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_135 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_146 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_157 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14822_ _00676_ net3 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_168 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_179 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14753_ _00607_ net3 mod.u_cpu.rf_ram.memory\[311\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11965_ _05460_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11816__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13704_ _06470_ _06711_ _06480_ _06320_ _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__14588__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10916_ _04740_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13018__A1 _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14684_ _00538_ net3 mod.u_cpu.rf_ram.memory\[345\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11896_ _05309_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07180__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08209__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13635_ _06642_ _06645_ _06646_ _06647_ _06648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10847_ _04692_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13566_ _06602_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10778_ mod.u_cpu.rf_ram.memory\[397\]\[1\] _04532_ _04645_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15305_ _00066_ net4 mod.u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08996__A2 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12517_ _05806_ _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13497_ _06556_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15236_ _01089_ net3 mod.u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12448_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _05784_ _05785_ _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10046__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15167_ _01020_ net3 mod.u_cpu.rf_ram.memory\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12379_ _05293_ _05726_ _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15213__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14118_ _07043_ mod.u_cpu.rf_ram.memory\[11\]\[0\] _07044_ _07045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15098_ _00952_ net3 mod.u_cpu.rf_ram.memory\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14049_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _06998_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15363__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13293__S _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08610_ mod.u_cpu.rf_ram.memory\[144\]\[1\] mod.u_cpu.rf_ram.memory\[145\]\[1\] mod.u_cpu.rf_ram.memory\[146\]\[1\]
+ mod.u_cpu.rf_ram.memory\[147\]\[1\] _02085_ _02049_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09590_ _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12304__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08541_ mod.u_cpu.rf_ram.memory\[295\]\[1\] _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13092__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08186__I _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08472_ mod.u_cpu.rf_ram.memory\[360\]\[1\] mod.u_cpu.rf_ram.memory\[361\]\[1\] mod.u_cpu.rf_ram.memory\[362\]\[1\]
+ mod.u_cpu.rf_ram.memory\[363\]\[1\] _02751_ _02748_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_63_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10866__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07487__A2 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08684__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _01729_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _01661_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07239__A2 _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11291__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ mod.u_cpu.rf_ram.memory\[496\]\[0\] mod.u_cpu.rf_ram.memory\[497\]\[0\] mod.u_cpu.rf_ram.memory\[498\]\[0\]
+ mod.u_cpu.rf_ram.memory\[499\]\[0\] _01540_ _01570_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13980__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] mod.u_cpu.cpu.bufreg.lsb\[1\]
+ mod.u_cpu.cpu.bufreg.lsb\[0\] _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09936__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13267__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09926_ _04051_ mod.u_cpu.rf_ram.memory\[52\]\[0\] _04059_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13496__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07265__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13496__B2 _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ _03999_ mod.u_cpu.rf_ram.memory\[540\]\[1\] _04010_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08808_ _02337_ _03097_ _03114_ _02380_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08762__I2 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14730__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13799__A2 _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _02043_ _03042_ _03045_ _01695_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10482__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10701_ _04511_ _03933_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14880__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11681_ _05262_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13420_ _06354_ mod.u_cpu.rf_ram.memory\[339\]\[1\] _06506_ _06508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10632_ _01754_ _04548_ _04549_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12223__A2 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11282__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10563_ _04498_ mod.u_cpu.rf_ram.memory\[432\]\[1\] _04500_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13351_ _06441_ _06390_ _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08978__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13971__A2 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11982__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15236__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _05667_ _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13282_ _06328_ _06379_ _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10494_ _04456_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14220__I0 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15021_ _00875_ net3 mod.u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13723__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12233_ _05639_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12164_ _05592_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14260__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15386__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11115_ _04878_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12095_ _05533_ mod.u_cpu.rf_ram.memory\[66\]\[1\] _05544_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07175__I _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_30 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11046_ _04830_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_41 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_63 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_74 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11626__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_85 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_96 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14805_ _00659_ net3 mod.u_cpu.rf_ram.memory\[285\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11425__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12997_ _06166_ _03404_ _06167_ _05780_ _03373_ _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14736_ _00590_ net3 mod.u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07469__A2 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _02407_ _05447_ _05449_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12462__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14667_ _00521_ net3 mod.u_cpu.rf_ram.memory\[354\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11879_ _05383_ mod.u_cpu.rf_ram.memory\[71\]\[1\] _05398_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08418__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13618_ _06581_ mod.u_cpu.rf_ram.memory\[319\]\[1\] _06633_ _06635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14598_ _00452_ net3 mod.u_cpu.rf_ram.memory\[388\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13549_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] mod.u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _06589_ _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14603__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15219_ _01072_ net3 mod.u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08402__C _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ _02148_ _02232_ _02279_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14753__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _02480_ _03897_ _03900_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07157__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09642_ _03845_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15109__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09573_ _03790_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08524_ _01879_ mod.u_cpu.rf_ram.memory\[342\]\[1\] _02830_ _01867_ _02831_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08657__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13650__A1 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08455_ _01496_ mod.u_cpu.rf_ram.memory\[380\]\[1\] _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08752__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15259__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07406_ _01524_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08386_ mod.u_cpu.rf_ram.memory\[421\]\[1\] _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13402__A1 _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10216__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07337_ _01644_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11070__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _01556_ mod.u_cpu.rf_ram.memory\[468\]\[0\] _01575_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14283__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ _03308_ _03309_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11016__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13705__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07199_ _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10519__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08312__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09137__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ _04048_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12141__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__S _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12920_ _05888_ _04704_ _06102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07538__I3 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12692__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12851_ _06052_ _06055_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11802_ _05346_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15570_ _01341_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09696__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13641__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12782_ _05919_ _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14521_ _00375_ net3 mod.u_cpu.rf_ram.memory\[427\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11733_ _05298_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07320__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14452_ _00306_ net3 mod.u_cpu.rf_ram.memory\[461\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11664_ _05250_ mod.u_cpu.rf_ram.memory\[257\]\[1\] _05247_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10058__I1 mod.u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13403_ _06432_ _06403_ _06496_ _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14626__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10615_ _04537_ mod.u_cpu.rf_ram.memory\[424\]\[1\] _04535_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12076__I _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14383_ _00237_ net3 mod.u_cpu.rf_ram.memory\[496\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ _05204_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09586__S _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13334_ _06133_ _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10546_ _04490_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07623__A2 _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13265_ _06362_ _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10477_ _04423_ mod.u_cpu.rf_ram.memory\[446\]\[0\] _04444_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11707__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09385__I _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12755__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14776__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15004_ _00858_ net3 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12216_ _05627_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13196_ _05782_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _06303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12147_ _05487_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12078_ _05534_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11029_ _01903_ _04816_ _04818_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08887__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11155__I _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09687__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A1 _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15401__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14719_ _00573_ net3 mod.u_cpu.rf_ram.memory\[328\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13370__I _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07311__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08240_ _02509_ _02547_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10049__I1 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ _01925_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15551__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09064__B2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07122_ _01428_ _01429_ _01430_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_119_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13699__A1 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08413__B _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12746__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10234__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__I1 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07955_ _02249_ mod.u_cpu.rf_ram.memory\[246\]\[0\] _02262_ _02252_ _02263_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11266__S _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08878__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07886_ _02191_ _02192_ _02193_ _01666_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07543__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _03763_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10685__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13218__A4 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15081__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09556_ _03764_ mod.u_cpu.rf_ram.memory\[573\]\[1\] _03772_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14649__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08507_ _01540_ mod.u_cpu.rf_ram.memory\[326\]\[1\] _02813_ _02453_ _02814_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07302__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _03712_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08438_ mod.u_cpu.rf_ram.memory\[388\]\[1\] mod.u_cpu.rf_ram.memory\[389\]\[1\] mod.u_cpu.rf_ram.memory\[390\]\[1\]
+ mod.u_cpu.rf_ram.memory\[391\]\[1\] _02020_ _01995_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_168_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13926__A2 _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ _02668_ _02671_ _02675_ _01687_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10400_ _04392_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14799__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11380_ _05046_ mod.u_cpu.rf_ram.memory\[302\]\[0\] _05059_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _04176_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10345__S _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07718__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10262_ _04186_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13050_ _06199_ mod.u_cpu.rf_ram.memory\[79\]\[1\] _06201_ _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _05483_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _03737_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07464__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13952_ _03430_ _03433_ _03438_ _06925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15424__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12903_ _06091_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09530__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13883_ _06468_ _06874_ _06875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15622_ _01393_ net3 mod.u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12834_ _06045_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15553_ _01324_ net3 mod.u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15574__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12765_ _03950_ _05978_ _06000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14504_ _00358_ net3 mod.u_cpu.rf_ram.memory\[435\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _05249_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15484_ _01255_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12696_ _05955_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14435_ _00289_ net3 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13917__A2 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09046__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11647_ _04195_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09597__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14366_ _00220_ net3 mod.u_cpu.rf_ram.memory\[504\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11578_ _05193_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13317_ _03271_ _06358_ _06411_ _06414_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10529_ _04184_ _04447_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14297_ _00151_ net3 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09349__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13248_ _06349_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10054__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13179_ _06122_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _06286_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08887__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12105__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07780__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07740_ _02047_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13853__A1 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13853__B2 mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__I1 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12900__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07671_ _01914_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09410_ _03642_ _03638_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13605__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12408__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09341_ _03386_ mod.u_scanchain_local.module_data_in\[54\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\]
+ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09285__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09272_ _03488_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14941__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07391__S0 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08223_ _02527_ mod.u_cpu.rf_ram.memory\[516\]\[0\] _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11219__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09037__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14030__A1 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11919__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08154_ _02116_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07599__A1 _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08085_ _02126_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14321__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15447__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__I _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _03281_ _03283_ _03285_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_102_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07771__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07938_ mod.u_cpu.rf_ram.memory\[237\]\[0\] _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14471__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ _02157_ _02176_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15597__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09608_ _03787_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10880_ _04716_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11458__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09539_ _03761_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12619__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09276__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12550_ _05806_ _05858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07382__S0 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11501_ _05128_ mod.u_cpu.rf_ram.memory\[283\]\[1\] _05140_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12481_ _05657_ _04309_ _05814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14220_ _03735_ mod.u_cpu.rf_ram.memory\[249\]\[1\] _07106_ _07108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09579__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11432_ _04817_ _05093_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07876__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11386__A2 _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14151_ _02261_ _07064_ _07065_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11363_ _05046_ mod.u_cpu.rf_ram.memory\[305\]\[0\] _05048_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13102_ _06236_ _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10314_ _04333_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14082_ _06577_ _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11294_ _04978_ mod.u_cpu.rf_ram.memory\[316\]\[0\] _05001_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__B _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13033_ _06184_ mod.u_cpu.rf_ram.memory\[108\]\[1\] _06190_ _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10245_ _04267_ mod.u_cpu.rf_ram.memory\[482\]\[1\] _04282_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07892__B _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09663__I _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _04217_ mod.u_cpu.rf_ram.memory\[492\]\[0\] _04235_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14088__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08500__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14814__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14984_ _00838_ net3 mod.u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13935_ _06909_ _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09503__A2 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11634__S _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13866_ _06791_ _06672_ _06858_ _06859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14964__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15605_ _01376_ net3 mod.u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12817_ _06034_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13797_ _06383_ _06364_ _06790_ _06395_ _06797_ _06798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15536_ _01307_ net3 mod.u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12748_ _05395_ _05422_ _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08943__S _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15467_ _01241_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14012__A1 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _05312_ _05940_ _05944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08490__A2 _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09838__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14418_ _00272_ net3 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15398_ _01173_ net3 mod.u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14349_ _00203_ net3 mod.u_cpu.rf_ram.memory\[513\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14344__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08898__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08910_ mod.u_cpu.rf_ram.memory\[525\]\[1\] _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09890_ _02567_ _04034_ _04035_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10188__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09573__I _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08841_ mod.u_cpu.rf_ram.memory\[45\]\[1\] _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10888__A1 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14494__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ mod.u_cpu.rf_ram.memory\[117\]\[1\] _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13826__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ _01857_ mod.u_cpu.rf_ram.memory\[270\]\[0\] _02029_ _02030_ _02031_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08928__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07505__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07654_ _01752_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07821__I _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13054__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07585_ _01856_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _03436_ mod.u_scanchain_local.module_data_in\[51\] _03402_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12801__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10812__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _03507_ _03508_ _03503_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14003__A1 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09748__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _02484_ _02513_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09186_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] _03464_
+ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13357__A3 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07696__C _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13601__I1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ _02337_ _02425_ _02444_ _01591_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08233__A2 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__I2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10040__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__A2 _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08068_ _02352_ _02372_ _02375_ _02361_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12317__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13365__I0 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14837__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08601__B _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12868__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10030_ _04117_ mod.u_cpu.rf_ram.memory\[512\]\[0\] _04129_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09733__A2 _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07744__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08320__C _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11540__A2 _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13817__A1 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14987__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08919__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11981_ _05422_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13720_ _06726_ _06314_ _06725_ _06441_ _06727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10932_ _04751_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07731__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13651_ _06661_ _06662_ _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10863_ _04700_ _04704_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12602_ _03796_ _05882_ _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13582_ _06611_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10794_ _04641_ mod.u_cpu.rf_ram.memory\[394\]\[1\] _04655_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15321_ mod.u_cpu.rf_ram_if.rtrig0 net3 mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12533_ _01775_ _05846_ _05847_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11851__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14367__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15252_ _00077_ net4 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12464_ _05790_ _05799_ _05801_ _03686_ _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__15612__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14203_ _06152_ _06150_ _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13753__B1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ _05071_ mod.u_cpu.rf_ram.memory\[296\]\[0\] _05082_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15183_ _01036_ net3 mod.u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12395_ _05749_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09421__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14134_ _07054_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ _05036_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12308__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14065_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] _06919_ _07010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09024__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11277_ _04988_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13016_ _06180_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10228_ _03960_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10332__I _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13808__A1 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ _04221_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10590__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13808__B2 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14967_ _00821_ net3 mod.u_cpu.rf_ram.memory\[215\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13918_ _06451_ _06874_ _06487_ _06814_ _06897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_14898_ _00752_ net3 mod.u_cpu.rf_ram.memory\[235\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08160__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13849_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06455_ _06843_ _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15142__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13036__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12095__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07370_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15519_ _01290_ net3 mod.u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09660__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15292__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _03342_ _03259_ _03343_ _03344_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_129_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12547__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13744__B1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09412__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ _04017_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07816__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _03915_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11338__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07726__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11522__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08824_ mod.u_cpu.rf_ram.memory\[16\]\[1\] mod.u_cpu.rf_ram.memory\[17\]\[1\] mod.u_cpu.rf_ram.memory\[18\]\[1\]
+ mod.u_cpu.rf_ram.memory\[19\]\[1\] _02403_ _02367_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _02532_ mod.u_cpu.rf_ram.memory\[100\]\[1\] _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11274__S _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ _01998_ mod.u_cpu.rf_ram.memory\[260\]\[0\] _02013_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10333__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08686_ mod.u_cpu.rf_ram.memory\[206\]\[1\] mod.u_cpu.rf_ram.memory\[207\]\[1\] _01545_
+ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08151__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07637_ mod.u_cpu.rf_ram.memory\[288\]\[0\] mod.u_cpu.rf_ram.memory\[289\]\[0\] mod.u_cpu.rf_ram.memory\[290\]\[0\]
+ mod.u_cpu.rf_ram.memory\[291\]\[0\] _01774_ _01932_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07568_ mod.u_cpu.rf_ram.memory\[373\]\[0\] _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15635__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09307_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13983__B1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10636__I1 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_139_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09238_ _03498_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10261__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13929__S _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ _03454_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09403__A1 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__S0 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11200_ _04935_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10013__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11210__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09954__A2 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12180_ _05583_ mod.u_cpu.rf_ram.memory\[204\]\[1\] _05601_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13728__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ _04880_ mod.u_cpu.rf_ram.memory\[342\]\[1\] _04888_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15015__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11062_ _04796_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07717__A1 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10013_ _03969_ _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_103 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_114 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_125 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_136 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08390__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_147 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14821_ _00675_ net3 mod.u_cpu.rf_ram.memory\[277\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_158 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__15165__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_169 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_151_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11184__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14752_ _00606_ net3 mod.u_cpu.rf_ram.memory\[311\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11964_ _05442_ mod.u_cpu.rf_ram.memory\[539\]\[0\] _05459_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10324__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09190__I0 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13703_ _06371_ _06389_ _06711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _04739_ mod.u_cpu.rf_ram.memory\[375\]\[1\] _04737_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12079__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14683_ _00537_ net3 mod.u_cpu.rf_ram.memory\[346\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11895_ _05411_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13018__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13634_ _06455_ _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12077__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ _04679_ mod.u_cpu.rf_ram.memory\[385\]\[0\] _04691_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13565_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] mod.u_arbiter.i_wb_cpu_dbus_adr\[17\]
+ _06599_ _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10777_ _04646_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11711__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15304_ _00065_ net4 mod.u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07410__B _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12516_ _02137_ _05835_ _05836_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13496_ _03635_ _06551_ _06552_ _03642_ _06556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15235_ _01088_ net3 mod.u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12447_ _03412_ _03400_ _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15166_ _01019_ net3 mod.u_cpu.rf_ram.memory\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12378_ _05738_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07956__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14117_ _06181_ _03911_ _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11329_ _04741_ _05011_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15097_ _00951_ net3 mod.u_cpu.rf_ram.memory\[479\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14048_ _06963_ _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07708__A1 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15508__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13574__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10563__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10997__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _01807_ mod.u_cpu.rf_ram.memory\[292\]\[1\] _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14532__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10315__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07371__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__I0 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _01991_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14206__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11822__S _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ mod.u_cpu.rf_ram.memory\[407\]\[0\] _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14682__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09633__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11621__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15240__D _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07320__B _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07284_ _01445_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09023_ _03306_ _03269_ _03268_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08135__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15038__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07947__A1 _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12452__I _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09925_ _04013_ _03843_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15188__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09856_ _04011_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _03102_ _03104_ _03113_ _02664_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09787_ _03870_ _03939_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13283__I _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08738_ _02632_ mod.u_cpu.rf_ram.memory\[254\]\[1\] _03044_ _01702_ _03045_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _02711_ _02974_ _02975_ _01723_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10700_ _04594_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12059__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11680_ _05253_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12759__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13956__B1 _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ _04414_ _04548_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11531__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13350_ _06358_ _06419_ _06420_ _06446_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11431__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _04501_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__I1 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13708__B1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12301_ _05685_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11982__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13281_ _03501_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _06378_ _06379_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10493_ _04450_ mod.u_cpu.rf_ram.memory\[444\]\[1\] _04454_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13184__A1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15020_ _00874_ net3 mod.u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12232_ mod.u_cpu.rf_ram.memory\[197\]\[1\] _05617_ _05637_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14405__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12163_ mod.u_cpu.rf_ram.memory\[73\]\[1\] _05468_ _05590_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11114_ _04864_ mod.u_cpu.rf_ram.memory\[344\]\[0\] _04877_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _05545_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08996__B _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_20 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__12534__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_31 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11045_ _04825_ mod.u_cpu.rf_ram.memory\[355\]\[1\] _04828_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11498__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_42 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__14555__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10545__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_53 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08363__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_64 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_75 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_86 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_97 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14804_ _00658_ net3 mod.u_cpu.rf_ram.memory\[285\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12298__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08287__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07191__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12996_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11947_ _05448_ _05447_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14735_ _00589_ net3 mod.u_cpu.rf_ram.memory\[320\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14666_ _00520_ net3 mod.u_cpu.rf_ram.memory\[354\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11670__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11878_ _02357_ _05398_ _05399_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13617_ _01926_ _06633_ _06634_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10258__S _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10829_ _04679_ mod.u_cpu.rf_ram.memory\[388\]\[0\] _04680_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09615__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14597_ _00451_ net3 mod.u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13548_ _06592_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__A3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12981__B _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13479_ _06539_ _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15218_ _01071_ net3 mod.u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13368__I _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11089__S _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15330__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15149_ _01002_ net3 mod.u_cpu.rf_ram.memory\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10784__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07971_ _01739_ _02256_ _02278_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _03899_ _03897_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10536__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07157__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15480__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ _03802_ mod.u_cpu.rf_ram.memory\[564\]\[0\] _03844_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12289__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08197__I _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09572_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09154__I0 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _01864_ _02829_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09854__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08657__A2 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ mod.u_cpu.rf_ram.memory\[381\]\[1\] _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07969__C _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13789__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07405_ _01711_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07960__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08385_ _02220_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10216__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07336_ _01494_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11264__I1 mod.u_cpu.rf_ram.memory\[320\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14428__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07267_ _01573_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09006_ _03306_ _03307_ _03310_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_152_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07198_ mod.u_cpu.raddr\[0\] _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12182__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14578__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07276__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08593__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11727__S _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04023_ mod.u_cpu.rf_ram.memory\[532\]\[0\] _04047_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08345__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07779__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12141__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _03999_ mod.u_cpu.rf_ram.memory\[543\]\[1\] _03997_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10430__I _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12850_ _02505_ _06054_ _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _05329_ mod.u_cpu.rf_ram.memory\[232\]\[1\] _05344_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12781_ _05962_ _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14520_ _00374_ net3 mod.u_cpu.rf_ram.memory\[427\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11732_ _05289_ mod.u_cpu.rf_ram.memory\[241\]\[0\] _05297_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15203__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14451_ _00305_ net3 mod.u_cpu.rf_ram.memory\[462\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11663_ _05249_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13402_ _06381_ _06439_ _06495_ _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10614_ _04497_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14382_ _00236_ net3 mod.u_cpu.rf_ram.memory\[496\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13897__B _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11594_ _05199_ mod.u_cpu.rf_ram.memory\[267\]\[0\] _05203_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07703__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13333_ _06318_ _06428_ _06429_ _06430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15353__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10545_ _04481_ mod.u_cpu.rf_ram.memory\[435\]\[1\] _04488_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08820__A2 _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13264_ _06361_ _06362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10476_ _04299_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15003_ _00857_ net3 mod.u_cpu.rf_ram.memory\[211\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _05605_ mod.u_cpu.rf_ram.memory\[198\]\[0\] _05626_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14224__D _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13195_ _06126_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _06302_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08584__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07186__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ _05187_ _05552_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ _05533_ mod.u_cpu.rf_ram.memory\[64\]\[1\] _05531_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08336__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _04817_ _04816_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11436__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13880__A2 _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11891__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_8 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12979_ _01453_ _06152_ _06153_ _06154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14718_ _00572_ net3 mod.u_cpu.rf_ram.memory\[328\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07311__A2 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14649_ _00503_ net3 mod.u_cpu.rf_ram.memory\[363\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11171__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13396__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _02477_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09064__A2 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07121_ mod.u_cpu.cpu.csr_d_sel _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14720__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13699__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08575__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A1 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14870__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07954_ _02180_ _02261_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07885_ _01682_ mod.u_cpu.rf_ram.memory\[220\]\[0\] _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09624_ _03831_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10685__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15226__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11882__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14120__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _02497_ _03772_ _03776_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08506_ _02672_ _02812_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12682__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09486_ _03702_ _03711_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14250__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15376__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ _01680_ _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08368_ _01567_ mod.u_cpu.rf_ram.memory\[486\]\[1\] _02674_ _02109_ _02675_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_165_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07319_ _01577_ mod.u_cpu.rf_ram.memory\[486\]\[0\] _01626_ _01582_ _01627_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08299_ _01533_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10330_ _04343_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10261_ _04294_ _04068_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10748__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12000_ _05404_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08566__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10192_ _04246_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07734__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13951_ _06923_ _06924_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08869__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13862__A2 _06849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10160__I mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12902_ _06086_ mod.u_cpu.rf_ram.memory\[96\]\[1\] _06089_ _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13882_ _06858_ _06873_ _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14111__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15621_ _01392_ net3 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12833_ _06038_ mod.u_cpu.rf_ram.memory\[124\]\[1\] _06043_ _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15552_ _01323_ net3 mod.u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12764_ _05999_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14503_ _00357_ net3 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _05286_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15483_ _01254_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12695_ mod.u_cpu.rf_ram.memory\[141\]\[1\] _05950_ _05953_ _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14434_ _00288_ net3 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12425__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14743__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11646_ _05238_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09046__A2 _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11928__A2 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14365_ _00219_ net3 mod.u_cpu.rf_ram.memory\[505\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12050__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11577_ _05180_ mod.u_cpu.rf_ram.memory\[270\]\[0\] _05192_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13316_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _06413_ _06357_ _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14178__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10528_ _04478_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14296_ _00150_ net3 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14893__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10335__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13247_ _06273_ mod.u_cpu.rf_ram.memory\[92\]\[0\] _06348_ _06349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10459_ _04431_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13178_ _06284_ _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13646__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12550__I _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _05300_ _05568_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15249__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08309__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07644__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07780__A2 _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13853__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _01832_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14273__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15399__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12198__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ _03571_ _03585_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11616__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09285__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _03506_ _03526_ _03527_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11830__S _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _02528_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07391__S1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11919__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _02115_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07819__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08084_ _02384_ _02387_ _02389_ _02390_ _02391_ _01720_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10355__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _03289_ _03290_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07554__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _01681_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10107__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14616__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11076__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07868_ mod.u_cpu.rf_ram.memory\[205\]\[0\] _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10902__I0 _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08720__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _03817_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07799_ _01854_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11804__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09538_ _03732_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08385__I _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14766__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07287__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ mod.u_cpu.rf_ram_if.wdata1_r\[0\] mod.u_cpu.rf_ram_if.wdata0_r _01449_ _03695_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12280__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ _05141_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07382__S1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12480_ _05812_ _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11431_ _04412_ _05062_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10356__S _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08787__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13780__A1 _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14150_ _07026_ _07064_ _07065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11362_ _05047_ _05038_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13101_ _06017_ _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10313_ _04326_ mod.u_cpu.rf_ram.memory\[472\]\[0\] _04332_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14081_ _07020_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12571__S _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11293_ _04859_ _04990_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08539__A1 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13032_ _06191_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10244_ _04283_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08003__A3 _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13466__I _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08634__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ _04233_ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14088__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09880__S _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14296__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14983_ _00837_ net3 mod.u_cpu.rf_ram.memory\[213\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15541__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13835__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13934_ _03394_ _03280_ _06907_ _06908_ _05800_ _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_93_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13865_ _06282_ _06294_ _06305_ _06858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13599__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15604_ _01375_ net3 mod.u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07413__B _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12816_ _06019_ mod.u_cpu.rf_ram.memory\[127\]\[1\] _06031_ _06034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13796_ _06321_ _06683_ _06797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15535_ _01306_ net3 mod.u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12746__S _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12747_ _05988_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12678_ _05943_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15466_ _01240_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14417_ _00271_ net3 mod.u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12023__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _05226_ _05210_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15397_ _01172_ net3 mod.u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08778__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13771__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14348_ _00202_ net3 mod.u_cpu.rf_ram.memory\[513\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14279_ _00133_ net3 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15071__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10337__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13376__I _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14639__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ mod.u_cpu.rf_ram.memory\[46\]\[1\] mod.u_cpu.rf_ram.memory\[47\]\[1\] _01577_
+ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10888__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ mod.u_cpu.rf_ram.memory\[112\]\[1\] mod.u_cpu.rf_ram.memory\[113\]\[1\] mod.u_cpu.rf_ram.memory\[114\]\[1\]
+ mod.u_cpu.rf_ram.memory\[115\]\[1\] _01664_ _02323_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07722_ _01782_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14789__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07505__A2 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08702__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07584_ mod.u_cpu.rf_ram.memory\[360\]\[0\] mod.u_cpu.rf_ram.memory\[361\]\[0\] mod.u_cpu.rf_ram.memory\[362\]\[0\]
+ mod.u_cpu.rf_ram.memory\[363\]\[0\] _01843_ _01838_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12637__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09323_ _03569_ _03571_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _03506_ _03512_ _03513_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08205_ mod.u_cpu.rf_ram.memory\[567\]\[0\] _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09185_ _03451_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08313__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07549__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08769__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15414__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13762__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _02149_ _02434_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_147_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__I3 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ _02356_ mod.u_cpu.rf_ram.memory\[78\]\[0\] _02374_ _02359_ _02375_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09764__I _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12317__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13365__I1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__A2 _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11376__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15564__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08601__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07744__A2 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13278__B1 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ _01421_ mod.u_cpu.cpu.branch_op mod.u_cpu.cpu.csr_d_sel _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11980_ _05412_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14111__S _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _04728_ mod.u_cpu.rf_ram.memory\[372\]\[0\] _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13650_ _06320_ _06368_ _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10862_ _04703_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ _05892_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13581_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] mod.u_arbiter.i_wb_cpu_dbus_adr\[24\]
+ _06609_ _06611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _04656_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08847__I2 mod.u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12532_ _05642_ _05846_ _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15320_ _01099_ net3 mod.u_cpu.raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07887__C _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15251_ _00076_ net4 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12463_ _05800_ _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07680__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15094__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13753__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14202_ _06152_ _06151_ _07097_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11414_ _04804_ _05058_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13753__B2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15182_ _01035_ net3 mod.u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12394_ _05745_ mod.u_cpu.rf_ram.memory\[509\]\[1\] _05747_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10567__A1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14133_ _07043_ mod.u_cpu.rf_ram.memory\[115\]\[0\] _07053_ _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11345_ _05032_ mod.u_cpu.rf_ram.memory\[308\]\[1\] _05034_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12308__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14064_ _07008_ _07009_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11276_ _03755_ _04701_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09024__I2 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13015_ _06105_ mod.u_cpu.rf_ram.memory\[85\]\[1\] _06178_ _06180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10227_ _04271_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14931__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13108__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _04215_ mod.u_cpu.rf_ram.memory\[494\]\[1\] _04219_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11645__S _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10089_ _04171_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14966_ _00820_ net3 mod.u_cpu.rf_ram.memory\[215\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07922__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08535__I1 mod.u_cpu.rf_ram.memory\[297\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13917_ _06647_ _06791_ _06640_ _06896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14897_ _00751_ net3 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07594__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13848_ _06334_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _06843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13779_ _06777_ _06780_ _06331_ _06781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14311__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15437__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15518_ _01289_ net3 mod.u_cpu.rf_ram.memory\[309\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09660__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15449_ _01223_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07369__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12547__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__B2 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15587__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14461__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07423__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09941_ _02552_ _04069_ _04070_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09872_ _04022_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10030__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _02365_ _03122_ _03129_ _02185_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10730__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08754_ _02171_ _03060_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07705_ _01711_ _02012_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _02972_ _02978_ _02985_ _02991_ _01489_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08782__S0 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07636_ _01791_ _01931_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12235__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07567_ _01825_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09100__A1 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _03546_ _03553_ _03556_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13983__A1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13983__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07498_ _01603_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09237_ mod.u_cpu.cpu.genblk1.align.ctrl_misal _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14804__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09168_ mod.u_arbiter.i_wb_cpu_rdt\[12\] mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] _03452_
+ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08837__S1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08119_ mod.u_cpu.rf_ram.memory\[37\]\[0\] _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09099_ _03399_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14954__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11130_ _04889_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _04840_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10021__I0 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _03995_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08914__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A2 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_104 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_115 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_126 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_137 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14820_ _00674_ net3 mod.u_cpu.rf_ram.memory\[277\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_148 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_159 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12474__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14751_ _00605_ net3 mod.u_cpu.rf_ram.memory\[312\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11963_ _05139_ _03996_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10324__I1 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14334__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13702_ _06710_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10914_ _04719_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14682_ _00536_ net3 mod.u_cpu.rf_ram.memory\[346\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11894_ _05406_ mod.u_cpu.rf_ram.memory\[226\]\[1\] _05409_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09890__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13633_ mod.u_arbiter.i_wb_cpu_rdt\[31\] _03458_ _03503_ _06646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11029__A2 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10845_ _04285_ _04687_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13564_ _06601_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10776_ mod.u_cpu.rf_ram.memory\[397\]\[0\] _04396_ _04645_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14484__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15303_ _00064_ net4 mod.u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12515_ _05759_ _05835_ _05836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13026__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07410__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13495_ _06555_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13726__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12446_ _05783_ _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15234_ _01087_ net3 mod.u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07405__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12377_ _05729_ mod.u_cpu.rf_ram.memory\[17\]\[1\] _05736_ _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15165_ _01018_ net3 mod.u_cpu.rf_ram.memory\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14116_ _06577_ _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11328_ _05024_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15096_ _00950_ net3 mod.u_cpu.rf_ram.memory\[479\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10960__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14151__A1 _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14047_ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] _06989_ _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11259_ _04951_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07652__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14949_ _00803_ net3 mod.u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11174__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08133__A2 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _02765_ _02767_ _02776_ _01849_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14206__A2 _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07421_ _01519_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14827__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08516__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13965__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07352_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09633__A2 _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _01458_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09022_ mod.u_cpu.cpu.mem_if.signbit _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14977__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10454__S _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _04058_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09855_ _04001_ mod.u_cpu.rf_ram.memory\[540\]\[0\] _04010_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14357__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08806_ _02665_ _03105_ _03112_ _02677_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09786_ _03915_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15602__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07562__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ _02084_ _03043_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ _01567_ mod.u_cpu.rf_ram.memory\[216\]\[1\] _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13256__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07619_ _01507_ _01926_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _01672_ _02905_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08607__B _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13956__A1 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10630_ _04412_ _04528_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__12759__A2 _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10561_ _04486_ mod.u_cpu.rf_ram.memory\[432\]\[0\] _04500_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13008__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11431__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12300_ _05677_ mod.u_cpu.rf_ram.memory\[187\]\[1\] _05683_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13280_ _06377_ _03424_ _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10492_ _04455_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12231_ _02158_ _05637_ _05638_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13184__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12643__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12162_ _05591_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15132__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11990__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _04732_ _04869_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12093_ _05539_ mod.u_cpu.rf_ram.memory\[66\]\[0\] _05544_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_10 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08996__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ _04829_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_21 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_32 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_43 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11742__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_54 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_65 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__09560__A1 _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_76 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_87 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15282__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_98 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14803_ _00657_ net3 mod.u_cpu.rf_ram.memory\[286\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12447__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12995_ _03686_ _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14734_ _00588_ net3 mod.u_cpu.rf_ram.memory\[320\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11946_ _05132_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07874__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14665_ _00519_ net3 mod.u_cpu.rf_ram.memory\[355\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13247__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12818__I _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11670__A2 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11877_ _05348_ _05398_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08517__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13616_ _06249_ _06633_ _06634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10828_ _04272_ _04669_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14596_ _00450_ net3 mod.u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13547_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] mod.u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _06589_ _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10759_ _04633_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13478_ _06537_ _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13649__I _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15217_ _01070_ net3 mod.u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12429_ _01796_ _05771_ _05772_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15148_ _01001_ net3 mod.u_cpu.rf_ram.memory\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10784__I1 mod.u_cpu.rf_ram.memory\[396\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07970_ _01791_ _02265_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08679__S _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15079_ _00933_ net3 mod.u_cpu.rf_ram.memory\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15625__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09926__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12686__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10536__I1 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09640_ _03814_ _03843_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09571_ _03786_ _03788_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08106__A2 mod.u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ mod.u_cpu.rf_ram.memory\[343\]\[1\] _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09854__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08453_ mod.u_cpu.rf_ram.memory\[382\]\[1\] mod.u_cpu.rf_ram.memory\[383\]\[1\] _02125_
+ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13238__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11632__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07404_ mod.u_cpu.rf_ram.memory\[415\]\[0\] _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13938__A1 _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15005__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13789__I1 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08384_ mod.u_cpu.rf_ram.memory\[416\]\[1\] mod.u_cpu.rf_ram.memory\[417\]\[1\] mod.u_cpu.rf_ram.memory\[418\]\[1\]
+ mod.u_cpu.rf_ram.memory\[419\]\[1\] _02559_ _02155_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07960__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07335_ _01604_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10472__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07266_ mod.u_cpu.rf_ram.memory\[469\]\[0\] _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09005_ _03308_ _03309_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15155__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__I _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07197_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13410__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11972__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09790__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09907_ _03843_ _04038_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10527__I1 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08345__A2 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11807__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07779__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _03889_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09769_ _02463_ _03943_ _03946_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _05345_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12780_ _06009_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09213__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13229__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11731_ _05047_ _05284_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10359__S _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14450_ _00304_ net3 mod.u_cpu.rf_ram.memory\[462\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11662_ _05106_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13401_ _06438_ _06493_ _06494_ _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08056__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ _04536_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14381_ _00235_ net3 mod.u_cpu.rf_ram.memory\[497\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11593_ _04930_ _05191_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10463__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08900__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10544_ _04489_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13332_ _06417_ _06326_ _06330_ _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07703__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08281__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13469__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13263_ _06359_ _06360_ _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10475_ _04442_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09883__S _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14522__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15002_ _00856_ net3 mod.u_cpu.rf_ram.memory\[211\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12214_ _05355_ _05611_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08033__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13194_ _06298_ _06300_ _06301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14106__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09781__A1 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12145_ _05579_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12076_ _05483_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14672__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11027_ _03898_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15028__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_9 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13093__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12978_ _03268_ _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A2 _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A3 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14717_ _00571_ net3 mod.u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11929_ _05426_ mod.u_cpu.rf_ram.memory\[221\]\[1\] _05434_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11452__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14648_ _00502_ net3 mod.u_cpu.rf_ram.memory\[363\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15178__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14579_ _00433_ net3 mod.u_cpu.rf_ram.memory\[398\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07120_ mod.u_cpu.cpu.bne_or_bge _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10454__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10906__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11954__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ mod.u_cpu.rf_ram.memory\[247\]\[0\] _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07884_ mod.u_cpu.rf_ram.memory\[221\]\[0\] _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11182__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09623_ _03802_ mod.u_cpu.rf_ram.memory\[566\]\[0\] _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09554_ _03775_ _03772_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07840__I _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ mod.u_cpu.rf_ram.memory\[327\]\[1\] _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07838__A1 _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09485_ _03704_ _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10693__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08436_ mod.u_cpu.rf_ram.memory\[384\]\[1\] mod.u_cpu.rf_ram.memory\[385\]\[1\] mod.u_cpu.rf_ram.memory\[386\]\[1\]
+ mod.u_cpu.rf_ram.memory\[387\]\[1\] _01994_ _02010_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _02672_ _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11398__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09767__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07318_ _01578_ _01625_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14545__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08298_ _02487_ _02601_ _02604_ _02196_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07249_ mod.u_cpu.rf_ram.memory\[477\]\[0\] _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10706__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _04250_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14695__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _04245_ mod.u_cpu.rf_ram.memory\[490\]\[1\] _04243_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14114__S _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__I0 mod.u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11570__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09208__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13950_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _06906_ _06911_ _03433_ _06924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12370__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12901_ _06090_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13881_ _06426_ _06670_ _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15620_ _01391_ net3 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12832_ _06044_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__B _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13075__A1 _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07750__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15551_ _01322_ net3 mod.u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _05998_ mod.u_cpu.rf_ram.memory\[135\]\[1\] _05996_ _05999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15320__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09878__S _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14502_ _00356_ net3 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11714_ _05268_ mod.u_cpu.rf_ram.memory\[248\]\[0\] _05285_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15482_ _01253_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12694_ _05954_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14433_ _00287_ net3 mod.u_cpu.rf_ram.memory\[471\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11645_ _05234_ mod.u_cpu.rf_ram.memory\[25\]\[1\] _05236_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__I _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15470__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14364_ _00218_ net3 mod.u_cpu.rf_ram.memory\[505\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12050__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11576_ _04775_ _05191_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13315_ _06412_ _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08514__C _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10527_ _04467_ mod.u_cpu.rf_ram.memory\[438\]\[1\] _04476_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14295_ _00149_ net3 mod.u_cpu.rf_ram.memory\[540\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07197__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10458_ _04430_ mod.u_cpu.rf_ram.memory\[44\]\[1\] _04427_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13246_ _03781_ _06344_ _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13927__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13177_ mod.u_arbiter.i_wb_cpu_rdt\[11\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _05781_ _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10389_ _04233_ _04373_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12128_ _05422_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09506__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12059_ _05521_ mod.u_cpu.rf_ram.memory\[62\]\[0\] _05522_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14418__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12113__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11616__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14568__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _03516_ mod.u_scanchain_local.module_data_in\[43\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_33_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08221_ mod.u_cpu.rf_ram.memory\[517\]\[0\] _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13611__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12416__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11910__I _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08152_ _02456_ mod.u_cpu.rf_ram.memory\[548\]\[0\] _02459_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08245__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10978__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08424__C _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _01679_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08985_ mod.u_cpu.cpu.state.o_cnt_r\[1\] mod.u_cpu.cpu.state.o_cnt_r\[0\] mod.u_cpu.cpu.state.o_cnt_r\[3\]
+ mod.u_cpu.cpu.state.o_cnt_r\[2\] _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_60_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07936_ _01806_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11304__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15343__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07867_ _02134_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09606_ _03800_ mod.u_cpu.rf_ram.memory\[568\]\[1\] _03815_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07798_ _01672_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09537_ _03760_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12188__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09468_ _03683_ _03691_ _03694_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15493__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07531__I0 mod.u_cpu.rf_ram.memory\[324\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _02534_ mod.u_cpu.rf_ram.memory\[412\]\[1\] _02725_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09399_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__B _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09497__I _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11430_ _05092_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10969__I1 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08787__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _03864_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13780__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10312_ _04168_ _04327_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11791__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13100_ _06235_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11292_ _05000_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14080_ _06904_ mod.u_cpu.rf_ram.memory\[299\]\[1\] _07018_ _07020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10243_ _04276_ mod.u_cpu.rf_ram.memory\[482\]\[0\] _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13031_ _06186_ mod.u_cpu.rf_ram.memory\[108\]\[0\] _06190_ _06191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12591__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _04136_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14982_ _00836_ net3 mod.u_cpu.rf_ram.memory\[213\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12343__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13933_ _06153_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03390_ _06908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13864_ _06856_ _06857_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13048__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14710__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14096__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15603_ _01374_ net3 mod.u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12815_ _02317_ _06031_ _06033_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07413__C _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13795_ _06331_ _06794_ _06795_ _06735_ _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15534_ _01305_ net3 mod.u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09511__I1 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12746_ _05984_ mod.u_cpu.rf_ram.memory\[219\]\[1\] _05986_ _05988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08475__A1 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14860__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15465_ _01239_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12677_ _05938_ mod.u_cpu.rf_ram.memory\[143\]\[1\] _05941_ _05943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14416_ _00270_ net3 mod.u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11628_ _04106_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13220__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12023__A2 _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15396_ _01171_ net3 mod.u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08617__I3 mod.u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09975__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14347_ _00201_ net3 mod.u_cpu.rf_ram.memory\[514\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13771__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11559_ _05047_ _05171_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15216__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14278_ _00132_ net3 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13229_ mod.u_arbiter.i_wb_cpu_rdt\[30\] _03456_ _06335_ _06336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08086__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14240__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15366__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08770_ _02293_ _03069_ _03076_ _02321_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12334__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ _02027_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10896__I0 _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08702__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14390__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12002__S _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _01749_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07583_ _01890_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09322_ _03542_ _03538_ _03570_ _03559_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_80_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08466__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09253_ _03479_ mod.u_scanchain_local.module_data_in\[40\] _03408_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08204_ _02478_ mod.u_cpu.rf_ram.memory\[564\]\[0\] _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09184_ _03463_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13062__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08608__I3 mod.u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08135_ _02150_ _02435_ _02442_ _02185_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08313__S1 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13762__A2 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08066_ _01823_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10820__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12471__I _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11087__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13278__A1 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ mod.u_arbiter.i_wb_cpu_dbus_we _03263_ mod.u_cpu.cpu.immdec.imm24_20\[0\]
+ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13278__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14733__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12325__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13817__A3 _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07919_ _02070_ mod.u_cpu.rf_ram.memory\[212\]\[0\] _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11828__A2 _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08899_ _02039_ _03186_ _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15434__D _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11815__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10930_ _04749_ _04733_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14078__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14883__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10861_ _04702_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12600_ _05891_ mod.u_cpu.rf_ram.memory\[155\]\[1\] _05889_ _05892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13580_ _06610_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13450__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10792_ _04637_ mod.u_cpu.rf_ram.memory\[394\]\[0\] _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12531_ _05593_ _04528_ _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15239__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15250_ _00075_ net4 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12462_ mod.u_arbiter.i_wb_cpu_ack _03406_ _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14201_ _06152_ _06151_ _06056_ _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09957__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11413_ _05081_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15181_ _01034_ net3 mod.u_cpu.rf_ram.memory\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12393_ _01609_ _05747_ _05748_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11764__A1 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14132_ _03850_ _05631_ _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11344_ _05035_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14263__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15389__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14063_ mod.u_arbiter.i_wb_cpu_rdt\[29\] _06937_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11275_ _04987_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10319__A2 _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07475__I _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09024__I3 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13014_ _06179_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10226_ mod.u_cpu.rf_ram.memory\[485\]\[1\] _04111_ _04269_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10157_ _04220_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10088_ _04157_ mod.u_cpu.rf_ram.memory\[504\]\[1\] _04169_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14965_ _00819_ net3 mod.u_cpu.rf_ram.memory\[569\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11725__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13916_ _06894_ _06895_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08696__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14896_ _00750_ net3 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13847_ _06803_ _06841_ _06842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13816__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12757__S _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13778_ _06404_ _06744_ _06779_ _06426_ _06780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10255__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15517_ _01288_ net3 mod.u_cpu.rf_ram.memory\[309\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12729_ _05966_ mod.u_cpu.rf_ram.memory\[78\]\[1\] _05975_ _05977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15448_ _01222_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14606__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10076__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13744__A2 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15379_ _01154_ net3 mod.u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08702__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _04044_ _04069_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12291__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14756__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09871_ _04018_ mod.u_cpu.rf_ram.memory\[538\]\[1\] _04020_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _02405_ _03125_ _03128_ _02415_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13336__B _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08753_ mod.u_cpu.rf_ram.memory\[101\]\[1\] _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07704_ mod.u_cpu.rf_ram.memory\[261\]\[0\] _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14011__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08684_ _02230_ _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13680__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09105__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08782__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ _01915_ _01933_ _01942_ _01768_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13807__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08439__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12235__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _01665_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14167__B _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _03554_ mod.u_scanchain_local.module_data_in\[49\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\]
+ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13983__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07497_ _01517_ mod.u_cpu.rf_ram.memory\[444\]\[0\] _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07111__A1 mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10797__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09976__S _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09236_ _03414_ _03400_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14286__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09939__A1 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13735__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09167_ _03453_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15531__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12794__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09775__I _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08118_ mod.u_cpu.rf_ram.memory\[32\]\[0\] mod.u_cpu.rf_ram.memory\[33\]\[0\] mod.u_cpu.rf_ram.memory\[34\]\[0\]
+ mod.u_cpu.rf_ram.memory\[35\]\[0\] _02403_ _02383_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08611__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09098_ _03398_ mod.u_cpu.cpu.state.ibus_cyc _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08049_ mod.u_cpu.rf_ram.memory\[71\]\[0\] _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07295__I _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11060_ _04827_ mod.u_cpu.rf_ram.memory\[352\]\[0\] _04839_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10011_ _04050_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_105 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_116 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_127 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_138 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_149 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__11545__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14750_ _00604_ net3 mod.u_cpu.rf_ram.memory\[312\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11962_ _05458_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08678__A1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12474__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13701_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _06708_ _06709_ _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _01880_ _04737_ _04738_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14681_ _00535_ net3 mod.u_cpu.rf_ram.memory\[347\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11893_ _05410_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13632_ _06319_ _06324_ _06643_ _06644_ _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__15061__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10844_ _04690_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07898__C _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14629__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13563_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] mod.u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _06599_ _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10775_ _04643_ _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15302_ _00062_ net4 mod.u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12514_ _05395_ _05667_ _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08850__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13494_ _03631_ _06551_ _06552_ _03635_ _06555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15233_ _01086_ net3 mod.u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12445_ _05782_ _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__S _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09685__I _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14779__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15164_ _01017_ net3 mod.u_cpu.rf_ram.memory\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08602__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12376_ _05737_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14115_ _07042_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11327_ _05014_ mod.u_cpu.rf_ram.memory\[311\]\[1\] _05021_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15095_ _00949_ net3 mod.u_cpu.rf_ram.memory\[509\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09158__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14046_ _06995_ _06996_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ _04975_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13935__I _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10209_ _03942_ _04173_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08461__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11189_ _04928_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08669__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14948_ _00802_ net3 mod.u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15404__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10476__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14879_ _00733_ net3 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07341__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07420_ _01604_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__A2 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08516__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ mod.u_cpu.raddr\[2\] _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15554__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ _01486_ _01554_ _01589_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09021_ _03298_ _03255_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13717__A2 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09641__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08432__C _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09923_ _04054_ mod.u_cpu.rf_ram.memory\[530\]\[1\] _04056_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12153__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10003__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _03782_ _04003_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07843__I _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _02063_ _03108_ _03111_ _01669_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09785_ _03957_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11365__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08736_ mod.u_cpu.rf_ram.memory\[255\]\[1\] _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15084__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12700__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08667_ mod.u_cpu.rf_ram.memory\[217\]\[1\] _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__B _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07618_ mod.u_cpu.rf_ram.memory\[319\]\[0\] _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08598_ mod.u_cpu.rf_ram.memory\[263\]\[1\] _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07549_ _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_195_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10560_ _04209_ _04487_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07635__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14921__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09219_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ _04453_ mod.u_cpu.rf_ram.memory\[444\]\[0\] _04454_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12230_ _05322_ _05637_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07399__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12392__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12161_ mod.u_cpu.rf_ram.memory\[73\]\[0\] _05437_ _05590_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08691__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11112_ _04876_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12092_ _05408_ _05543_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_11 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11043_ _04827_ mod.u_cpu.rf_ram.memory\[355\]\[0\] _04828_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08899__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_22 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14301__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_33 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__15427__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13892__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_44 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_55 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_66 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_77 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_88 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_99 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14802_ _00656_ net3 mod.u_cpu.rf_ram.memory\[286\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12994_ _06165_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14733_ _00587_ net3 mod.u_cpu.rf_ram.memory\[321\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14451__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11945_ _04983_ _03837_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15577__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14664_ _00518_ net3 mod.u_cpu.rf_ram.memory\[355\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11876_ _05395_ _05397_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13615_ _04844_ _05020_ _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10827_ _04621_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10619__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14595_ _00449_ net3 mod.u_cpu.rf_ram.memory\[390\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11958__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ _06591_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10758_ _04626_ mod.u_cpu.rf_ram.memory\[400\]\[1\] _04631_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08823__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10630__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13477_ _06544_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ _04587_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15216_ _01069_ net3 mod.u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12428_ _05759_ _05771_ _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09623__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15147_ _01000_ net3 mod.u_cpu.rf_ram.memory\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10354__I _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12359_ _05666_ _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15078_ _00932_ net3 mod.u_cpu.rf_ram.memory\[182\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14029_ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] _06978_ _06984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13883__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12686__A2 _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09570_ _03787_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08521_ _01893_ mod.u_cpu.rf_ram.memory\[340\]\[1\] _02827_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _01615_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14944__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13938__A2 _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08383_ _02687_ _02689_ _02077_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09067__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14060__A1 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07334_ _01607_ mod.u_cpu.rf_ram.memory\[492\]\[0\] _01641_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09862__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10621__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07265_ _01510_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _03303_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07196_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13410__I1 mod.u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12374__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14324__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09790__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13174__I0 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09906_ _04046_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13874__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12921__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09837_ _02576_ _03997_ _03998_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14474__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09768_ _03945_ _03943_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ _02751_ mod.u_cpu.rf_ram.memory\[230\]\[1\] _03025_ _02154_ _03026_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07305__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09699_ _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _05296_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13229__I1 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10860__A1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07241__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09058__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11661_ _05248_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13400_ _06434_ _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10612_ _04523_ mod.u_cpu.rf_ram.memory\[424\]\[0\] _04535_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14380_ _00234_ net3 mod.u_cpu.rf_ram.memory\[497\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08805__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11592_ _05202_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _06424_ _06370_ _06427_ _06417_ _06428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08900__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10543_ _04486_ mod.u_cpu.rf_ram.memory\[435\]\[0\] _04488_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10375__S _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11660__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09449__B _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13262_ _05782_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10474_ _04435_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15001_ _00855_ net3 mod.u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11412__I0 mod.u_cpu.rf_ram.memory\[297\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12213_ _05625_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13193_ _06299_ _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08033__A2 _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12144_ _05566_ mod.u_cpu.rf_ram.memory\[75\]\[1\] _05577_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13165__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14817__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__I1 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08416__S0 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12075_ _05532_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10679__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _04412_ _04780_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11934__S _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14967__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12977_ _03269_ _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13093__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A4 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11928_ _02192_ _05434_ _05435_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14716_ _00570_ net3 mod.u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10151__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09203__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14647_ _00501_ net3 mod.u_cpu.rf_ram.memory\[364\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14042__A1 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11859_ _05310_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13396__A3 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14578_ _00432_ net3 mod.u_cpu.rf_ram.memory\[398\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10603__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10454__I1 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13529_ _06236_ _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11651__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10285__S _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14347__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10084__I _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__A2 mod.u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09873__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11954__I1 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14497__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07952_ _02175_ mod.u_cpu.rf_ram.memory\[244\]\[0\] _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07393__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07883_ _02190_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09622_ _03814_ _03829_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10390__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09553_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08504_ _02041_ mod.u_cpu.rf_ram.memory\[324\]\[1\] _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11095__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07838__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09484_ _03707_ _03709_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_169_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09113__I mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15122__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08435_ _02609_ _02732_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08366_ mod.u_cpu.rf_ram.memory\[487\]\[1\] _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08952__I _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11398__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07317_ mod.u_cpu.rf_ram.memory\[487\]\[0\] _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _02191_ mod.u_cpu.rf_ram.memory\[454\]\[1\] _02603_ _02093_ _02604_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_164_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15272__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07248_ _01539_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12347__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12198__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _01419_ _01443_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _04177_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07774__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11570__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12370__I1 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12900_ _06088_ mod.u_cpu.rf_ram.memory\[96\]\[0\] _06089_ _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13880_ _06811_ _06871_ _06872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12831_ _06035_ mod.u_cpu.rf_ram.memory\[124\]\[0\] _06043_ _06044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13075__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15550_ _01321_ net3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12762_ _05937_ _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14501_ _00355_ net3 mod.u_cpu.rf_ram.memory\[437\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11713_ _05283_ _05284_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08067__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15481_ _00004_ net3 mod.u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12693_ mod.u_cpu.rf_ram.memory\[141\]\[0\] _05622_ _05953_ _05954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14432_ _00286_ net3 mod.u_cpu.rf_ram.memory\[471\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11644_ _05237_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09826__I0 _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15615__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14363_ _00217_ net3 mod.u_cpu.rf_ram.memory\[506\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11575_ _05119_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07688__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13314_ _06138_ _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10526_ _04477_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14294_ _00148_ net3 mod.u_cpu.rf_ram.memory\[540\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__S _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13245_ _06347_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10457_ _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11936__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09754__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13176_ _06282_ _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10388_ _04384_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12127_ _05567_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12058_ _05428_ _03878_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08102__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _04804_ _04788_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07941__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08190__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15145__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12113__I1 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11077__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07376__S0 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14015__A1 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14015__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08220_ _01538_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15295__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12577__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08151_ _02457_ _02458_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11624__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10807__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07388__I _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08082_ mod.u_cpu.rf_ram.memory\[8\]\[0\] mod.u_cpu.rf_ram.memory\[9\]\[0\] mod.u_cpu.rf_ram.memory\[10\]\[0\]
+ mod.u_cpu.rf_ram.memory\[11\]\[0\] _02171_ _02267_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08721__B _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11001__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08984_ _03286_ _03287_ _03288_ _01421_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_87_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09108__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07935_ mod.u_cpu.rf_ram.memory\[232\]\[0\] mod.u_cpu.rf_ram.memory\[233\]\[0\] mod.u_cpu.rf_ram.memory\[234\]\[0\]
+ mod.u_cpu.rf_ram.memory\[235\]\[0\] _02242_ _02172_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07508__A1 _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _02154_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10363__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09605_ _03816_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ _01488_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _03740_ mod.u_cpu.rf_ram.memory\[574\]\[0\] _03759_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14512__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15638__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09467_ _03693_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08484__A2 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07531__I1 mod.u_cpu.rf_ram.memory\[325\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08418_ _02526_ _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ _03632_ _03633_ _03634_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14662__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _01841_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11360_ _05045_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _04331_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11791__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11291_ _04999_ mod.u_cpu.rf_ram.memory\[317\]\[1\] _04997_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08619__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15018__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13030_ _03904_ _06092_ _06190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09736__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _04281_ _04263_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12040__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10173_ _03904_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15168__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14981_ _00835_ net3 mod.u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13932_ _03268_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03279_ _03269_ _06907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13863_ mod.u_cpu.cpu.immdec.imm24_20\[2\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[3\]
+ _06857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14096__I1 mod.u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11059__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15602_ _01373_ net3 mod.u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12814_ _06032_ _06031_ _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13794_ _06726_ _06407_ _06486_ _06795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15533_ _01304_ net3 mod.u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12745_ _02199_ _05986_ _05987_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11854__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08475__A2 mod.u_cpu.rf_ram.memory\[364\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10282__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15464_ _01238_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12676_ _05942_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14415_ _00269_ net3 mod.u_cpu.rf_ram.memory\[480\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _05225_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15395_ _01170_ net3 mod.u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13220__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14346_ _00200_ net3 mod.u_cpu.rf_ram.memory\[514\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10034__A2 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09975__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11558_ _05143_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _04466_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14277_ _00131_ net3 mod.u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11489_ _01999_ _05131_ _05134_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13228_ _06334_ _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08086__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _06268_ _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07720_ mod.u_cpu.rf_ram.memory\[271\]\[0\] _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11298__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10345__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14535__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07671__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ mod.u_cpu.rf_ram.memory\[296\]\[0\] mod.u_cpu.rf_ram.memory\[297\]\[0\] mod.u_cpu.rf_ram.memory\[298\]\[0\]
+ mod.u_cpu.rf_ram.memory\[299\]\[0\] _01957_ _01958_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12098__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07582_ _01487_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09321_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03570_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13995__B1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14685__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _03507_ _03511_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08203_ _02509_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09183_ mod.u_arbiter.i_wb_cpu_rdt\[18\] mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _03459_
+ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08134_ _02155_ _02438_ _02441_ _02166_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12270__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07977__A1 _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08065_ mod.u_cpu.rf_ram.memory\[79\]\[0\] _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07846__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09718__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15310__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08967_ mod.u_arbiter.i_wb_cpu_dbus_we _03271_ _03263_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13522__I0 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07918_ mod.u_cpu.rf_ram.memory\[213\]\[0\] _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08898_ _03195_ _03204_ _02520_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15460__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07849_ _01681_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14078__I1 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12089__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10860_ _03992_ _04134_ _04701_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _03703_ _03742_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10791_ _04242_ _04648_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12530_ _05845_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08345__C _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07760__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10447__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12461_ _03359_ _03355_ _05798_ _05799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09406__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14200_ _06046_ _06151_ _07096_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_11412_ mod.u_cpu.rf_ram.memory\[297\]\[1\] _05065_ _05079_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09957__A2 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12261__I0 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15180_ _01033_ net3 mod.u_cpu.rf_ram.memory\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12392_ _05581_ _05747_ _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14408__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07968__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14131_ _07052_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11764__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _05028_ mod.u_cpu.rf_ram.memory\[308\]\[0\] _05034_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14062_ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] _07000_ _07008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11274_ _04976_ mod.u_cpu.rf_ram.memory\[31\]\[1\] _04985_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11278__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13013_ _06107_ mod.u_cpu.rf_ram.memory\[85\]\[0\] _06178_ _06179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10225_ _01622_ _04269_ _04270_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10575__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14558__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09971__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10156_ _04217_ mod.u_cpu.rf_ram.memory\[494\]\[0\] _04219_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10087_ _04170_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14964_ _00818_ net3 mod.u_cpu.rf_ram.memory\[569\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13915_ _05790_ _06413_ _06811_ _06465_ _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08535__I3 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14895_ _00749_ net3 mod.u_cpu.rf_ram.memory\[237\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13846_ _06437_ _06662_ _06840_ _06841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13816__I1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13777_ _06667_ _06778_ _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10989_ _04790_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11741__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08536__B _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10255__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15516_ _01287_ net3 mod.u_cpu.rf_ram.memory\[319\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12728_ _05976_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12659_ _05930_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15447_ _01221_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12252__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15378_ _01153_ net3 mod.u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__S _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15333__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14329_ _00183_ net3 mod.u_cpu.rf_ram.memory\[523\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08620__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09870_ _04021_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15483__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _02410_ mod.u_cpu.rf_ram.memory\[30\]\[1\] _03127_ _01830_ _03128_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ mod.u_cpu.rf_ram.memory\[96\]\[1\] mod.u_cpu.rf_ram.memory\[97\]\[1\] mod.u_cpu.rf_ram.memory\[98\]\[1\]
+ mod.u_cpu.rf_ram.memory\[99\]\[1\] _02211_ _02386_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_97_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08136__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ mod.u_cpu.rf_ram.memory\[256\]\[0\] mod.u_cpu.rf_ram.memory\[257\]\[0\] mod.u_cpu.rf_ram.memory\[258\]\[0\]
+ mod.u_cpu.rf_ram.memory\[259\]\[0\] _01994_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08683_ _02594_ _02986_ _02989_ _02591_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07634_ _01918_ _01937_ _01941_ _01929_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13807__I1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13968__B1 _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07565_ mod.u_cpu.rf_ram.memory\[368\]\[0\] mod.u_cpu.rf_ram.memory\[369\]\[0\] mod.u_cpu.rf_ram.memory\[370\]\[0\]
+ mod.u_cpu.rf_ram.memory\[371\]\[0\] _01843_ _01844_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08439__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09304_ _03407_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11294__I1 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07496_ _01802_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__A2 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07742__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10267__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09939__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ mod.u_arbiter.i_wb_cpu_rdt\[11\] mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _03452_
+ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12243__I0 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13578__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12943__A1 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ _02420_ _02422_ _02423_ _02424_ _02391_ _01552_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08998__I0 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11746__A2 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09097_ net5 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08611__A2 _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07576__I _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14700__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08048_ _01993_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10010_ _04116_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09999_ _04077_ _04108_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_106 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__13019__S _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14850__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_117 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_128 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_139 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13120__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__B1 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11961_ _05450_ mod.u_cpu.rf_ram.memory\[529\]\[1\] _05456_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__A2 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13700_ _06655_ _06709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10912_ _04611_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15206__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14680_ _00534_ net3 mod.u_cpu.rf_ram.memory\[347\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11682__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _05385_ mod.u_cpu.rf_ram.memory\[226\]\[0\] _05409_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13631_ _06371_ _06310_ _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10843_ _04682_ mod.u_cpu.rf_ram.memory\[386\]\[1\] _04688_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08356__B _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13562_ _06600_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12482__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10774_ _03723_ _04225_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_34_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14230__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12513_ _05834_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15301_ _00061_ net4 mod.u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15356__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13493_ _06554_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08850__A2 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12444_ _05781_ _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_145_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15232_ _01085_ net3 mod.u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13488__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15163_ _01016_ net3 mod.u_cpu.rf_ram.memory\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12375_ _05731_ mod.u_cpu.rf_ram.memory\[17\]\[0\] _05736_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10905__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14380__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11002__S _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14114_ _07041_ mod.u_cpu.rf_ram.memory\[87\]\[1\] _07039_ _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11326_ _01939_ _05021_ _05023_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15094_ _00948_ net3 mod.u_cpu.rf_ram.memory\[509\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14045_ mod.u_arbiter.i_wb_cpu_rdt\[24\] _06987_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _06996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11257_ _04961_ mod.u_cpu.rf_ram.memory\[321\]\[0\] _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _04258_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11188_ _04918_ mod.u_cpu.rf_ram.memory\[332\]\[0\] _04927_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08461__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11736__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _04199_ mod.u_cpu.rf_ram.memory\[497\]\[1\] _04206_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09166__I0 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14947_ _00801_ net3 mod.u_cpu.rf_ram.memory\[220\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13662__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12465__A3 _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14878_ _00732_ net3 mod.u_cpu.rf_ram.memory\[248\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07341__A2 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13829_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_arbiter.i_wb_cpu_rdt\[13\] _06335_
+ _06827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07350_ _01657_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07281_ _01446_ _01566_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09876__I _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _03323_ _03324_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14723__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13398__I _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I1 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10787__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14873__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09922_ _04057_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12153__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _04009_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10164__A1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _01511_ mod.u_cpu.rf_ram.memory\[70\]\[1\] _03110_ _02109_ _03111_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09784_ _03936_ mod.u_cpu.rf_ram.memory\[54\]\[1\] _03955_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15229__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09116__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A2 _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ _02179_ mod.u_cpu.rf_ram.memory\[252\]\[1\] _03041_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13653__A2 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ mod.u_cpu.rf_ram.memory\[218\]\[1\] mod.u_cpu.rf_ram.memory\[219\]\[1\] _02294_
+ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10711__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07999__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14253__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07617_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15379__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08597_ _02070_ mod.u_cpu.rf_ram.memory\[260\]\[1\] _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09609__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13405__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09987__S _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07548_ _01603_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07479_ mod.u_cpu.raddr\[3\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08832__A2 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _03482_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10490_ _04315_ _04443_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10725__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13101__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08596__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12160_ _05588_ _05589_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08691__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11111_ _04862_ mod.u_cpu.rf_ram.memory\[345\]\[1\] _04874_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14133__S _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12091_ _05387_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11042_ _04277_ _04822_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_12 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_23 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10155__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_34 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13892__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_45 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_56 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_67 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10950__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_78 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_89 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14801_ _00655_ net3 mod.u_cpu.rf_ram.memory\[287\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12993_ _06162_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _06164_ _06165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14732_ _00586_ net3 mod.u_cpu.rf_ram.memory\[321\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11944_ _05446_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13704__C _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10702__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08520__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14663_ _00517_ net3 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11875_ _05396_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13614_ _03313_ _03378_ _06632_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14746__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10826_ _04678_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14594_ _00448_ net3 mod.u_cpu.rf_ram.memory\[390\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11958__A2 _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12080__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13545_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] mod.u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _06589_ _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10757_ _04632_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08823__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10630__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13476_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _06538_ _06540_ _03598_ _06544_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _04579_ mod.u_cpu.rf_ram.memory\[412\]\[1\] _04585_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08533__C _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12427_ _05019_ _04442_ _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15215_ _01068_ net3 mod.u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14896__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__A3 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09623__I1 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15146_ _00999_ net3 mod.u_cpu.rf_ram.memory\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12358_ _05724_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _04989_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15077_ _00931_ net3 mod.u_cpu.rf_ram.memory\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12289_ _05677_ mod.u_cpu.rf_ram.memory\[18\]\[1\] _05675_ _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08339__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13332__A1 _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14028_ _06981_ _06983_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09000__A2 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11194__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13883__A2 _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14276__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15521__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08520_ _01858_ _02826_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _02630_ _02681_ _02722_ _02757_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08708__C _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07402_ _01509_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08382_ mod.u_cpu.rf_ram.memory\[424\]\[1\] mod.u_cpu.rf_ram.memory\[425\]\[1\] mod.u_cpu.rf_ram.memory\[426\]\[1\]
+ mod.u_cpu.rf_ram.memory\[427\]\[1\] _02688_ _02475_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_177_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09067__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14060__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07333_ _01608_ _01640_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09862__I1 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07264_ _01504_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ mod.u_cpu.cpu.alu.i_rs1 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07195_ _01498_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12374__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15051__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13323__A1 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ _04036_ mod.u_cpu.rf_ram.memory\[533\]\[1\] _04042_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14619__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13874__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09836_ _03945_ _03997_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14123__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09767_ _03944_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12201__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14769__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08718_ _01704_ _03024_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09698_ _03762_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08649_ _02130_ _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12000__I _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _05243_ mod.u_cpu.rf_ram.memory\[257\]\[0\] _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _04255_ _04534_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12935__I _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11591_ _05194_ mod.u_cpu.rf_ram.memory\[268\]\[1\] _05200_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10999__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08805__A2 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13330_ _06316_ _06426_ _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10542_ _04352_ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13261_ _06126_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _06359_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10473_ _04441_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15000_ _00854_ net3 mod.u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12212_ mod.u_cpu.rf_ram.memory\[1\]\[1\] _05617_ _05623_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13192_ mod.u_arbiter.i_wb_cpu_rdt\[15\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _03499_ _06299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11412__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07241__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12670__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12143_ _05578_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14299__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12074_ _05521_ mod.u_cpu.rf_ram.memory\[64\]\[0\] _05531_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08416__S1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11286__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15544__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__I _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11025_ _04815_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10679__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11876__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08741__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14114__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08592__I1 mod.u_cpu.rf_ram.memory\[265\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13617__A2 _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11479__I1 mod.u_cpu.rf_ram.memory\[286\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12976_ _06150_ _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14715_ _00569_ net3 mod.u_cpu.rf_ram.memory\[330\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _05348_ _05434_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10151__I1 mod.u_cpu.rf_ram.memory\[495\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11950__S _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14646_ _00500_ net3 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11858_ _05384_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14042__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10809_ _04667_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11789_ _05329_ mod.u_cpu.rf_ram.memory\[234\]\[1\] _05336_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14577_ _00431_ net3 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10603__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13528_ _06580_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08263__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13459_ _06533_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15074__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09221__A2 _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15129_ _00982_ net3 mod.u_cpu.rf_ram.memory\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07951_ _02245_ _02258_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13856__A2 _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ _02026_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14911__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09621_ _03828_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11924__I _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09552_ _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12667__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08503_ _01520_ _02809_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11095__A2 _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09483_ _01531_ _03708_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12292__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07342__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08434_ _02687_ _02733_ _02740_ _01658_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12044__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08365_ _02026_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_07316_ _01556_ mod.u_cpu.rf_ram.memory\[484\]\[0\] _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15417__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__A1 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__B2 _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08296_ _02066_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09460__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ mod.u_cpu.rf_ram.memory\[472\]\[0\] mod.u_cpu.rf_ram.memory\[473\]\[0\] mod.u_cpu.rf_ram.memory\[474\]\[0\]
+ mod.u_cpu.rf_ram.memory\[475\]\[0\] _01540_ _01501_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_165_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12347__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _01485_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14441__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15567__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08971__A1 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11158__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14591__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09819_ _03983_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10530__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12830_ _03781_ _05721_ _06043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09304__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12761_ _05997_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11330__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14500_ _00354_ net3 mod.u_cpu.rf_ram.memory\[437\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _05254_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15480_ _01252_ net3 mod.u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12692_ _04643_ _05952_ _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14431_ _00285_ net3 mod.u_cpu.rf_ram.memory\[472\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11643_ _05222_ mod.u_cpu.rf_ram.memory\[25\]\[0\] _05236_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13083__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12665__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15097__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07759__I _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14362_ _00216_ net3 mod.u_cpu.rf_ram.memory\[506\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11574_ _05190_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__A2 _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10525_ _04469_ mod.u_cpu.rf_ram.memory\[438\]\[0\] _04476_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13313_ _06338_ _06363_ _06400_ _06410_ _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14293_ _00147_ net3 mod.u_cpu.rf_ram.memory\[541\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13244_ _06276_ mod.u_cpu.rf_ram.memory\[93\]\[1\] _06345_ _06347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10456_ _04176_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10349__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07214__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13175_ _06281_ _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10387_ mod.u_cpu.rf_ram.memory\[461\]\[1\] _04383_ _04381_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07494__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07765__A2 _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14934__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12126_ _05566_ mod.u_cpu.rf_ram.memory\[20\]\[1\] _05564_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07427__C _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13838__A2 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12057_ _05520_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _03931_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11077__A2 _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10124__I1 mod.u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12959_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _05783_ _06136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14314__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07376__S1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14629_ _00483_ net3 mod.u_cpu.rf_ram.memory\[373\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08274__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07669__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08150_ mod.u_cpu.rf_ram.memory\[549\]\[0\] _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14464__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__I3 mod.u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07453__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08081_ mod.u_cpu.rf_ram.memory\[12\]\[0\] mod.u_cpu.rf_ram.memory\[13\]\[0\] mod.u_cpu.rf_ram.memory\[14\]\[0\]
+ mod.u_cpu.rf_ram.memory\[15\]\[0\] _02266_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13526__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07205__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08721__C _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11001__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ mod.u_cpu.cpu.branch_op _03254_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__10760__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07934_ _01604_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12888__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07865_ mod.u_cpu.rf_ram.memory\[200\]\[0\] mod.u_cpu.rf_ram.memory\[201\]\[0\] mod.u_cpu.rf_ram.memory\[202\]\[0\]
+ mod.u_cpu.rf_ram.memory\[203\]\[0\] _02171_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08449__B _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ _03802_ mod.u_cpu.rf_ram.memory\[568\]\[0\] _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07796_ _01458_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09535_ _03752_ _03758_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10115__I1 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13802__C _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08417_ mod.u_cpu.rf_ram.memory\[413\]\[1\] _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12017__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07692__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13065__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14807__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09397_ _03386_ mod.u_scanchain_local.module_data_in\[63\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__B _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07579__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08348_ mod.u_cpu.rf_ram.memory\[494\]\[1\] mod.u_cpu.rf_ram.memory\[495\]\[1\] _01709_
+ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08279_ mod.u_cpu.rf_ram.memory\[462\]\[1\] mod.u_cpu.rf_ram.memory\[463\]\[1\] _02585_
+ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10310_ _04330_ mod.u_cpu.rf_ram.memory\[473\]\[1\] _04328_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14957__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11290_ _04951_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08619__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10241_ _03974_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10051__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09992__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _04232_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14980_ _00834_ net3 mod.u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12879__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13931_ _05801_ _06906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14337__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13862_ _06814_ _06849_ _06855_ _06704_ _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_74_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__I mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15601_ _01372_ net3 mod.u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11059__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12813_ _03774_ _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13793_ _06779_ _06792_ _06793_ _06776_ _06794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15532_ _01303_ net3 mod.u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12744_ _05843_ _05986_ _05987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13712__C _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14487__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08806__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15463_ _01237_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12675_ _05934_ mod.u_cpu.rf_ram.memory\[143\]\[0\] _05941_ _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07710__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14414_ _00268_ net3 mod.u_cpu.rf_ram.memory\[480\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13756__A1 _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11606__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11626_ _05208_ mod.u_cpu.rf_ram.memory\[262\]\[1\] _05223_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15394_ _01169_ net3 mod.u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14345_ _00199_ net3 mod.u_cpu.rf_ram.memory\[515\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11557_ _05179_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10508_ _04453_ mod.u_cpu.rf_ram.memory\[441\]\[0\] _04465_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14276_ _00130_ net3 mod.u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11488_ _05133_ _05131_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13227_ _03502_ _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10439_ _04418_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08113__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13158_ _06270_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15112__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12109_ _05555_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13089_ _02287_ _06227_ _06228_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07650_ _01827_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15262__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07581_ _01849_ _01871_ _01888_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09320_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09112__A1 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13995__A1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09251_ _03508_ _03510_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08202_ mod.u_cpu.rf_ram.memory\[565\]\[0\] _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09182_ _03462_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08133_ _02161_ mod.u_cpu.rf_ram.memory\[46\]\[0\] _02440_ _01828_ _02441_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07426__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__S1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ _02302_ mod.u_cpu.rf_ram.memory\[76\]\[0\] _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10981__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07285__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11585__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08966_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07862__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15605__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12486__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07917_ _01518_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08897_ _02471_ _03196_ _03203_ _02518_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09351__A1 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07848_ _01635_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12238__A1 _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07779_ mod.u_cpu.rf_ram.memory\[180\]\[0\] mod.u_cpu.rf_ram.memory\[181\]\[0\] mod.u_cpu.rf_ram.memory\[182\]\[0\]
+ mod.u_cpu.rf_ram.memory\[183\]\[0\] _02085_ _02086_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09789__I _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _01418_ _01498_ _01518_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10790_ _04654_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ _03675_ _03676_ _03677_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_169_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07760__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12460_ _05792_ _05796_ _05797_ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _05798_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _05080_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12391_ _03770_ _04142_ _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12410__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14136__S _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _04749_ _05011_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14130_ _07041_ mod.u_cpu.rf_ram.memory\[118\]\[1\] _07050_ _07052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15135__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14061_ _07006_ _07007_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11273_ _02398_ _04985_ _04986_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08917__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09029__I _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09965__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10224_ _04230_ _04269_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13910__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13012_ _03837_ _06080_ _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A2 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _04218_ _04202_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15285__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07772__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10086_ _04162_ mod.u_cpu.rf_ram.memory\[504\]\[0\] _04169_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14963_ _00817_ net3 mod.u_cpu.rf_ram.memory\[559\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13674__B1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13674__C2 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08089__B _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09342__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13914_ _06476_ _06892_ _06893_ _06894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14894_ _00748_ net3 mod.u_cpu.rf_ram.memory\[237\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12229__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13723__B _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13845_ _06775_ _06839_ _06450_ _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09699__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13776_ _06322_ _06714_ _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10988_ _04774_ mod.u_cpu.rf_ram.memory\[363\]\[0\] _04789_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15515_ _01286_ net3 mod.u_cpu.rf_ram.memory\[319\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12727_ _05963_ mod.u_cpu.rf_ram.memory\[78\]\[0\] _05975_ _05976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15446_ _01220_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12658_ _05923_ mod.u_cpu.rf_ram.memory\[145\]\[1\] _05928_ _05930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11609_ _05213_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12853__I _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15377_ _01152_ net3 mod.u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12589_ _05869_ mod.u_cpu.rf_ram.memory\[156\]\[0\] _05883_ _05884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14328_ _00182_ net3 mod.u_cpu.rf_ram.memory\[523\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11469__I _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08271__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14259_ _00113_ net3 mod.u_cpu.rf_ram.memory\[558\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14502__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08908__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15628__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13901__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08820_ _02411_ _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _01670_ _03057_ _02230_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14652__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11515__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07702_ _01581_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08682_ _02477_ _02987_ _02988_ _01638_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ _01938_ mod.u_cpu.rf_ram.memory\[310\]\[0\] _01940_ _01783_ _01941_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13968__A1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15008__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07564_ _01851_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09402__I _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09303_ _03495_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07495_ mod.u_cpu.rf_ram.memory\[445\]\[0\] _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07742__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09234_ _03405_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15158__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13196__A2 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09165_ _03451_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12243__I1 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ mod.u_cpu.rf_ram.memory\[56\]\[0\] mod.u_cpu.rf_ram.memory\[57\]\[0\] mod.u_cpu.rf_ram.memory\[58\]\[0\]
+ mod.u_cpu.rf_ram.memory\[59\]\[0\] _02242_ _02267_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12943__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08998__I1 _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09096_ mod.u_cpu.cpu.state.init_done _03391_ _03393_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_163_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ _02135_ mod.u_cpu.rf_ram.memory\[68\]\[0\] _02354_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09947__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09998_ _04107_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_107 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_118 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__12459__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_129 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08949_ mod.u_cpu.cpu.decode.opcode\[0\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11506__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__A1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13120__A2 _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11960_ _05457_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10911_ _04172_ _04713_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07886__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11682__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11891_ _05408_ _05401_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11842__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08637__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13630_ _06485_ _06284_ _06322_ _06305_ _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_10842_ _04689_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13561_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] mod.u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _06599_ _06600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12631__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _03895_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_158_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15300_ _00060_ net4 mod.u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10493__I0 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12512_ _05822_ mod.u_cpu.rf_ram.memory\[168\]\[1\] _05832_ _05834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13492_ _03624_ _06551_ _06552_ _03631_ _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_157_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15231_ _01084_ net3 mod.u_cpu.rf_ram.memory\[229\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12443_ _03498_ _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12673__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09468__B _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08372__B _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11198__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10245__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14525__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15162_ _01015_ net3 mod.u_cpu.rf_ram.memory\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12934__A2 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08063__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12374_ _05563_ _03866_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10193__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14113_ _06903_ _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07810__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ _05022_ _05021_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15093_ _00947_ net3 mod.u_cpu.rf_ram.memory\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14044_ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] _06989_ _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _04973_ _04969_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14675__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09563__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _04245_ mod.u_cpu.rf_ram.memory\[488\]\[1\] _04256_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11187_ _04784_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _04207_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09315__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10069_ _04157_ mod.u_cpu.rf_ram.memory\[507\]\[1\] _04155_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14946_ _00800_ net3 mod.u_cpu.rf_ram.memory\[220\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11122__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12465__A4 _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14877_ _00731_ net3 mod.u_cpu.rf_ram.memory\[253\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08547__B _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13828_ _06283_ _06824_ _06825_ _06642_ _06826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07629__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13759_ _06492_ _06712_ _06762_ _06475_ _06412_ _06763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__15300__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07280_ _01536_ _01571_ _01585_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15429_ _01204_ net3 mod.u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15450__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08054__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14127__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _04051_ mod.u_cpu.rf_ram.memory\[530\]\[0\] _04056_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13886__B1 _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09554__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10831__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _03999_ mod.u_cpu.rf_ram.memory\[541\]\[1\] _04007_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _02190_ _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09783_ _03956_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07345__C _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08109__A2 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08734_ _02197_ _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11113__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08665_ _02561_ _02968_ _02971_ _01696_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11662__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10711__I1 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _01634_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08596_ _01858_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09132__I mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10278__I _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07547_ _01854_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14548__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08293__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _01773_ _01777_ _01784_ _01785_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ mod.u_scanchain_local.module_data_in\[35\] mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _03479_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13413__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _03440_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14698__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _03379_ _03304_ _03380_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _04875_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12090_ _05542_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11041_ _04802_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10741__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_13 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10155__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__A3 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_24 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_35 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_46 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_57 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__07651__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_68 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__I1 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_79 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_14800_ _00654_ net3 mod.u_cpu.rf_ram.memory\[287\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12992_ _06163_ _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14731_ _00585_ net3 mod.u_cpu.rf_ram.memory\[322\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11943_ _05426_ mod.u_cpu.rf_ram.memory\[220\]\[1\] _05444_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07859__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15323__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14662_ _00516_ net3 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11874_ _05386_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13613_ _03378_ _06631_ _06632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _04666_ mod.u_cpu.rf_ram.memory\[38\]\[1\] _04676_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14593_ _00447_ net3 mod.u_cpu.rf_ram.memory\[391\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13801__B1 _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13544_ _06590_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15473__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12080__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10756_ _04622_ mod.u_cpu.rf_ram.memory\[400\]\[0\] _04631_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13499__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13475_ _06543_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10687_ _04586_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15214_ _01067_ net3 mod.u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12426_ _05770_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10918__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11966__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15145_ _00998_ net3 mod.u_cpu.rf_ram.memory\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12357_ _05711_ mod.u_cpu.rf_ram.memory\[122\]\[1\] _05722_ _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11308_ _05010_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15076_ _00930_ net3 mod.u_cpu.rf_ram.memory\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12288_ _05634_ _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14027_ mod.u_arbiter.i_wb_cpu_rdt\[19\] _06976_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11239_ _04961_ mod.u_cpu.rf_ram.memory\[324\]\[0\] _04962_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14929_ _00783_ net3 mod.u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08277__B _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08450_ _02742_ _02756_ _01483_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07401_ _01516_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08381_ _01879_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_195_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08114__I2 mod.u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09887__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07332_ mod.u_cpu.rf_ram.memory\[493\]\[0\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08275__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07263_ mod.u_cpu.rf_ram.memory\[464\]\[0\] mod.u_cpu.rf_ram.memory\[465\]\[0\] mod.u_cpu.rf_ram.memory\[466\]\[0\]
+ mod.u_cpu.rf_ram.memory\[467\]\[0\] _01567_ _01570_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14840__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09002_ _01430_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08027__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07194_ mod.u_cpu.rf_ram.memory\[448\]\[0\] mod.u_cpu.rf_ram.memory\[449\]\[0\] mod.u_cpu.rf_ram.memory\[450\]\[0\]
+ mod.u_cpu.rf_ram.memory\[451\]\[0\] _01496_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07200__I _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10385__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11582__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14990__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07250__A2 _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11709__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09904_ _02563_ _04042_ _04045_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14033__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09127__I mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12382__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09835_ _03991_ _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12689__S _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15346__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09766_ _03697_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13087__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08717_ mod.u_cpu.rf_ram.memory\[231\]\[1\] _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09697_ _03888_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14370__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10696__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08648_ mod.u_cpu.rf_ram.memory\[165\]\[1\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15496__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13821__B _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08579_ _01711_ _02885_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _04436_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08266__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11590_ _05201_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _04442_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13260_ _06357_ _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _04430_ mod.u_cpu.rf_ram.memory\[447\]\[1\] _04438_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12211_ _05624_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13191_ _05782_ _03456_ _06297_ _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_163_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12142_ _05575_ mod.u_cpu.rf_ram.memory\[75\]\[0\] _05577_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13268__B _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12073_ _05417_ _05388_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11325__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11024_ _04797_ mod.u_cpu.rf_ram.memory\[358\]\[1\] _04813_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11876__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14713__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12825__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12975_ _03389_ mod.u_cpu.cpu.state.o_cnt\[2\] _06150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14714_ _00568_ net3 mod.u_cpu.rf_ram.memory\[330\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _04994_ _05433_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14645_ _00499_ net3 mod.u_cpu.rf_ram.memory\[365\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14863__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11857_ _05383_ mod.u_cpu.rf_ram.memory\[6\]\[1\] _05381_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08257__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10808_ _04666_ mod.u_cpu.rf_ram.memory\[392\]\[1\] _04664_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14576_ _00430_ net3 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11788_ _05337_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__I _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__C _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13527_ _06578_ mod.u_cpu.rf_ram.memory\[129\]\[0\] _06579_ _06580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ _04619_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15219__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13458_ _03552_ _06531_ _06532_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _06533_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12409_ _05487_ _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12861__I _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10582__S _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13389_ _06377_ _03449_ _06484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11564__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15128_ _00981_ net3 mod.u_cpu.rf_ram.memory\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14243__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15369__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11477__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13893__S _06882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10381__I _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ mod.u_cpu.rf_ram.memory\[245\]\[0\] _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15059_ _00913_ net3 mod.u_cpu.rf_ram.memory\[190\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11316__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07881_ mod.u_cpu.rf_ram.memory\[222\]\[0\] mod.u_cpu.rf_ram.memory\[223\]\[0\] _02048_
+ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09620_ _03827_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14393__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13069__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07690__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__C _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09551_ _03695_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07623__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08502_ mod.u_cpu.rf_ram.memory\[325\]\[1\] _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12101__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09482_ _01659_ _03703_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08433_ _02654_ _02736_ _02739_ _02730_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12419__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _02638_ mod.u_cpu.rf_ram.memory\[484\]\[1\] _02670_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12044__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13241__A1 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10055__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _01573_ _01622_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09996__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__A2 _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10556__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08295_ mod.u_cpu.rf_ram.memory\[455\]\[1\] _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _01489_ _01535_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _01484_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12355__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14736__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09818_ mod.u_cpu.rf_ram.memory\[545\]\[1\] _03929_ _03981_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09920__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12212__S _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09749_ mod.u_cpu.rf_ram.memory\[553\]\[1\] _03929_ _03926_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12807__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13855__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14886__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12760_ _05992_ mod.u_cpu.rf_ram.memory\[135\]\[0\] _05996_ _05997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08487__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07534__I0 mod.u_cpu.rf_ram.memory\[320\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I1 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _03803_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12691_ _03723_ _05319_ _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08645__B _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14430_ _00284_ net3 mod.u_cpu.rf_ram.memory\[472\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11642_ _05110_ _04026_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14361_ _00215_ net3 mod.u_cpu.rf_ram.memory\[507\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13783__A2 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10466__I _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _05178_ mod.u_cpu.rf_ram.memory\[271\]\[1\] _05188_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13312_ _06401_ _06408_ _06409_ _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12991__B1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10524_ _04180_ _04464_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14292_ _00146_ net3 mod.u_cpu.rf_ram.memory\[541\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14266__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15511__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13243_ _06346_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10455_ _04428_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07775__I _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11546__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13174_ mod.u_arbiter.i_wb_cpu_rdt\[10\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _05781_ _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07214__A2 _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10386_ _03928_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07845__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12125_ _05549_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12056_ _05309_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11961__S _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13017__I _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08478__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12958_ _06134_ _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ _04300_ _05371_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12889_ _06082_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14628_ _00482_ net3 mod.u_cpu.rf_ram.memory\[373\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15041__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09230__I mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10037__A1 _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14609__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11085__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14559_ _00413_ net3 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08080_ _02126_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08650__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15191__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13526__A2 _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07685__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12585__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14759__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08982_ mod.u_cpu.cpu.decode.co_mem_word mod.u_cpu.cpu.csr_d_sel _03287_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10760__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ _02170_ _02233_ _02240_ _02168_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12032__S _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07864_ _01614_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09603_ _03814_ _03805_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07795_ _02089_ _02101_ _02102_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09534_ _03757_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08469__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09130__A2 _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09465_ _03292_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07141__A1 _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08416_ mod.u_cpu.rf_ram.memory\[408\]\[1\] mod.u_cpu.rf_ram.memory\[409\]\[1\] mod.u_cpu.rf_ram.memory\[410\]\[1\]
+ mod.u_cpu.rf_ram.memory\[411\]\[1\] _02225_ _02325_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12017__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09396_ _03631_ _03627_ _03493_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14289__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15534__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _02218_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10823__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08278_ _01636_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08641__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08492__I1 mod.u_cpu.rf_ram.memory\[329\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ _01515_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11528__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11111__S _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ _04280_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10051__I1 mod.u_cpu.rf_ram.memory\[510\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ mod.u_cpu.rf_ram.memory\[493\]\[1\] _04111_ _04229_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__S _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12450__B _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13930_ _06905_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11700__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13861_ _06853_ _06854_ _06855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15600_ _01371_ net3 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _04844_ _06030_ _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08004__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15064__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13792_ _06425_ _06373_ _06402_ _06683_ _06793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_28_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12500__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15531_ _01302_ net3 mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12743_ _03790_ _05552_ _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07132__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15462_ _01236_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12674_ _04913_ _05940_ _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09050__I _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14413_ _00267_ net3 mod.u_cpu.rf_ram.memory\[481\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08094__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11625_ _05224_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15393_ _01168_ net3 mod.u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11767__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14344_ _00198_ net3 mod.u_cpu.rf_ram.memory\[515\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11556_ _05178_ mod.u_cpu.rf_ram.memory\[274\]\[1\] _05175_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14901__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _04163_ _04464_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13508__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14275_ _00129_ net3 mod.u_cpu.rf_ram.memory\[550\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10924__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11487_ _05132_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13226_ _06139_ _06332_ _06333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_171_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _04400_ mod.u_cpu.rf_ram.memory\[452\]\[0\] _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12192__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13157_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _06268_ _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10369_ _04311_ _04370_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12108_ _05550_ mod.u_cpu.rf_ram.memory\[211\]\[1\] _05553_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13088_ _06032_ _06227_ _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12039_ _05443_ _03810_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08699__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15407__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07580_ _01872_ _01873_ _01885_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13444__B2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09112__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14431__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13995__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15557__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _01682_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09181_ mod.u_arbiter.i_wb_cpu_rdt\[17\] mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _03459_
+ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11758__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _01819_ _02439_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10805__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14581__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08063_ _02369_ _02370_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08304__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07729__A3 _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07285__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08965_ _03269_ mod.u_cpu.cpu.state.o_cnt\[2\] _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14041__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07916_ _01651_ _02223_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15087__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ _02476_ _03199_ _03202_ _02489_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12486__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _02154_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08974__I mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07752__I3 mod.u_cpu.rf_ram.memory\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07778_ _01854_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08907__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09517_ _01461_ _01778_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08537__S1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07811__C _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__A1 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11997__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _03334_ _03668_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14924__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _03602_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03586_ _03594_ _03618_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_178_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11410_ mod.u_cpu.rf_ram.memory\[297\]\[0\] _04954_ _05079_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12797__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12390_ _05746_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12410__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11341_ _05033_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14060_ mod.u_arbiter.i_wb_cpu_rdt\[28\] _06998_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14163__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11272_ _04746_ _04985_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07258__C _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13371__B1 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13011_ _06177_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08917__A2 _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10223_ _04108_ _04228_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14304__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _03885_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11575__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14962_ _00816_ net3 mod.u_cpu.rf_ram.memory\[559\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10085_ _04168_ _04164_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13674__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13674__B2 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13913_ _06398_ _06452_ _06695_ _06893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14454__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14893_ _00747_ net3 mod.u_cpu.rf_ram.memory\[239\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13844_ _06367_ _06743_ _06839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12229__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13775_ _06776_ _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10987_ _04238_ _04788_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11988__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11016__S _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15514_ _01285_ net3 mod.u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12726_ _03885_ _05576_ _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08853__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15445_ _01219_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12657_ _05929_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11608_ mod.u_cpu.rf_ram.memory\[265\]\[1\] _05065_ _05211_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08605__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15376_ _01151_ net3 mod.u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09653__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12588_ _05443_ _05882_ _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14327_ _00181_ net3 mod.u_cpu.rf_ram.memory\[524\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11460__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _05167_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14258_ _00112_ net3 mod.u_cpu.rf_ram.memory\[558\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13209_ _06117_ _06300_ _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08908__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13901__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14189_ _07090_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11912__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ mod.u_cpu.rf_ram.memory\[104\]\[1\] mod.u_cpu.rf_ram.memory\[105\]\[1\] mod.u_cpu.rf_ram.memory\[106\]\[1\]
+ mod.u_cpu.rf_ram.memory\[107\]\[1\] _02106_ _02107_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08216__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13665__A1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07701_ _01978_ _01990_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08681_ _02632_ mod.u_cpu.rf_ram.memory\[208\]\[1\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07344__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07632_ _01507_ _01939_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13417__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14947__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13968__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _01852_ _01853_ _01869_ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14090__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ _03552_ _03549_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08844__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07647__A2 _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07494_ _01752_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__07203__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09233_ _03491_ _03494_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13141__S _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__B _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12779__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09164_ _03413_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08115_ mod.u_cpu.rf_ram.memory\[60\]\[0\] mod.u_cpu.rf_ram.memory\[61\]\[0\] mod.u_cpu.rf_ram.memory\[62\]\[0\]
+ mod.u_cpu.rf_ram.memory\[63\]\[0\] _02369_ _02218_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14036__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ _03394_ _03395_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14327__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08046_ _02266_ _02353_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11596__S _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10006__I1 mod.u_cpu.rf_ram.memory\[516\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09947__I1 mod.u_cpu.rf_ram.memory\[526\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09021__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14477__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09997_ _04106_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_108 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08948_ _01422_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13656__A1 _06312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12459__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_119 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ _03176_ _03185_ _02609_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08918__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10910_ _04736_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11890_ _03973_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10890__A1 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _04679_ mod.u_cpu.rf_ram.memory\[386\]\[0\] _04688_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13560_ _06583_ _06599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_125_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _04642_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09883__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12631__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12511_ _05833_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15102__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11690__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13491_ _06553_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_157_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15230_ _01083_ net3 mod.u_cpu.rf_ram.memory\[229\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12442_ _01433_ _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09635__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08438__I1 mod.u_cpu.rf_ram.memory\[389\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08372__C _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10474__I _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15161_ _01014_ net3 mod.u_cpu.rf_ram.memory\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12373_ _05735_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12934__A3 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15252__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14112_ _07040_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__I1 mod.u_cpu.rf_ram.memory\[569\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11324_ _04541_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15092_ _00946_ net3 mod.u_cpu.rf_ram.memory\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14043_ _06992_ _06994_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _04125_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10206_ _04257_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09563__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11186_ _04905_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10137_ _04193_ mod.u_cpu.rf_ram.memory\[497\]\[0\] _04206_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09315__A2 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _04090_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14945_ _00799_ net3 mod.u_cpu.rf_ram.memory\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12170__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14876_ _00730_ net3 mod.u_cpu.rf_ram.memory\[253\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10881__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13827_ _06319_ _06324_ _06643_ _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10649__I _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14072__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13758_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_arbiter.i_wb_cpu_rdt\[3\] _03509_
+ _06762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08826__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__A2 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12709_ _05870_ _04668_ _05964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13689_ _06695_ _06698_ _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15428_ _01203_ net3 mod.u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09626__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__C _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15359_ _01134_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13695__I _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09920_ _03859_ _04038_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13886__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09851_ _02573_ _04007_ _04008_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08802_ mod.u_cpu.rf_ram.memory\[71\]\[1\] _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12104__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09782_ _03916_ mod.u_cpu.rf_ram.memory\[54\]\[0\] _03955_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ mod.u_cpu.rf_ram.memory\[253\]\[1\] _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12161__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08664_ _02566_ mod.u_cpu.rf_ram.memory\[222\]\[1\] _02970_ _01703_ _02971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07615_ _01643_ mod.u_cpu.rf_ram.memory\[316\]\[0\] _01922_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15125__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14063__A1 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08595_ mod.u_cpu.rf_ram.memory\[261\]\[1\] _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__I0 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ _01499_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08029__I _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08817__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _01765_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09490__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15275__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _03481_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09617__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13413__I1 mod.u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _03438_ _03439_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09078_ mod.u_cpu.cpu.alu.add_cy_r _03356_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13177__I0 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _02057_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13877__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11040_ _04826_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_14 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_25 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_36 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_47 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_58 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07651__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_69 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12991_ _06062_ _03375_ _03337_ _03336_ _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07308__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11942_ _05445_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14730_ _00584_ net3 mod.u_cpu.rf_ram.memory\[322\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__A2 _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10469__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14661_ _00515_ net3 mod.u_cpu.rf_ram.memory\[357\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10863__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11873_ _03940_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13612_ _06624_ _06628_ _06629_ _06630_ _06631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10824_ _04677_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15618__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14592_ _00446_ net3 mod.u_cpu.rf_ram.memory\[391\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08808__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13543_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] mod.u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _06589_ _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10755_ _04209_ _04623_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08383__B _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13474_ _03588_ _06538_ _06540_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _06543_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10686_ _04584_ mod.u_cpu.rf_ram.memory\[412\]\[0\] _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15213_ _01066_ net3 mod.u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12425_ _05761_ mod.u_cpu.rf_ram.memory\[174\]\[1\] _05768_ _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14642__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11415__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15144_ _00997_ net3 mod.u_cpu.rf_ram.memory\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12356_ _05723_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13317__B1 _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13168__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__A1 _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11307_ _04999_ mod.u_cpu.rf_ram.memory\[314\]\[1\] _05008_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08830__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15075_ _00929_ net3 mod.u_cpu.rf_ram.memory\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12287_ _05676_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14792__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14026_ _06970_ _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11238_ _04821_ _04945_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__S _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11169_ _04901_ mod.u_cpu.rf_ram.memory\[335\]\[0\] _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15148__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11763__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14928_ _00782_ net3 mod.u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10379__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14045__A1 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14859_ _00713_ net3 mod.u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14045__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _01705_ mod.u_cpu.rf_ram.memory\[412\]\[0\] _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15298__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08380_ _02591_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09847__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07331_ mod.u_cpu.rf_ram.memory\[488\]\[0\] mod.u_cpu.rf_ram.memory\[489\]\[0\] mod.u_cpu.rf_ram.memory\[490\]\[0\]
+ mod.u_cpu.rf_ram.memory\[491\]\[0\] _01636_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08114__I3 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12594__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09001_ _03299_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11406__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ _01500_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08027__A2 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13159__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11938__I _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08740__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12035__S _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13859__B2 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12906__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _04044_ _04042_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12531__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09765_ _03834_ _03942_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08716_ _01608_ mod.u_cpu.rf_ram.memory\[228\]\[1\] _03022_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10145__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09696_ _03877_ mod.u_cpu.rf_ram.memory\[558\]\[0\] _03887_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14515__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ mod.u_cpu.rf_ram.memory\[160\]\[1\] mod.u_cpu.rf_ram.memory\[161\]\[1\] mod.u_cpu.rf_ram.memory\[162\]\[1\]
+ mod.u_cpu.rf_ram.memory\[163\]\[1\] _02125_ _02127_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10845__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08578_ mod.u_cpu.rf_ram.memory\[285\]\[1\] _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08915__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14665__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07529_ _01510_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11645__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _04452_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _01808_ _04438_ _04440_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12210_ mod.u_cpu.rf_ram.memory\[1\]\[0\] _05622_ _05623_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13190_ _06116_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _06297_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_191_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12141_ _04930_ _05576_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09518__A2 _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12072_ _05530_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11325__A2 _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11023_ _04814_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13570__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__B _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12974_ _06149_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15440__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14713_ _00567_ net3 mod.u_cpu.rf_ram.memory\[331\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14027__A1 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11925_ _05432_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07701__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14644_ _00498_ net3 mod.u_cpu.rf_ram.memory\[365\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11856_ _05328_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _04640_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14575_ _00429_ net3 mod.u_cpu.rf_ram.memory\[400\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08257__A2 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15590__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11787_ _05311_ mod.u_cpu.rf_ram.memory\[234\]\[0\] _05336_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13303__I _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ _04608_ mod.u_cpu.rf_ram.memory\[403\]\[1\] _04617_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13526_ _03980_ _05373_ _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11959__S _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13457_ _06513_ _06532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10669_ _04573_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12408_ _05187_ _05757_ _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12061__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13388_ _06482_ _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07768__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15127_ _00980_ net3 mod.u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12339_ _05711_ mod.u_cpu.rf_ram.memory\[183\]\[1\] _05707_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15058_ _00912_ net3 mod.u_cpu.rf_ram.memory\[190\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08980__A3 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13973__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14009_ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] _06966_ _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13561__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07880_ _01582_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10375__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14538__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13069__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07940__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__I1 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _03767_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10127__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08501_ mod.u_cpu.rf_ram.memory\[320\]\[1\] mod.u_cpu.rf_ram.memory\[321\]\[1\] mod.u_cpu.rf_ram.memory\[322\]\[1\]
+ mod.u_cpu.rf_ram.memory\[323\]\[1\] _01920_ _02666_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09481_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _01441_ _03706_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14688__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _02692_ mod.u_cpu.rf_ram.memory\[406\]\[1\] _02738_ _01918_ _02739_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07920__B _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _01561_ _02669_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07314_ mod.u_cpu.rf_ram.memory\[485\]\[0\] _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10055__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _02585_ mod.u_cpu.rf_ram.memory\[452\]\[1\] _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _01536_ _01541_ _01549_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__B _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _01450_ _01456_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11668__I _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__C _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08042__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12355__I1 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08184__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15463__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _03982_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07931__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11109__S _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12807__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13855__I1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13832__B _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11866__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14009__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ _03847_ mod.u_cpu.rf_ram.memory\[560\]\[0\] _03874_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A2 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11710_ _05282_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12690_ _05951_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12448__B _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11641_ _05235_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09436__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14360_ _00214_ net3 mod.u_cpu.rf_ram.memory\[507\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08217__I _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11572_ _02028_ _05188_ _05189_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07121__I mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13311_ _06134_ _06409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10523_ _04475_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14291_ _00145_ net3 mod.u_cpu.rf_ram.memory\[542\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13242_ _06273_ mod.u_cpu.rf_ram.memory\[93\]\[0\] _06345_ _06346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10454_ _04423_ mod.u_cpu.rf_ram.memory\[44\]\[0\] _04427_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12743__A1 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07277__B _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13173_ mod.u_cpu.cpu.bufreg.i_sh_signed _06140_ _06280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10385_ _01542_ _04381_ _04382_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08411__A2 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07845__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _05565_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12055_ _05519_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11006_ _04620_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09372__B1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14830__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12957_ _06064_ _06133_ _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08478__A2 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11908_ _05420_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14980__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12888_ _06073_ mod.u_cpu.rf_ram.memory\[89\]\[0\] _06081_ _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13759__B1 _06762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14627_ _00481_ net3 mod.u_cpu.rf_ram.memory\[374\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11839_ _03662_ _04223_ _03753_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11085__I1 mod.u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14558_ _00412_ net3 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15336__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13509_ _06562_ _03302_ _03260_ _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14489_ _00343_ net3 mod.u_cpu.rf_ram.memory\[443\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09159__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10392__I _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08402__A2 _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14360__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15486__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13917__B _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ _01428_ _01429_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13534__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07932_ _02155_ _02236_ _02239_ _02166_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07863_ _01806_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09602_ _03757_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07794_ _02057_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09533_ _03756_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13998__B1 _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09464_ _03685_ _03690_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10520__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07141__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08415_ _01459_ _02701_ _02721_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09395_ _03631_ _03624_ _03620_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__09418__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08346_ _01592_ _02643_ _02652_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11599__S _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12973__A1 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12782__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08277_ _01466_ _02038_ _02448_ _02584_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__12973__B2 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07228_ _01492_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14703__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__A2 _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _01463_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _01467_ mod.u_cpu.cpu.immdec.imm24_20\[4\]
+ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10587__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10170_ _01640_ _04229_ _04231_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14853__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11700__A2 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12022__I _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13860_ _06465_ _06744_ _06840_ _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15209__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _05630_ _06030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13791_ _06791_ _06714_ _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08004__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11861__I _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15530_ _01301_ net3 mod.u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12742_ _05985_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14233__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15359__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12673_ _05919_ _05940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15461_ _01235_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09409__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14412_ _00266_ net3 mod.u_cpu.rf_ram.memory\[481\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11216__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11624_ _05222_ mod.u_cpu.rf_ram.memory\[262\]\[0\] _05223_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12264__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15392_ _01167_ net3 mod.u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12964__A1 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11767__A2 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__A4 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14343_ _00197_ net3 mod.u_cpu.rf_ram.memory\[516\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11555_ _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08391__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14383__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10506_ _04442_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14274_ _00128_ net3 mod.u_cpu.rf_ram.memory\[550\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11486_ _03773_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13225_ _06331_ _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _04272_ _04407_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11101__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13156_ _06269_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10368_ _04369_ _04335_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__I3 mod.u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12107_ _02210_ _05553_ _05554_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13087_ _03941_ _06030_ _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10299_ _04322_ _04303_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12038_ _05508_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11972__S _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13989_ _06942_ _06954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11771__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10502__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08320__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ mod.u_cpu.rf_ram.memory\[560\]\[0\] mod.u_cpu.rf_ram.memory\[561\]\[0\] mod.u_cpu.rf_ram.memory\[562\]\[0\]
+ mod.u_cpu.rf_ram.memory\[563\]\[0\] _02507_ _02473_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09180_ _03461_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14726__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12255__I0 _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ mod.u_cpu.rf_ram.memory\[47\]\[0\] _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11758__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08062_ mod.u_cpu.rf_ram.memory\[77\]\[0\] _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14876__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08387__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13380__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13139__S _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11946__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10850__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ mod.u_cpu.cpu.mem_bytecnt\[0\] _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08139__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14180__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07915_ _02066_ mod.u_cpu.rf_ram.memory\[214\]\[0\] _02222_ _01821_ _02223_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08895_ _02483_ mod.u_cpu.rf_ram.memory\[566\]\[1\] _03201_ _02487_ _03202_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13683__A2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07846_ _01749_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14256__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07777_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11681__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15501__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _03739_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08311__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__A2 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08195__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11997__A2 _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09447_ _03323_ _03324_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09378_ _03610_ _03608_ _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08329_ _02421_ _02635_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11340_ _05032_ mod.u_cpu.rf_ram.memory\[30\]\[1\] _05029_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _04983_ _04984_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13010_ _06105_ mod.u_cpu.rf_ram.memory\[86\]\[1\] _06175_ _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10222_ _04268_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13371__A1 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11856__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10153_ _04147_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15031__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07440__I3 mod.u_cpu.rf_ram.memory\[419\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14961_ _00815_ net3 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10084_ _03804_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13674__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13912_ _06471_ _06823_ _06390_ _06660_ _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_43_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09342__A3 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14892_ _00746_ net3 mod.u_cpu.rf_ram.memory\[239\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08550__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13843_ _06677_ _06838_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15181__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11437__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14749__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13774_ _06289_ _06775_ _06643_ _06317_ _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_10986_ _04703_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09061__I mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__S0 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15513_ _01284_ net3 mod.u_cpu.rf_ram.memory\[329\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12725_ _05974_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15444_ _01218_ net3 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12656_ _05918_ mod.u_cpu.rf_ram.memory\[145\]\[0\] _05928_ _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14899__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12937__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10935__I _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11607_ _05212_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12587_ _05373_ _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15375_ _01150_ net3 mod.u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13311__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14326_ _00180_ net3 mod.u_cpu.rf_ram.memory\[524\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _05162_ mod.u_cpu.rf_ram.memory\[277\]\[1\] _05165_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14257_ _00111_ net3 mod.u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10871__S _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ _05118_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08369__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13208_ _06311_ _06314_ _06315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14188_ _03699_ mod.u_cpu.rf_ram.memory\[244\]\[0\] _07089_ _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11766__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11912__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10670__I _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13139_ mod.u_arbiter.i_wb_cpu_rdt\[21\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _06258_ _06260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10971__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14279__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08216__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13665__A2 _06659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15524__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ _01992_ _01996_ _02006_ _02007_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08680_ mod.u_cpu.rf_ram.memory\[209\]\[1\] _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07631_ mod.u_cpu.rf_ram.memory\[311\]\[0\] _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13417__A2 _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07562_ _01550_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07493_ mod.u_cpu.rf_ram.memory\[440\]\[0\] mod.u_cpu.rf_ram.memory\[441\]\[0\] mod.u_cpu.rf_ram.memory\[442\]\[0\]
+ mod.u_cpu.rf_ram.memory\[443\]\[0\] _01753_ _01771_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11006__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _03492_ _03493_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08743__C _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12928__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09163_ _03450_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08114_ mod.u_cpu.rf_ram.memory\[48\]\[0\] mod.u_cpu.rf_ram.memory\[49\]\[0\] mod.u_cpu.rf_ram.memory\[50\]\[0\]
+ mod.u_cpu.rf_ram.memory\[51\]\[0\] _02421_ _02350_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _03349_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ mod.u_cpu.rf_ram.memory\[69\]\[0\] _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15054__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10167__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ _03702_ _03939_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09146__I _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13105__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08780__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_109 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08947_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12703__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11667__A1 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08878_ _02592_ _03177_ _03184_ _01836_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_151_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__A1 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07829_ mod.u_cpu.rf_ram.memory\[167\]\[0\] _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11419__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _04281_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13813__C1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10890__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12092__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10771_ _04641_ mod.u_cpu.rf_ram.memory\[398\]\[1\] _04638_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07194__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12510_ _05827_ mod.u_cpu.rf_ram.memory\[168\]\[0\] _05832_ _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13490_ _03616_ _06551_ _06552_ _03624_ _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_185_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12441_ _05779_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08653__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08225__I _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12372_ _05729_ mod.u_cpu.rf_ram.memory\[499\]\[1\] _05733_ _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15160_ _01013_ net3 mod.u_cpu.rf_ram.memory\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14111_ _07021_ mod.u_cpu.rf_ram.memory\[87\]\[0\] _07039_ _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11323_ _05019_ _05020_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15091_ _00945_ net3 mod.u_cpu.rf_ram.memory\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12970__I _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14042_ mod.u_arbiter.i_wb_cpu_rdt\[23\] _06987_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11254_ _04972_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14421__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10205_ _04249_ mod.u_cpu.rf_ram.memory\[488\]\[0\] _04256_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15547__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11185_ _04925_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _03866_ _04202_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10067_ _04156_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14944_ _00798_ net3 mod.u_cpu.rf_ram.memory\[169\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14571__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14875_ _00729_ net3 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13826_ _06471_ _06823_ _06695_ _06490_ _06824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_63_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10881__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14072__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13757_ _06492_ _06319_ _06713_ _06744_ _06365_ _06761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10866__S _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10969_ _04774_ mod.u_cpu.rf_ram.memory\[366\]\[0\] _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08382__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12708_ _05962_ _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13688_ _06494_ _06644_ _06696_ _06697_ _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__08563__C _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15427_ _01202_ net3 mod.u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12639_ _05907_ mod.u_cpu.rf_ram.memory\[148\]\[1\] _05915_ _05917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09626__I1 mod.u_cpu.rf_ram.memory\[566\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15077__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15358_ _01133_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10397__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09251__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14309_ _00163_ net3 mod.u_cpu.rf_ram.memory\[533\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14073__S _07015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15289_ _00048_ net4 mod.u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10149__A1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13886__A2 _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _03945_ _04007_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14914__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08801_ _02204_ mod.u_cpu.rf_ram.memory\[68\]\[1\] _03107_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _03878_ _03829_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13638__A2 _06648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08732_ mod.u_cpu.rf_ram.memory\[248\]\[1\] mod.u_cpu.rf_ram.memory\[249\]\[1\] mod.u_cpu.rf_ram.memory\[250\]\[1\]
+ mod.u_cpu.rf_ram.memory\[251\]\[1\] _03001_ _01525_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_61_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ _02711_ _02969_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08738__C _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13216__I _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _01920_ _01921_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08594_ mod.u_cpu.rf_ram.memory\[256\]\[1\] mod.u_cpu.rf_ram.memory\[257\]\[1\] mod.u_cpu.rf_ram.memory\[258\]\[1\]
+ mod.u_cpu.rf_ram.memory\[259\]\[1\] _01837_ _02252_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08117__I1 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07545_ mod.u_cpu.rf_ram.memory\[376\]\[0\] mod.u_cpu.rf_ram.memory\[377\]\[0\] mod.u_cpu.rf_ram.memory\[378\]\[0\]
+ mod.u_cpu.rf_ram.memory\[379\]\[0\] _01837_ _01838_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13810__A2 _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07476_ _01689_ mod.u_cpu.rf_ram.memory\[430\]\[0\] _01781_ _01783_ _01784_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11821__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09215_ mod.u_scanchain_local.module_data_in\[34\] mod.u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _03479_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _03405_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12621__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14444__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09077_ mod.u_cpu.cpu.alu.add_cy_r _03308_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12129__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _02104_ _02311_ _02335_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14594__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_15 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_26 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13835__B _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_37 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09979_ _04095_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10560__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_48 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_59 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12990_ _05780_ _06161_ _03373_ _06162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07308__A2 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11941_ _05442_ mod.u_cpu.rf_ram.memory\[220\]\[0\] _05444_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10312__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13126__I _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14660_ _00514_ net3 mod.u_cpu.rf_ram.memory\[357\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10863__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11872_ _05394_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13611_ mod.u_cpu.cpu.alu.cmp_r _03687_ _03305_ _06624_ _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10823_ _04663_ mod.u_cpu.rf_ram.memory\[38\]\[0\] _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14591_ _00445_ net3 mod.u_cpu.rf_ram.memory\[392\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08808__A2 _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13801__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13542_ _06583_ _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10754_ _04630_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__A1 _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10685_ _04315_ _04575_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13473_ _06542_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08116__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15212_ _01065_ net3 mod.u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12424_ _05769_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15143_ _00996_ net3 mod.u_cpu.rf_ram.memory\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12355_ _05713_ mod.u_cpu.rf_ram.memory\[122\]\[0\] _05722_ _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07794__I _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13317__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14937__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11306_ _05009_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12286_ _05662_ mod.u_cpu.rf_ram.memory\[18\]\[0\] _05675_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15074_ _00928_ net3 mod.u_cpu.rf_ram.memory\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14025_ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] _06978_ _06981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11237_ _04960_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08744__A1 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11168_ _04913_ _04906_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10119_ _04147_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11099_ _04867_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09514__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14927_ _00781_ net3 mod.u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14317__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14858_ _00712_ net3 mod.u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14045__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13809_ _06401_ _06808_ _06809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14789_ _00643_ net3 mod.u_cpu.rf_ram.memory\[293\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08355__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07330_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11803__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14467__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07261_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ mod.u_cpu.cpu.alu.add_cy_r mod.u_cpu.cpu.alu.i_rs1 _03304_ _03305_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_164_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12603__I0 _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07192_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07235__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09902_ _04043_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12115__I _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07209__I _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08735__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14108__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12531__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ _03994_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10542__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08468__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08715_ _02027_ _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09695_ _03855_ _03886_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08594__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08646_ _01670_ _02945_ _02952_ _02122_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15242__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10845__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08577_ mod.u_cpu.rf_ram.memory\[280\]\[1\] mod.u_cpu.rf_ram.memory\[281\]\[1\] mod.u_cpu.rf_ram.memory\[282\]\[1\]
+ mod.u_cpu.rf_ram.memory\[283\]\[1\] _02020_ _01995_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _01677_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12842__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09463__A2 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15392__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07459_ _01751_ _01756_ _01764_ _01766_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_167_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _04439_ _04438_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ _03392_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12140_ _05387_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10781__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ _05518_ mod.u_cpu.rf_ram.memory\[63\]\[1\] _05528_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07119__I mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ _04803_ mod.u_cpu.rf_ram.memory\[358\]\[0\] _04813_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08726__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08378__C _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12973_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie _06145_ _06148_ _03353_ _06149_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14712_ _00566_ net3 mod.u_cpu.rf_ram.memory\[331\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _05421_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14643_ _00497_ net3 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11855_ _05382_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08394__B _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07789__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08337__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _04665_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12833__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14574_ _00428_ net3 mod.u_cpu.rf_ram.memory\[400\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11786_ _05334_ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13525_ _06577_ _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _04618_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13456_ _06510_ _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10668_ _04560_ mod.u_cpu.rf_ram.memory\[415\]\[1\] _04571_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12407_ _05725_ _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10943__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13387_ _06064_ _06482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10599_ _04514_ mod.u_cpu.rf_ram.memory\[426\]\[1\] _04524_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10072__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07768__A2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15126_ _00979_ net3 mod.u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12338_ _05710_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15115__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13010__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15057_ _00911_ net3 mod.u_cpu.rf_ram.memory\[191\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12269_ _05664_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__A4 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14008_ _06967_ _06968_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13710__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15265__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07940__A2 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10127__I1 mod.u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08500_ _02778_ _02799_ _02806_ _01870_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09480_ _01461_ _03705_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12029__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ _02244_ _02737_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__C _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07699__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ mod.u_cpu.rf_ram.memory\[485\]\[1\] _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09445__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07313_ mod.u_cpu.rf_ram.memory\[480\]\[0\] mod.u_cpu.rf_ram.memory\[481\]\[0\] mod.u_cpu.rf_ram.memory\[482\]\[0\]
+ mod.u_cpu.rf_ram.memory\[483\]\[0\] _01605_ _01570_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07456__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08293_ _01607_ _02599_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11014__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11949__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _01482_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10063__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08708__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15608__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08184__A2 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09816_ mod.u_cpu.rf_ram.memory\[545\]\[0\] _03925_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08198__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _03733_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14632__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09133__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09678_ _03855_ _03873_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11866__I1 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08926__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08629_ mod.u_cpu.rf_ram.memory\[180\]\[1\] mod.u_cpu.rf_ram.memory\[181\]\[1\] mod.u_cpu.rf_ram.memory\[182\]\[1\]
+ mod.u_cpu.rf_ram.memory\[183\]\[1\] _02085_ _02086_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07695__A1 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13768__A1 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13768__B2 _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14782__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11640_ _05234_ mod.u_cpu.rf_ram.memory\[260\]\[1\] _05232_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09436__A2 _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__A1 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _05133_ _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_168_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ _06403_ _06407_ _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10522_ _04467_ mod.u_cpu.rf_ram.memory\[43\]\[1\] _04473_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14290_ _00144_ net3 mod.u_cpu.rf_ram.memory\[542\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12464__B _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15138__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11859__I _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10453_ _04251_ _03905_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13241_ _03771_ _06344_ _06345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10384_ _04230_ _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13172_ _06047_ _06279_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12123_ _05559_ mod.u_cpu.rf_ram.memory\[20\]\[0\] _05564_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15288__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12054_ _05518_ mod.u_cpu.rf_ram.memory\[61\]\[1\] _05516_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _04801_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09124__A1 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13742__C _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12956_ _06121_ _06130_ _06132_ _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09675__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11907_ _05406_ mod.u_cpu.rf_ram.memory\[224\]\[1\] _05418_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12887_ _05896_ _06080_ _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13759__A1 _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14626_ _00480_ net3 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13759__B2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11838_ _05370_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14557_ _00411_ net3 mod.u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11769_ mod.u_cpu.rf_ram.memory\[237\]\[1\] _05230_ _05321_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ mod.u_cpu.cpu.ctrl.i_jump _03325_ _06563_ _06564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14488_ _00342_ net3 mod.u_cpu.rf_ram.memory\[443\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10993__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13439_ _06521_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13189__C _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09239__I _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14505__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08143__I _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15109_ _00963_ net3 mod.u_cpu.rf_ram.memory\[173\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08980_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _03284_ mod.u_cpu.cpu.genblk3.csr.o_new_irq
+ _01422_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_170_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07931_ _02179_ mod.u_cpu.rf_ram.memory\[230\]\[0\] _02238_ _02164_ _02239_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__C _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14655__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _01741_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _03813_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13933__B _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07793_ _01836_ _02095_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13998__A1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09532_ _03753_ _03755_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09702__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09666__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09463_ _03252_ _03276_ _03689_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11473__A2 _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10520__I1 mod.u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ _02609_ _02710_ _02720_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09394_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09418__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07429__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _02631_ _02644_ _02651_ _02377_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12422__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ _01464_ _01465_ _02522_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_165_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07227_ _01493_ _01502_ _01530_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13922__A1 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ _01449_ _01465_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__15430__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10587__I1 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15580__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08937__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12810_ _06029_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13790_ _06291_ _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09657__A2 _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12459__B _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09612__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12741_ _05984_ mod.u_cpu.rf_ram.memory\[209\]\[1\] _05982_ _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07668__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07560__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15460_ _01234_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12672_ _05939_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14411_ _00265_ net3 mod.u_cpu.rf_ram.memory\[482\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11623_ _04812_ _05214_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15391_ _01166_ net3 mod.u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11216__A2 _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10275__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14528__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14342_ _00196_ net3 mod.u_cpu.rf_ram.memory\[516\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12964__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11554_ _05106_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10975__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08391__C _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _04463_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14273_ _00127_ net3 mod.u_cpu.rf_ram.memory\[551\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11485_ _04994_ _05130_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13224_ _06323_ _06326_ _06330_ _06331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13913__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10436_ _04416_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14678__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13155_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _06268_ _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _04066_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12106_ _05488_ _05553_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13086_ _06226_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10298_ _03796_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12037_ mod.u_cpu.rf_ram.memory\[5\]\[1\] _05468_ _05506_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13988_ _06951_ _06953_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12939_ _05781_ _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15303__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13979__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14609_ _00463_ net3 mod.u_cpu.rf_ram.memory\[383\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15589_ _01360_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08130_ _02156_ mod.u_cpu.rf_ram.memory\[44\]\[0\] _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15453__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14157__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08061_ _01644_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13904__A1 _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13380__A2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11391__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ mod.u_cpu.cpu.mem_bytecnt\[1\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11518__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13219__I _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08139__A2 _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07914_ _02220_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08894_ _02484_ _03200_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07898__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07845_ mod.u_cpu.rf_ram.memory\[192\]\[0\] mod.u_cpu.rf_ram.memory\[193\]\[0\] mod.u_cpu.rf_ram.memory\[194\]\[0\]
+ mod.u_cpu.rf_ram.memory\[195\]\[0\] _02151_ _02152_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13155__S _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _01671_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09515_ _03738_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08311__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08048__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _03371_ mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09377_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08328_ mod.u_cpu.rf_ram.memory\[501\]\[1\] _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08259_ mod.u_cpu.rf_ram.memory\[535\]\[0\] _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14820__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10009__I0 _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13838__B _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11270_ _04844_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10221_ _04267_ mod.u_cpu.rf_ram.memory\[486\]\[1\] _04264_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13371__A2 _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10152_ _04216_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14970__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11509__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ _04167_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14960_ _00814_ net3 mod.u_cpu.rf_ram.memory\[216\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13911_ _06641_ _06890_ _06891_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14891_ _00745_ net3 mod.u_cpu.rf_ram.memory\[238\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15326__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08550__A2 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13842_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[1\]
+ _06838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10488__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13773_ _06309_ _06666_ _06775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10985_ _04787_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15512_ _01283_ net3 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14350__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__S1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12724_ mod.u_cpu.rf_ram.memory\[137\]\[1\] _05950_ _05972_ _05974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15476__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15443_ _01217_ net3 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12655_ _05742_ _05920_ _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07797__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08066__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11606_ mod.u_cpu.rf_ram.memory\[265\]\[0\] _04954_ _05211_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15374_ _01149_ net3 mod.u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12586_ _05881_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14139__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14325_ _00179_ net3 mod.u_cpu.rf_ram.memory\[525\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07813__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11537_ _01982_ _05165_ _05166_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12208__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14256_ _00110_ net3 mod.u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11468_ _03993_ _04701_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13207_ _06313_ _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08369__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10419_ _04311_ _04404_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14187_ _03842_ _05263_ _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12144__S _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11399_ _05071_ mod.u_cpu.rf_ram.memory\[2\]\[0\] _05072_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11373__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13138_ _06259_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07672__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11983__S _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10971__I1 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13069_ _05742_ _06193_ _06215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12173__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11920__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07630_ _01825_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07561_ _01855_ _01861_ _01868_ _01631_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09300_ _03546_ _03550_ _03551_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07492_ _01770_ _01792_ _01799_ _01768_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09231_ _03487_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14843__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10239__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12928__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _03449_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] _03442_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _01919_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09093_ _03297_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14993__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08044_ _01882_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__A2 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10861__I _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09995_ _04105_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15349__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14223__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13105__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__A2 _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08946_ _01421_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13393__B _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08877_ _02476_ _03180_ _03183_ _02083_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11667__A2 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11692__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08532__A2 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10302__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14373__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07828_ _01862_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15499__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ _02042_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13813__B1 _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08296__A1 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12092__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08934__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _03417_ mod.u_scanchain_local.module_data_in\[68\] _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12440_ _05761_ mod.u_cpu.rf_ram.memory\[172\]\[1\] _05777_ _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13041__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__A2 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12371_ _05734_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14110_ _03823_ _05397_ _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10650__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11322_ _04995_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15090_ _00944_ net3 mod.u_cpu.rf_ram.memory\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14041_ _06970_ _06993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11253_ _04952_ mod.u_cpu.rf_ram.memory\[322\]\[1\] _04970_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10402__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ _04255_ _04234_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11184_ mod.u_cpu.rf_ram.memory\[333\]\[1\] _04819_ _04923_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10135_ _04205_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14716__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10066_ _04148_ mod.u_cpu.rf_ram.memory\[507\]\[0\] _04155_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14943_ _00797_ net3 mod.u_cpu.rf_ram.memory\[221\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08523__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14874_ _00728_ net3 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09072__I _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13825_ _06664_ _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14866__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10011__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13756_ _01479_ _06657_ _06760_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10968_ _04775_ _04759_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10094__A1 _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12707_ _05694_ _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08382__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13687_ _06292_ _06485_ _06294_ _06305_ _06697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11043__S _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _04163_ _04709_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15426_ _01201_ net3 mod.u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12638_ _05916_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14080__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15357_ _01132_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07637__I1 mod.u_cpu.rf_ram.memory\[289\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12569_ _04982_ _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14308_ _00162_ net3 mod.u_cpu.rf_ram.memory\[533\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15288_ _00047_ net4 mod.u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14246__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14239_ _00093_ net3 mod.u_cpu.rf_ram.memory\[568\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12394__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _03001_ _03106_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14396__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09780_ _03954_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07990__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15641__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _03017_ _03030_ _03037_ _02852_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07923__C _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12846__A1 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08514__A2 _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08662_ mod.u_cpu.rf_ram.memory\[223\]\[1\] _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12401__I _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07613_ mod.u_cpu.rf_ram.memory\[317\]\[0\] _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08593_ _01979_ _02899_ _01788_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__I2 _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10085__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11821__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07475_ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13232__I _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09214_ _03480_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15021__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08326__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09145_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12621__I1 mod.u_cpu.rf_ram.memory\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09076_ _03377_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15171__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08027_ _01693_ _02322_ _02334_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__B _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14739__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08061__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_16 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_89_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_27 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09978_ mod.u_cpu.rf_ram.memory\[521\]\[1\] _03929_ _04093_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_38 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12137__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_49 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08929_ mod.u_cpu.rf_ram.memory\[533\]\[1\] _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12837__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14889__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10699__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11940_ _05443_ _05423_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12311__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13851__B _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _05383_ mod.u_cpu.rf_ram.memory\[72\]\[1\] _05392_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13610_ _03365_ _06625_ _06627_ _06629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08269__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ _04511_ _03951_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14590_ _00444_ net3 mod.u_cpu.rf_ram.memory\[392\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09620__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__C _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13541_ _06588_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10753_ _04626_ mod.u_cpu.rf_ram.memory\[401\]\[1\] _04628_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10871__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13472_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _06538_ _06540_ _03588_ _06542_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10684_ _04522_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07492__A2 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14269__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15211_ _01064_ net3 mod.u_cpu.rf_ram.memory\[199\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12423_ _05753_ mod.u_cpu.rf_ram.memory\[174\]\[0\] _05768_ _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08116__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15514__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11576__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15142_ _00995_ net3 mod.u_cpu.rf_ram.memory\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12354_ _05452_ _05721_ _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11305_ _05007_ mod.u_cpu.rf_ram.memory\[314\]\[0\] _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15073_ _00927_ net3 mod.u_cpu.rf_ram.memory\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12285_ _05563_ _03859_ _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14024_ _06979_ _06980_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11236_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10000__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11167_ _04067_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _04192_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11098_ _04862_ mod.u_cpu.rf_ram.memory\[347\]\[1\] _04865_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12221__I _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ _04117_ mod.u_cpu.rf_ram.memory\[510\]\[0\] _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14926_ _00780_ net3 mod.u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14857_ _00711_ net3 mod.u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15044__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13808_ _06418_ _06449_ _06807_ _06442_ _06808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14788_ _00642_ net3 mod.u_cpu.rf_ram.memory\[293\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12300__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13739_ _06713_ _06744_ _06745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08355__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11803__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13052__I _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08146__I _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _01497_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15194__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15409_ _01184_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07191_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14084__S _07022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11501__S _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07985__I _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08432__A1 _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08983__A2 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09901_ _03697_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09832_ _01478_ _03993_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08735__A2 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08291__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12119__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09705__I _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__C _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12819__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08714_ mod.u_cpu.rf_ram.memory\[229\]\[1\] _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08499__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09694_ _03885_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08043__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07225__I _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08645_ _02110_ _02948_ _02951_ _02141_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08594__S1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08576_ _01979_ _02875_ _02882_ _01989_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14411__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09999__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07527_ _01818_ _01834_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15537__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10853__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08671__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07389_ _01633_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14561__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _03416_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__S _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ _03315_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09816__S _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12070_ _05529_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07609__S0 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11021_ _04812_ _04788_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15067__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08034__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12972_ _06142_ _06146_ _06147_ _06145_ _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _05431_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14711_ _00565_ net3 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14642_ _00496_ net3 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13235__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11854_ _05366_ mod.u_cpu.rf_ram.memory\[6\]\[0\] _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _04663_ mod.u_cpu.rf_ram.memory\[392\]\[0\] _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13786__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14573_ _00427_ net3 mod.u_cpu.rf_ram.memory\[401\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11785_ _05262_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13524_ _03923_ _06577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ _04598_ mod.u_cpu.rf_ram.memory\[403\]\[0\] _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14904__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13455_ _06530_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10667_ _01712_ _04571_ _04572_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12597__I0 _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12406_ _05756_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08414__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13386_ _06480_ _06447_ _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04525_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15125_ _00978_ net3 mod.u_cpu.rf_ram.memory\[459\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12337_ _05709_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11120__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15056_ _00910_ net3 mod.u_cpu.rf_ram.memory\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12268_ _05662_ mod.u_cpu.rf_ram.memory\[192\]\[0\] _05663_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14007_ _03456_ _06964_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _06968_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09914__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _04936_ mod.u_cpu.rf_ram.memory\[327\]\[1\] _04946_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13710__A2 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12199_ _05616_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12521__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14434__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14909_ _00763_ net3 mod.u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12886__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ mod.u_cpu.rf_ram.memory\[407\]\[1\] _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13226__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12029__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08361_ _01960_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ _01592_ _01601_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14584__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ mod.u_cpu.rf_ram.memory\[453\]\[1\] _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07456__A2 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08653__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _01550_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _01472_ _01473_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10063__I1 mod.u_cpu.rf_ram.memory\[508\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11260__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11030__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11012__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12760__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ _03757_ _03980_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08479__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _03927_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08016__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12512__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08628_ _02090_ _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13217__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14927__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08559_ _01963_ _02865_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11779__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08644__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__A2 _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11570_ _05187_ _05130_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10521_ _04474_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07839__B _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12464__C _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13240_ _05396_ _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10452_ _04426_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14193__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11251__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13171_ _03510_ _06278_ _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10383_ _04377_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14307__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12122_ _05563_ _03843_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11875__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12053_ _05483_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12751__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11004_ mod.u_cpu.rf_ram.memory\[361\]\[1\] _04661_ _04799_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14457__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07383__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12700__S _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07773__I3 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12955_ _06131_ _06132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11906_ _05419_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13208__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12886_ _05396_ _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13759__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10690__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14625_ _00479_ net3 mod.u_cpu.rf_ram.memory\[375\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11837_ _05364_ mod.u_cpu.rf_ram.memory\[228\]\[1\] _05368_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14556_ _00410_ net3 mod.u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08635__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11768_ _02246_ _05321_ _05323_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10442__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13507_ mod.u_cpu.cpu.ctrl.i_jump _03296_ _06562_ _06563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10719_ _04598_ mod.u_cpu.rf_ram.memory\[406\]\[0\] _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10954__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11490__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14487_ _00341_ net3 mod.u_cpu.rf_ram.memory\[444\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11699_ _05275_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13438_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _06519_ _06520_ _03520_ _06521_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_13369_ _06464_ _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15232__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15108_ _00962_ net3 mod.u_cpu.rf_ram.memory\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11785__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15039_ _00893_ net3 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07930_ _01819_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07861_ _02150_ _02153_ _02167_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15382__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09600_ _03800_ mod.u_cpu.rf_ram.memory\[56\]\[1\] _03811_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07792_ _02097_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09531_ _03754_ _03721_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13998__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07931__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11226__S _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09462_ _03686_ _03687_ _03688_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _02539_ _02712_ _02719_ _01678_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09393_ _03623_ _03629_ _03630_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08344_ _02597_ _02647_ _02650_ _01651_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08626__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12422__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10433__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08275_ _01459_ _02558_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13240__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ _01533_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07157_ _01464_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11933__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14071__I _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13686__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09165__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12733__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08788__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08002__C _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13438__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09729_ _03890_ mod.u_cpu.rf_ram.memory\[555\]\[1\] _03912_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12110__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11136__S _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12459__C _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12740_ _05937_ _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07668__A2 _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15105__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10672__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12671_ _05938_ mod.u_cpu.rf_ram.memory\[121\]\[1\] _05935_ _05939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14410_ _00264_ net3 mod.u_cpu.rf_ram.memory\[482\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11622_ _05221_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15390_ _01165_ net3 mod.u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14341_ _00195_ net3 mod.u_cpu.rf_ram.memory\[517\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10424__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10275__I1 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11553_ _05176_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10975__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10504_ _04450_ mod.u_cpu.rf_ram.memory\[442\]\[1\] _04461_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15255__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14272_ _00126_ net3 mod.u_cpu.rf_ram.memory\[551\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11484_ _05119_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10027__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13223_ _06329_ _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13913__A2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ mod.u_cpu.rf_ram.memory\[453\]\[1\] _04383_ _04413_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13154_ _06252_ _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10366_ _04368_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12105_ _03850_ _05552_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13085_ _06217_ mod.u_cpu.rf_ram.memory\[104\]\[1\] _06224_ _06226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10297_ _04321_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09075__I _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12036_ _05507_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13987_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _06952_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _06953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13325__I _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12938_ _06115_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07323__I _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12869_ _06035_ mod.u_cpu.rf_ram.memory\[409\]\[0\] _06068_ _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14608_ _00462_ net3 mod.u_cpu.rf_ram.memory\[383\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15588_ _01359_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10684__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14539_ _00393_ net3 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08154__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ mod.u_cpu.rf_ram.memory\[72\]\[0\] mod.u_cpu.rf_ram.memory\[73\]\[0\] mod.u_cpu.rf_ram.memory\[74\]\[0\]
+ mod.u_cpu.rf_ram.memory\[75\]\[0\] _02366_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12168__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14622__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11391__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08962_ mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r _03266_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13668__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14772__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ mod.u_cpu.rf_ram.memory\[215\]\[0\] _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08893_ mod.u_cpu.rf_ram.memory\[567\]\[1\] _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07347__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07844_ _02126_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15128__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07775_ _01785_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ _03737_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09445_ _01451_ _03674_ mod.u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15278__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09376_ _03614_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10594__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08327_ mod.u_cpu.rf_ram.memory\[496\]\[1\] mod.u_cpu.rf_ram.memory\[497\]\[1\] mod.u_cpu.rf_ram.memory\[498\]\[1\]
+ mod.u_cpu.rf_ram.memory\[499\]\[1\] _02632_ _02633_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_36_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11454__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _02245_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12159__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__I1 mod.u_cpu.rf_ram.memory\[516\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _01516_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11206__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08189_ mod.u_cpu.rf_ram.memory\[573\]\[0\] _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10220_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07836__C _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _04215_ mod.u_cpu.rf_ram.memory\[495\]\[1\] _04213_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12314__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07408__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10082_ _04157_ mod.u_cpu.rf_ram.memory\[505\]\[1\] _04165_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13910_ _03679_ _06649_ _06891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14890_ _00744_ net3 mod.u_cpu.rf_ram.memory\[238\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10893__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13841_ _05787_ _06834_ _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10769__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13145__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13772_ _06773_ _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10984_ _04772_ mod.u_cpu.rf_ram.memory\[364\]\[1\] _04785_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13831__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15511_ _01282_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12723_ _05973_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11693__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15442_ _01216_ net3 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _05927_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14645__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11605_ _05078_ _05210_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11445__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15373_ _01148_ net3 mod.u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12585_ _05874_ mod.u_cpu.rf_ram.memory\[157\]\[1\] _05879_ _05881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09263__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14324_ _00178_ net3 mod.u_cpu.rf_ram.memory\[525\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14139__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11536_ _05133_ _05165_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13347__B1 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14255_ _00109_ net3 mod.u_cpu.rf_ram.memory\[560\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11467_ _05117_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13898__A1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13206_ _06312_ _06313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14795__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10418_ _03942_ _04335_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14186_ _07088_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11398_ _04196_ _03975_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12570__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13137_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _06258_ _06259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _04201_ _04353_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07672__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13068_ _06214_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12322__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12019_ _05496_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10184__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08621__S0 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09533__I _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07481__C _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07560_ _01863_ mod.u_cpu.rf_ram.memory\[382\]\[0\] _01866_ _01867_ _01868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08149__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15420__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13822__B2 _06820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07491_ _01773_ _01795_ _01798_ _01785_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07501__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08593__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09230_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ mod.u_arbiter.i_wb_cpu_rdt\[10\] _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15570__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09254__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11303__I _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08112_ mod.u_cpu.rf_ram.memory\[52\]\[0\] mod.u_cpu.rf_ram.memory\[53\]\[0\] mod.u_cpu.rf_ram.memory\[54\]\[0\]
+ mod.u_cpu.rf_ram.memory\[55\]\[0\] _02403_ _02152_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_148_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09092_ _03362_ _03392_ _03300_ _03279_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ mod.u_cpu.rf_ram.memory\[64\]\[0\] mod.u_cpu.rf_ram.memory\[65\]\[0\] mod.u_cpu.rf_ram.memory\[66\]\[0\]
+ mod.u_cpu.rf_ram.memory\[67\]\[0\] _02349_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09708__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09801__I0 _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09994_ _04091_ mod.u_cpu.rf_ram.memory\[518\]\[1\] _04103_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08945_ _01440_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08876_ _02483_ mod.u_cpu.rf_ram.memory\[558\]\[1\] _03182_ _02487_ _03183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14518__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08612__S0 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09443__I _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08487__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14066__A1 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14066__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13113__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _01704_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14668__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08296__A2 _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07689_ _01960_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09428_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _03657_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11427__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09359_ _03489_ _03600_ _03601_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13041__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11978__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12370_ _05731_ mod.u_cpu.rf_ram.memory\[499\]\[0\] _05733_ _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _03821_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10650__I1 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14040_ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _06989_ _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11252_ _04971_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10203_ _03932_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11183_ _04924_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07138__I _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _04199_ mod.u_cpu.rf_ram.memory\[498\]\[1\] _04203_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08678__B _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10065_ _03791_ _04143_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14942_ _00796_ net3 mod.u_cpu.rf_ram.memory\[221\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15443__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14057__A1 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14873_ _00727_ net3 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13824_ _06821_ _06822_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13755_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _06753_ _06709_ _06759_ _06760_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15593__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09484__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10967_ _03884_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13280__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10094__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12706_ _05961_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13686_ _06424_ _06682_ _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10898_ _04694_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15425_ _01200_ net3 mod.u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09236__A1 _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12637_ _05904_ mod.u_cpu.rf_ram.memory\[148\]\[0\] _05915_ _05916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14080__I1 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12568_ _05812_ _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15356_ _01131_ net3 mod.u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14307_ _00161_ net3 mod.u_cpu.rf_ram.memory\[534\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _05154_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10641__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12499_ _05825_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15287_ _00046_ net4 mod.u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09528__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12918__I0 mod.u_cpu.rf_ram.memory\[389\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14238_ _00092_ net3 mod.u_cpu.rf_ram.memory\[568\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07476__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14169_ _05780_ _07067_ _07077_ _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__A2 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07970__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _02043_ _03033_ _03036_ _01695_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12846__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08661_ _02450_ mod.u_cpu.rf_ram.memory\[220\]\[1\] _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14810__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07612_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08592_ mod.u_cpu.rf_ram.memory\[264\]\[1\] mod.u_cpu.rf_ram.memory\[265\]\[1\] mod.u_cpu.rf_ram.memory\[266\]\[1\]
+ mod.u_cpu.rf_ram.memory\[267\]\[1\] _01802_ _01932_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11657__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07543_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07474_ _01700_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14960__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09213_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] _03479_
+ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11033__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09144_ _03434_ _03435_ _03437_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08770__C _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15316__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ _03334_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09438__I _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08026_ _02293_ _02324_ _02333_ _02291_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14340__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15466__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_17 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_28 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09977_ _04094_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_39 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ mod.u_cpu.rf_ram.memory\[528\]\[1\] mod.u_cpu.rf_ram.memory\[529\]\[1\] mod.u_cpu.rf_ram.memory\[530\]\[1\]
+ mod.u_cpu.rf_ram.memory\[531\]\[1\] _02528_ _02543_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12837__A2 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14490__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08859_ _01471_ _03116_ _03165_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11870_ _05393_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09901__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _04675_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13262__A2 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13423__I _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10752_ _04629_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13540_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] mod.u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _06584_ _06588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11273__A1 _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ _06541_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10683_ _04583_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15210_ _01063_ net3 mod.u_cpu.rf_ram.memory\[199\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12422_ _05312_ _05767_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08453__S _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15141_ _00994_ net3 mod.u_cpu.rf_ram.memory\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12353_ _05720_ _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13298__C _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11304_ _04868_ _04990_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08252__I _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15072_ _00926_ net3 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12284_ _05674_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14023_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _06976_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11235_ _03737_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08824__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12703__S _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10000__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__A2 _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _04912_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14833__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _04178_ mod.u_cpu.rf_ram.memory\[500\]\[1\] _04190_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12502__I _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10139__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11097_ _04866_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09083__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10048_ _03752_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14925_ _00779_ net3 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14856_ _00710_ net3 mod.u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14983__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08855__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13807_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_arbiter.i_wb_cpu_rdt\[11\] _03509_
+ _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14787_ _00641_ net3 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11999_ _02221_ _05481_ _05482_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11054__S _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13738_ _06743_ _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15339__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13669_ _06658_ _06680_ _06681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15408_ _01183_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07190_ _01497_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08590__C _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13961__B1 _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11811__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15339_ _01114_ net3 mod.u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14363__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15489__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09258__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09900_ _03837_ _04033_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13713__B1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09831_ _03754_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08291__S1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12119__I1 mod.u_cpu.rf_ram.memory\[210\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07943__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12412__I _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09762_ _03818_ _03939_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12819__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08713_ mod.u_cpu.rf_ram.memory\[224\]\[1\] mod.u_cpu.rf_ram.memory\[225\]\[1\] mod.u_cpu.rf_ram.memory\[226\]\[1\]
+ mod.u_cpu.rf_ram.memory\[227\]\[1\] _01507_ _01763_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09693_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08043__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08644_ _02115_ mod.u_cpu.rf_ram.memory\[174\]\[1\] _02950_ _01771_ _02951_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10550__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _01981_ _02878_ _02881_ _01972_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09448__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ _01822_ _01824_ _01829_ _01831_ _01832_ _01833_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09999__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10302__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08120__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07457_ _01527_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14706__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07388_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_135_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09058_ _03306_ _03360_ _03346_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08072__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08009_ mod.u_cpu.rf_ram.memory\[127\]\[0\] _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14856__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__S1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13180__A1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _03949_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13862__B _06855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11869__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10978__S _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12971_ mod.u_cpu.cpu.genblk3.csr.mstatus_mpie _06142_ _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08034__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14710_ _00564_ net3 mod.u_cpu.rf_ram.memory\[332\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _05426_ mod.u_cpu.rf_ram.memory\[222\]\[1\] _05429_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09631__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14236__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14641_ _00495_ net3 mod.u_cpu.rf_ram.memory\[367\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11853_ _05239_ _03951_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13235__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10804_ _04255_ _04648_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08247__I _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11784_ _03917_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14572_ _00426_ net3 mod.u_cpu.rf_ram.memory\[401\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07151__I _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08111__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07545__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13523_ _06576_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10735_ _04352_ _04599_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14386__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11602__S _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10666_ _04542_ _04571_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13454_ _03547_ _06525_ _06526_ _03552_ _06530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__15631__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _05745_ mod.u_cpu.rf_ram.memory\[176\]\[1\] _05754_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13385_ _06397_ _06129_ _06480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10597_ _04523_ mod.u_cpu.rf_ram.memory\[426\]\[0\] _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09611__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15124_ _00977_ net3 mod.u_cpu.rf_ram.memory\[459\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12336_ _05105_ _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12267_ _05417_ _05650_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15055_ _00909_ net3 mod.u_cpu.rf_ram.memory\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13171__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09806__I _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14006_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _06966_ _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11218_ _04947_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08710__I _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12198_ mod.u_cpu.rf_ram.memory\[201\]\[0\] _05437_ _05615_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07754__C _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ _04882_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15011__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07326__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09678__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14908_ _00762_ net3 mod.u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11485__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09541__I _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15161__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14839_ _00693_ net3 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13226__A2 _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08360_ mod.u_cpu.rf_ram.memory\[480\]\[1\] mod.u_cpu.rf_ram.memory\[481\]\[1\] mod.u_cpu.rf_ram.memory\[482\]\[1\]
+ mod.u_cpu.rf_ram.memory\[483\]\[1\] _01963_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08157__I _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14729__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07311_ _01602_ _01606_ _01617_ _01618_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12985__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08291_ mod.u_cpu.rf_ram.memory\[448\]\[1\] mod.u_cpu.rf_ram.memory\[449\]\[1\] mod.u_cpu.rf_ram.memory\[450\]\[1\]
+ mod.u_cpu.rf_ram.memory\[451\]\[1\] _01508_ _02597_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09850__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07242_ mod.u_cpu.raddr\[3\] _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10460__A2 _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12737__A1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14879__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07173_ _01478_ _01479_ _01480_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12407__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10599__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09716__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07916__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09814_ _03979_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14259__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09745_ mod.u_cpu.rf_ram.memory\[553\]\[0\] _03925_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09669__A1 _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08016__S1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11981__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15504__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07680__B _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ mod.u_cpu.rf_ram.memory\[176\]\[1\] mod.u_cpu.rf_ram.memory\[177\]\[1\] mod.u_cpu.rf_ram.memory\[178\]\[1\]
+ mod.u_cpu.rf_ram.memory\[179\]\[1\] _02048_ _02086_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13217__A2 _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__A2 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12276__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08558_ mod.u_cpu.rf_ram.memory\[309\]\[1\] _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11779__A2 _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07509_ _01656_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ _02778_ _02788_ _02795_ _02677_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10520_ _04469_ mod.u_cpu.rf_ram.memory\[43\]\[0\] _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10451_ _04410_ mod.u_cpu.rf_ram.memory\[450\]\[1\] _04424_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13170_ _03492_ _03412_ _03400_ _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_184_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10382_ _04225_ _04379_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12121_ _04982_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15034__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ _05517_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11003_ _04800_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08580__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07383__A2 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15184__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12954_ _06125_ _06128_ _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11905_ _05413_ mod.u_cpu.rf_ram.memory\[224\]\[0\] _05418_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13208__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12885_ _06079_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14624_ _00478_ net3 mod.u_cpu.rf_ram.memory\[375\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10690__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11836_ _05369_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12967__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14555_ _00409_ net3 mod.u_cpu.rf_ram.memory\[410\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09832__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11767_ _05322_ _05321_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13506_ _06142_ _03250_ _06562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10718_ _04180_ _04599_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14486_ _00340_ net3 mod.u_cpu.rf_ram.memory\[444\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11698_ _05271_ mod.u_cpu.rf_ram.memory\[254\]\[1\] _05273_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13437_ _06513_ _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10649_ _04497_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13392__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13368_ _06388_ _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13767__B _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15107_ _00961_ net3 mod.u_cpu.rf_ram.memory\[439\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12319_ _05698_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12163__S _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13299_ _06328_ _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09199__I0 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15038_ _00892_ net3 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14401__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15527__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07860_ _01586_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10753__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08571__A1 _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07791_ mod.u_cpu.rf_ram.memory\[188\]\[0\] mod.u_cpu.rf_ram.memory\[189\]\[0\] mod.u_cpu.rf_ram.memory\[190\]\[0\]
+ mod.u_cpu.rf_ram.memory\[191\]\[0\] _02092_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09530_ _03716_ _03717_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14551__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09461_ _03681_ _03679_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ _02654_ _02715_ _02718_ _01992_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09392_ _03496_ mod.u_scanchain_local.module_data_in\[62\] _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08343_ _02638_ mod.u_cpu.rf_ram.memory\[510\]\[1\] _02649_ _01821_ _02650_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09823__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ _02571_ _02581_ _02520_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11630__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13907__B1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13758__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07225_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15057__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13383__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _01438_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12430__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11233__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11933__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13686__A2 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08562__A1 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07989_ _02091_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10321__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09728_ _03913_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12110__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09659_ _03858_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10672__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12670_ _05937_ _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _04959_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14340_ _00194_ net3 mod.u_cpu.rf_ram.memory\[517\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11552_ _05159_ mod.u_cpu.rf_ram.memory\[274\]\[0\] _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09290__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _04462_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14271_ _00125_ net3 mod.u_cpu.rf_ram.memory\[552\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11483_ _05129_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12177__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13222_ _06328_ _06129_ _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10434_ _01512_ _04413_ _04415_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14424__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11886__I _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10365_ _04363_ mod.u_cpu.rf_ram.memory\[464\]\[1\] _04366_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13153_ _06267_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12104_ _05432_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13084_ _06225_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10296_ _04313_ mod.u_cpu.rf_ram.memory\[475\]\[1\] _04319_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13677__A2 _06685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12724__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12035_ mod.u_cpu.rf_ram.memory\[5\]\[0\] _05437_ _05506_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14574__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11327__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13986_ _06937_ _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09091__I mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12937_ _06057_ _06114_ _06115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11160__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15821__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12868_ _05896_ _04687_ _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14607_ _00461_ net3 mod.u_cpu.rf_ram.memory\[384\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11819_ _05350_ mod.u_cpu.rf_ram.memory\[230\]\[1\] _05356_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15587_ _01358_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12799_ _06019_ mod.u_cpu.rf_ram.memory\[12\]\[1\] _06021_ _06023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14538_ _00392_ net3 mod.u_cpu.rf_ram.memory\[418\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07292__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14469_ _00323_ net3 mod.u_cpu.rf_ram.memory\[453\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11796__I _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14917__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08170__I _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08961_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _03265_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07912_ _01519_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08892_ _02478_ mod.u_cpu.rf_ram.memory\[564\]\[1\] _03198_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07347__A2 _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__A1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _01856_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07774_ _02080_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09513_ _03695_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11151__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09444_ _03353_ _03673_ _03674_ mod.u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10875__I _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09375_ _03486_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13251__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ _01637_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11454__I1 mod.u_cpu.rf_ram.memory\[290\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14447__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08257_ _02527_ mod.u_cpu.rf_ram.memory\[532\]\[0\] _02564_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07208_ _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12159__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ mod.u_cpu.rf_ram.memory\[568\]\[0\] mod.u_cpu.rf_ram.memory\[569\]\[0\] mod.u_cpu.rf_ram.memory\[570\]\[0\]
+ mod.u_cpu.rf_ram.memory\[571\]\[0\] _02494_ _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12403__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07139_ _01439_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09176__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14597__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ _04177_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08080__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10081_ _04166_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09583__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11147__S _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13426__I _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13840_ _06835_ _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10893__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13771_ _06415_ _06772_ _06773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_90_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10983_ _04786_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11142__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15510_ _01281_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ mod.u_cpu.rf_ram.memory\[137\]\[0\] _05971_ _05972_ _05973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15222__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12890__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08683__C _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15441_ _01215_ net3 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12653_ _05923_ mod.u_cpu.rf_ram.memory\[146\]\[1\] _05925_ _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11604_ _03723_ _04779_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15372_ _01147_ net3 mod.u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11445__I1 mod.u_cpu.rf_ram.memory\[291\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12584_ _05880_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14323_ _00177_ net3 mod.u_cpu.rf_ram.memory\[526\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15372__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11535_ _05164_ _05130_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13347__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13347__B2 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14254_ _00108_ net3 mod.u_cpu.rf_ram.memory\[560\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _05108_ mod.u_cpu.rf_ram.memory\[288\]\[1\] _05115_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13898__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13205_ mod.u_arbiter.i_wb_cpu_rdt\[8\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _03499_ _06312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10417_ _04403_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14185_ _07081_ mod.u_cpu.rf_ram.memory\[279\]\[1\] _07086_ _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11397_ _05045_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10956__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09086__I _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14147__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13136_ _06252_ _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12570__A2 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10348_ _04356_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10279_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13067_ _06199_ mod.u_cpu.rf_ram.memory\[106\]\[1\] _06212_ _06214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12322__A2 _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12018_ _05470_ mod.u_cpu.rf_ram.memory\[214\]\[0\] _05495_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08621__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13780__B _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10896__S _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12086__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13969_ _06936_ _06939_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13822__A2 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07490_ _01689_ mod.u_cpu.rf_ram.memory\[438\]\[0\] _01797_ _01763_ _01798_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15639_ _01410_ net3 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09160_ _03448_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08165__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08111_ _01693_ _02392_ _02418_ _02380_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_187_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09091_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ _01637_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13889__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09993_ _04104_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10572__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08944_ _03249_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08517__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08768__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _02484_ _03181_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08612__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12150__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07826_ _01634_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15245__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07244__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13113__I1 mod.u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07757_ _01849_ _02064_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12872__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ mod.u_cpu.rf_ram.memory\[280\]\[0\] mod.u_cpu.rf_ram.memory\[281\]\[0\] mod.u_cpu.rf_ram.memory\[282\]\[0\]
+ mod.u_cpu.rf_ram.memory\[283\]\[0\] _01994_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09493__A2 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09427_ mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15395__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12624__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09358_ _03554_ mod.u_scanchain_local.module_data_in\[57\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ _02532_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09289_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13329__A1 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11320_ _05018_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ _04961_ mod.u_cpu.rf_ram.memory\[322\]\[0\] _04970_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _04254_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11182_ mod.u_cpu.rf_ram.memory\[333\]\[0\] _04658_ _04923_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10133_ _04204_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08508__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08678__C _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10064_ _04154_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14941_ _00795_ net3 mod.u_cpu.rf_ram.memory\[222\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11363__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14872_ _00726_ net3 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14057__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07154__I _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13823_ mod.u_cpu.cpu.immdec.imm30_25\[3\] _06773_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[4\]
+ _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12068__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12995__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14612__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13754_ _06432_ _06755_ _06758_ _06065_ _06759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10618__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10966_ _04694_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12705_ mod.u_cpu.rf_ram.memory\[13\]\[1\] _05950_ _05959_ _05961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13685_ _06694_ _06398_ _06695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10897_ _04727_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15424_ _01199_ net3 mod.u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12615__I0 _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14762__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12636_ _05535_ _05900_ _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15355_ _01130_ net3 mod.u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12567_ _05868_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13759__C _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11340__S _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14306_ _00160_ net3 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11518_ _05144_ mod.u_cpu.rf_ram.memory\[280\]\[0\] _05153_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15286_ _00045_ net4 mod.u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12498_ _05813_ mod.u_cpu.rf_ram.memory\[459\]\[0\] _05824_ _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15118__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12918__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14237_ _00091_ net3 mod.u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11449_ _05104_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09745__S _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13740__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14168_ _05790_ _06166_ _03393_ _07073_ _07077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13119_ _06247_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15268__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14099_ _07032_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09544__I _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07492__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10306__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08660_ _02656_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14292__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07611_ _01743_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14098__S _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _02759_ _02894_ _02897_ _02764_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11515__S _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07542_ _01490_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11657__I1 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09475__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__A1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07473_ _01779_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09212_ _03414_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A2 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09143_ mod.u_arbiter.i_wb_cpu_rdt\[4\] _03436_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08986__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09074_ _03370_ _03376_ mod.u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08025_ _02325_ _02328_ _02332_ _01717_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13031__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13731__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07410__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ mod.u_cpu.rf_ram.memory\[521\]\[0\] _03925_ _04093_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_18 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_29 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08498__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08927_ _02523_ _03226_ _03233_ _02505_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14635__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _01475_ _03141_ _03164_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_73_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ mod.u_cpu.rf_ram.memory\[175\]\[0\] _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08789_ _01493_ _03095_ _01534_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ _04666_ mod.u_cpu.rf_ram.memory\[390\]\[1\] _04673_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14785__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _04622_ mod.u_cpu.rf_ram.memory\[401\]\[0\] _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11273__A2 _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11224__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _03578_ _06538_ _06540_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _06541_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_164_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _04579_ mod.u_cpu.rf_ram.memory\[413\]\[1\] _04581_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _05725_ _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12222__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11160__S _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15140_ _00993_ net3 mod.u_cpu.rf_ram.memory\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13970__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12352_ _05629_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11303_ _04960_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13022__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15071_ _00925_ net3 mod.u_cpu.rf_ram.memory\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12283_ _05660_ mod.u_cpu.rf_ram.memory\[190\]\[1\] _05672_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__I _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08729__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14022_ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] _06978_ _06979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15410__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13722__A1 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09777__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__A2 _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11234_ _04958_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10387__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11165_ _04896_ mod.u_cpu.rf_ram.memory\[336\]\[1\] _04910_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07952__A2 mod.u_cpu.rf_ram.memory\[244\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _04191_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11096_ _04864_ mod.u_cpu.rf_ram.memory\[347\]\[0\] _04865_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15560__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10047_ _04142_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14924_ _00778_ net3 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14855_ _00709_ net3 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _06735_ _06802_ _06805_ _06332_ _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14786_ _00640_ net3 mod.u_cpu.rf_ram.memory\[294\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11998_ _05448_ _05481_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09457__A2 _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07612__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13737_ _06288_ _06667_ _06669_ _06743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12461__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ _04511_ _03961_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13668_ _06677_ _06679_ _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14202__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15407_ _01182_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12619_ _05886_ _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07768__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13599_ _03694_ _06573_ _06620_ _03659_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__14508__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09539__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13961__A1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15338_ _01113_ net3 mod.u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10775__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07640__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15269_ _00026_ net4 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13013__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15090__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13713__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13713__B2 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14658__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08815__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09393__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ _03806_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _03746_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11327__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08111__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _03017_ _03018_ _01870_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09692_ _03856_ _03883_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _02116_ _02949_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13524__I _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08574_ _01697_ mod.u_cpu.rf_ram.memory\[278\]\[1\] _02880_ _01952_ _02881_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_148_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09448__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07459__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07525_ _01679_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08120__A2 _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07456_ _01689_ mod.u_cpu.rf_ram.memory\[422\]\[0\] _01761_ _01763_ _01764_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_168_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07387_ _01491_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08959__A1 _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15433__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _03423_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08353__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10766__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09057_ _03355_ mod.u_cpu.cpu.csr_imm _03358_ _03359_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13704__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08008_ _01924_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15583__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13180__A2 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09959_ _04082_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12970_ _03369_ _06146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13862__C _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11869__I1 mod.u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09912__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _05430_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07698__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12691__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14640_ _00494_ net3 mod.u_cpu.rf_ram.memory\[367\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09133__B _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11852_ _05380_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07432__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10803_ _04621_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14571_ _00425_ net3 mod.u_cpu.rf_ram.memory\[402\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _05333_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08972__B _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08111__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13522_ _03426_ _06575_ _06570_ _06576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07545__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10734_ _04616_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14196__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13453_ _06529_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10665_ _03991_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12404_ _05755_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13384_ _03663_ _06356_ _06416_ _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10596_ _04242_ _04507_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09611__A2 _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15123_ _00976_ net3 mod.u_cpu.rf_ram.memory\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07622__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12335_ _05708_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14800__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15054_ _00908_ net3 mod.u_cpu.rf_ram.memory\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12266_ _05604_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14005_ _06942_ _06966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11217_ _04938_ mod.u_cpu.rf_ram.memory\[327\]\[0\] _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12197_ _05588_ _05594_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09094__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14950__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07607__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _04900_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13545__S _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11079_ _04854_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09678__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09822__I _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07233__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14907_ _00761_ net3 mod.u_cpu.rf_ram.memory\[231\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07770__C _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11485__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15306__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13344__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14838_ _00692_ net3 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14769_ _00623_ net3 mod.u_cpu.rf_ram.memory\[303\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10296__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14330__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07310_ _01551_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15456__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ _01882_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09850__A2 _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14187__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07241_ _01505_ _01544_ _01548_ _01529_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12037__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09989__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07172_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _01467_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13934__A1 _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14480__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08106__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__I1 mod.u_cpu.rf_ram.memory\[425\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09813_ _03768_ _03966_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__I1 mod.u_cpu.rf_ram.memory\[398\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ _03714_ _03893_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09732__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09669__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09675_ _03870_ _03848_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08626_ _01486_ _02923_ _02932_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_54_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07252__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ mod.u_cpu.rf_ram.memory\[304\]\[1\] mod.u_cpu.rf_ram.memory\[305\]\[1\] mod.u_cpu.rf_ram.memory\[306\]\[1\]
+ mod.u_cpu.rf_ram.memory\[307\]\[1\] _01994_ _02010_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07508_ _01694_ _01737_ _01738_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08488_ _02668_ _02791_ _02794_ _02096_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10987__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07439_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07852__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14823__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13925__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10450_ _04425_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08083__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11787__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09109_ _03385_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07604__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ _04378_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14973__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12120_ _05562_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12051_ _05498_ mod.u_cpu.rf_ram.memory\[61\]\[0\] _05516_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11002_ mod.u_cpu.rf_ram.memory\[361\]\[0\] _04658_ _04799_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15329__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10911__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12953_ _06125_ _06129_ _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11904_ _05417_ _05401_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14353__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08258__I _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15479__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12884_ _06070_ mod.u_cpu.rf_ram.memory\[99\]\[1\] _06077_ _06079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__I _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07391__I0 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14623_ _00477_ net3 mod.u_cpu.rf_ram.memory\[376\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11835_ _05366_ mod.u_cpu.rf_ram.memory\[228\]\[0\] _05368_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14554_ _00408_ net3 mod.u_cpu.rf_ram.memory\[410\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _03944_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09832__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14169__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13505_ _06561_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10717_ _04605_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14485_ _00339_ net3 mod.u_cpu.rf_ram.memory\[445\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12508__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11697_ _05274_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13436_ _06510_ _06519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10648_ _04559_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13367_ _06308_ _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _04506_ mod.u_cpu.rf_ram.memory\[42\]\[0\] _04512_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15106_ _00960_ net3 mod.u_cpu.rf_ram.memory\[439\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12318_ _05696_ mod.u_cpu.rf_ram.memory\[189\]\[0\] _05697_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13298_ _06289_ _06390_ _06394_ _06373_ _06395_ _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_170_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09348__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15037_ _00891_ net3 mod.u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12249_ _05649_ _05650_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07337__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11950__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ _01637_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09552__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12655__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09520__A1 _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _03388_ _03337_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_149_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08168__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07382__I0 mod.u_cpu.rf_ram.memory\[396\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08411_ _02656_ mod.u_cpu.rf_ram.memory\[446\]\[1\] _02717_ _01961_ _02718_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14846__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] _03615_ _03628_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_145_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11523__S _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08342_ _02220_ _02648_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09823__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _02542_ _02572_ _02580_ _02491_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07834__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11630__A2 _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11322__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07224_ _01531_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14996__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13907__B2 _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13758__I1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13383__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__B _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14226__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08011__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13185__S _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11941__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__A2 _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14376__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08279__S _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ mod.u_cpu.rf_ram.memory\[104\]\[0\] mod.u_cpu.rf_ram.memory\[105\]\[0\] mod.u_cpu.rf_ram.memory\[106\]\[0\]
+ mod.u_cpu.rf_ram.memory\[107\]\[0\] _02294_ _02295_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__15621__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09727_ _03877_ mod.u_cpu.rf_ram.memory\[555\]\[0\] _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _03857_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08078__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08609_ _02040_ _02915_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09589_ _03779_ _03786_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11620_ _05220_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07825__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ _04758_ _05171_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10502_ _04453_ mod.u_cpu.rf_ram.memory\[442\]\[0\] _04461_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15001__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14270_ _00124_ net3 mod.u_cpu.rf_ram.memory\[552\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11482_ _05128_ mod.u_cpu.rf_ram.memory\[286\]\[1\] _05126_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13221_ _03501_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _06327_ _06328_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10433_ _04414_ _04413_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11385__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13152_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _06263_ _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10364_ _04367_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15151__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12103_ _05551_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13083_ _06205_ mod.u_cpu.rf_ram.memory\[104\]\[0\] _06224_ _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10295_ _04320_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14719__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08002__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12034_ _03728_ _04955_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11608__S _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13985_ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _06943_ _06951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14869__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09502__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10499__I0 _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12936_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _06111_ _06112_ _06113_ _06063_ _06114_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12867_ _03677_ _06066_ _06067_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11860__A2 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11343__S _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14606_ _00460_ net3 mod.u_cpu.rf_ram.memory\[384\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11818_ _05357_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15586_ _01357_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12798_ _06022_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14537_ _00391_ net3 mod.u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11749_ _03696_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14468_ _00322_ net3 mod.u_cpu.rf_ram.memory\[453\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14249__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13419_ _06507_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14399_ _00253_ net3 mod.u_cpu.rf_ram.memory\[488\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _03253_ _03261_ _03262_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__14399__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11128__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07911_ _01607_ _02215_ _02217_ _02218_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__15644__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ _02479_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12876__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08544__A2 _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07842_ _01741_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07773_ mod.u_cpu.rf_ram.memory\[176\]\[0\] mod.u_cpu.rf_ram.memory\[177\]\[0\] mod.u_cpu.rf_ram.memory\[178\]\[0\]
+ mod.u_cpu.rf_ram.memory\[179\]\[0\] _02048_ _02049_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09512_ _03736_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ _03391_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13532__I _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15024__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _03496_ mod.u_scanchain_local.module_data_in\[61\] _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07530__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08325_ _01495_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ _02528_ _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__A1 _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15174__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ mod.u_cpu.raddr\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08187_ _02393_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10414__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07138_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08361__I _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13200__C _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08783__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10080_ _04162_ mod.u_cpu.rf_ram.memory\[505\]\[0\] _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12867__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13770_ _03403_ _06771_ _03377_ _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10982_ _04774_ mod.u_cpu.rf_ram.memory\[364\]\[0\] _04785_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12721_ _05588_ _05952_ _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_43_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11163__S _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15440_ _00003_ net3 mod.u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12652_ _05926_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11603_ _05209_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15371_ _01146_ net3 mod.u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15517__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12583_ _05869_ mod.u_cpu.rf_ram.memory\[157\]\[0\] _05879_ _05880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14322_ _00176_ net3 mod.u_cpu.rf_ram.memory\[526\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10653__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11534_ _03835_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11897__I _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13347__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14253_ _00107_ net3 mod.u_cpu.rf_ram.memory\[561\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11465_ _05116_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13204_ _06310_ _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14541__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08223__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _04387_ mod.u_cpu.rf_ram.memory\[456\]\[1\] _04401_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14184_ _01985_ _07086_ _07087_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11396_ _05070_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13135_ _06257_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08774__A2 mod.u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _04345_ mod.u_cpu.rf_ram.memory\[467\]\[1\] _04354_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12722__S _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13066_ _06213_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10278_ _04301_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14691__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11905__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12017_ _05494_ _05471_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08526__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08909__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15047__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12086__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13968_ mod.u_arbiter.i_wb_cpu_rdt\[4\] _06938_ _06928_ _03444_ _06939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12919_ _06101_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13899_ _01453_ _06140_ _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15638_ _01409_ net3 mod.u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__I _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15197__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15569_ _01340_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08110_ _01592_ _02402_ _02417_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09090_ _03390_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08041_ _02058_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11349__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08181__I _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08214__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09962__A1 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _04096_ mod.u_cpu.rf_ram.memory\[518\]\[0\] _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12632__S _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08943_ mod.u_cpu.rf_ram_if.rdata0\[1\] _03248_ _01478_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12849__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08517__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08874_ mod.u_cpu.rf_ram.memory\[559\]\[1\] _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07525__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07825_ _02129_ mod.u_cpu.rf_ram.memory\[164\]\[0\] _02132_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07820__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11047__I _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07756_ mod.u_cpu.rf_ram.memory\[136\]\[0\] mod.u_cpu.rf_ram.memory\[137\]\[0\] mod.u_cpu.rf_ram.memory\[138\]\[0\]
+ mod.u_cpu.rf_ram.memory\[139\]\[0\] _02022_ _02063_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14414__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07687_ _01762_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12872__I1 mod.u_cpu.rf_ram.memory\[409\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09426_ _03654_ _03658_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07260__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09357_ _03598_ _03595_ _03599_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12624__I1 mod.u_cpu.rf_ram.memory\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11588__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ mod.u_cpu.rf_ram.memory\[479\]\[1\] _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14564__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A2 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ mod.u_cpu.rf_ram.memory\[525\]\[0\] _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11250_ _04831_ _04969_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _04245_ mod.u_cpu.rf_ram.memory\[48\]\[1\] _04252_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08024__C _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09953__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__I _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11181_ _04643_ _04922_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_162_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10132_ _04193_ mod.u_cpu.rf_ram.memory\[498\]\[0\] _04203_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11158__S _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13437__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12341__I _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10063_ _04140_ mod.u_cpu.rf_ram.memory\[508\]\[1\] _04152_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14940_ _00794_ net3 mod.u_cpu.rf_ram.memory\[222\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11512__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14871_ _00725_ net3 mod.u_cpu.rf_ram.memory\[251\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13822_ _06814_ _06815_ _06817_ _06820_ _06753_ _06821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__12068__A2 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10079__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12312__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13753_ _06726_ _06472_ _06283_ _06712_ _06757_ _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10796__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _04773_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12704_ _05960_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13684_ _06367_ _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08692__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14907__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07170__I _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10896_ _04720_ mod.u_cpu.rf_ram.memory\[378\]\[1\] _04725_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15423_ _01198_ net3 mod.u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12635_ _05914_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10626__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15354_ _01129_ net3 mod.u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12566_ _05858_ mod.u_cpu.rf_ram.memory\[160\]\[1\] _05866_ _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14305_ _00159_ net3 mod.u_cpu.rf_ram.memory\[535\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11517_ _04732_ _05149_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10237__S _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15285_ _00044_ net4 mod.u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12497_ _05606_ _04309_ _05824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09097__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14236_ _00090_ net3 mod.u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11448_ _05096_ mod.u_cpu.rf_ram.memory\[290\]\[0\] _05103_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__A2 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13740__A2 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14167_ _07071_ _07075_ _07076_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11379_ _04775_ _05058_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13118_ _06237_ mod.u_cpu.rf_ram.memory\[0\]\[1\] _06245_ _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14098_ _07028_ mod.u_cpu.rf_ram.memory\[120\]\[1\] _07030_ _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13879__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13049_ _02373_ _06201_ _06202_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14437__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _01750_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08590_ _02688_ _02895_ _02896_ _01698_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07541_ _01832_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14587__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ mod.u_cpu.rf_ram.memory\[431\]\[0\] _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08176__I _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07486__A2 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09211_ _03478_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10490__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08109__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09142_ _03409_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08435__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10242__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09073_ _03371_ _03375_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ _02329_ mod.u_cpu.rf_ram.memory\[118\]\[0\] _02331_ _01916_ _02332_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__S _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13031__I1 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A2 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13731__A2 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12362__S _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15212__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09735__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _03714_ _04077_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_130_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_19 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08926_ _02525_ _03229_ _03232_ _02539_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12542__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__I1 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _02102_ _03146_ _03163_ _01739_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15362__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _01862_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08788_ mod.u_cpu.rf_ram.memory\[92\]\[1\] mod.u_cpu.rf_ram.memory\[93\]\[1\] mod.u_cpu.rf_ram.memory\[94\]\[1\]
+ mod.u_cpu.rf_ram.memory\[95\]\[1\] _01636_ _01638_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09470__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13798__A2 _06798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07739_ _02026_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10856__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10750_ _04360_ _04623_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08674__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09409_ _03561_ _03643_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _01706_ _04581_ _04582_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12420_ _05766_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12351_ _05719_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13970__A2 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12336__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11302_ _05006_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15070_ _00924_ net3 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12282_ _05673_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14021_ _06942_ _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11233_ mod.u_cpu.rf_ram.memory\[325\]\[1\] _04819_ _04956_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13722__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09777__I1 mod.u_cpu.rf_ram.memory\[550\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09645__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11164_ _04911_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__C _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13167__I _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ _04162_ mod.u_cpu.rf_ram.memory\[500\]\[0\] _04190_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11095_ _04457_ _04848_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__I1 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10046_ _04135_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14923_ _00777_ net3 mod.u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10520__S _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14854_ _00708_ net3 mod.u_cpu.rf_ram.memory\[260\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13805_ _06468_ _06452_ _06779_ _06804_ _06776_ _06805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11997_ _05019_ _05433_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14785_ _00639_ net3 mod.u_cpu.rf_ram.memory\[295\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09457__A3 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13736_ _06726_ _06459_ _06741_ _06442_ _06381_ _06742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08665__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07468__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10948_ _04762_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13667_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _06678_ _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10879_ _04698_ mod.u_cpu.rf_ram.memory\[381\]\[1\] _04714_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15406_ _01181_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12618_ _05903_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13598_ mod.u_cpu.cpu.bufreg.i_sh_signed _03669_ _03693_ _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10224__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12549_ _05857_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15337_ _01112_ net3 mod.u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15235__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15268_ _00025_ net4 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07640__A2 mod.u_cpu.rf_ram.memory\[292\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11024__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13713__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14219_ _07107_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15199_ _01052_ net3 mod.u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15385__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _03747_ _03748_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09491__S _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08711_ mod.u_cpu.rf_ram.memory\[232\]\[1\] mod.u_cpu.rf_ram.memory\[233\]\[1\] mod.u_cpu.rf_ram.memory\[234\]\[1\]
+ mod.u_cpu.rf_ram.memory\[235\]\[1\] _01647_ _01732_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09691_ _03746_ _03710_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ mod.u_cpu.rf_ram.memory\[175\]\[1\] _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07803__I _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ _01949_ _02879_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ _01444_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08656__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07455_ _01762_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08408__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13401__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _01676_ _01692_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _03415_ _03422_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09056_ _03280_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09208__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08007_ _02297_ mod.u_cpu.rf_ram.memory\[124\]\[0\] _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14602__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09465__I _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12763__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09958_ _04073_ mod.u_cpu.rf_ram.memory\[524\]\[0\] _04081_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14752__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08909_ mod.u_cpu.rf_ram.memory\[520\]\[1\] mod.u_cpu.rf_ram.memory\[521\]\[1\] mod.u_cpu.rf_ram.memory\[522\]\[1\]
+ mod.u_cpu.rf_ram.memory\[523\]\[1\] _02507_ _02543_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_44_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__A1 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ _03945_ _04034_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13715__I mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _05413_ mod.u_cpu.rf_ram.memory\[222\]\[0\] _05429_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07537__I3 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12691__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15108__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11851_ _05364_ mod.u_cpu.rf_ram.memory\[149\]\[1\] _05378_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10802_ _04662_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14570_ _00424_ net3 mod.u_cpu.rf_ram.memory\[402\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08745__S _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11782_ _05329_ mod.u_cpu.rf_ram.memory\[235\]\[1\] _05331_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13640__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10733_ _04608_ mod.u_cpu.rf_ram.memory\[404\]\[1\] _04614_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13521_ _06573_ _06574_ _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15258__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13452_ _03541_ _06525_ _06526_ _03547_ _06529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10664_ _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12403_ _05753_ mod.u_cpu.rf_ram.memory\[176\]\[0\] _05754_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13383_ _03665_ _03391_ _03672_ _06478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_182_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15122_ _00975_ net3 mod.u_cpu.rf_ram.memory\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12334_ _05696_ mod.u_cpu.rf_ram.memory\[183\]\[0\] _05707_ _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A2 _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14282__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15053_ _00907_ net3 mod.u_cpu.rf_ram.memory\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12265_ _05661_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11706__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14004_ _06962_ _06965_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11216_ _04668_ _04945_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12196_ _05614_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ mod.u_cpu.rf_ram.memory\[33\]\[1\] _04819_ _04898_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12506__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11078_ _04843_ mod.u_cpu.rf_ram.memory\[350\]\[0\] _04853_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10029_ _03986_ _04118_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14906_ _00760_ net3 mod.u_cpu.rf_ram.memory\[231\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08886__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07233__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14837_ _00691_ net3 mod.u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12809__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14768_ _00622_ net3 mod.u_cpu.rf_ram.memory\[303\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13719_ _06320_ _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11493__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14699_ _00553_ net3 mod.u_cpu.rf_ram.memory\[338\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07240_ _01545_ mod.u_cpu.rf_ram.memory\[462\]\[0\] _01547_ _01525_ _01548_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14187__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07861__A2 _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11245__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14625__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09989__I1 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07171_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11945__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13698__A1 _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08403__B _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14775__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07377__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09812_ _03978_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09743_ _03924_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12122__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09674_ _03778_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13870__A1 _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07533__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _02925_ _02927_ _02929_ _02931_ _02077_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08556_ _01915_ _02855_ _02862_ _01812_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15400__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07507_ _01739_ _01790_ _01814_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08487_ _01496_ mod.u_cpu.rf_ram.memory\[358\]\[1\] _02793_ _02453_ _02794_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13270__I _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07438_ _01568_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07852__A2 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15550__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13925__A2 _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _01550_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09108_ _03407_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10380_ _03721_ _04134_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08801__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ mod.u_cpu.cpu.decode.op26 _01452_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12050_ _05515_ _03810_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07368__A1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ _04527_ _04780_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__12361__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10911__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13161__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08868__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12952_ _06128_ _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07443__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11903_ _03984_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12883_ _06078_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07391__I1 mod.u_cpu.rf_ram.memory\[409\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14622_ _00476_ net3 mod.u_cpu.rf_ram.memory\[376\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15080__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11834_ _05367_ _05335_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14648__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14553_ _00407_ net3 mod.u_cpu.rf_ram.memory\[411\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11765_ _04377_ _05320_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09293__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15312__D _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10716_ _04593_ mod.u_cpu.rf_ram.memory\[407\]\[1\] _04603_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13504_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _06557_ _06558_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14484_ _00338_ net3 mod.u_cpu.rf_ram.memory\[445\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11696_ _05268_ mod.u_cpu.rf_ram.memory\[254\]\[0\] _05273_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13377__B1 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ _04557_ mod.u_cpu.rf_ram.memory\[418\]\[0\] _04558_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13435_ _06518_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11927__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14798__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13366_ _06326_ _06391_ _06330_ _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10578_ _04511_ _03919_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15105_ _00959_ net3 mod.u_cpu.rf_ram.memory\[174\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__S _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12317_ _05515_ _05686_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13297_ _06301_ _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12727__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12248_ _05432_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15036_ _00890_ net3 mod.u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12179_ _05602_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__C _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13355__I _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13152__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13852__A1 _06842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15423__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07353__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10666__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09520__A2 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ _01709_ _02716_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _03564_ _03625_ _03627_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_17_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ mod.u_cpu.rf_ram.memory\[511\]\[1\] _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10418__A1 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11466__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15573__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ _02545_ _02575_ _02579_ _02555_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07223_ mod.u_cpu.raddr\[3\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10219__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13907__A2 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11769__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13383__A3 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12718__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07528__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09743__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11941__I1 mod.u_cpu.rf_ram.memory\[220\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07987_ _01854_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13143__I0 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09726_ _03902_ _03911_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13843__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10657__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09657_ _03856_ _03848_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08608_ mod.u_cpu.rf_ram.memory\[128\]\[1\] mod.u_cpu.rf_ram.memory\[129\]\[1\] mod.u_cpu.rf_ram.memory\[130\]\[1\]
+ mod.u_cpu.rf_ram.memory\[131\]\[1\] _02638_ _02067_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09588_ _03739_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _01843_ _02845_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11550_ _05174_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11082__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14940__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A2 mod.u_cpu.rf_ram.memory\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10501_ _04322_ _04443_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10129__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11481_ _05107_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13220_ _06122_ _06123_ _06327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _03898_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12582__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13151_ _06266_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10363_ _04365_ mod.u_cpu.rf_ram.memory\[464\]\[0\] _04366_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12102_ _05550_ mod.u_cpu.rf_ram.memory\[67\]\[1\] _05547_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13082_ _03932_ _06223_ _06224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10294_ _04298_ mod.u_cpu.rf_ram.memory\[475\]\[0\] _04319_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08978__B mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12033_ _05505_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08002__A2 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14320__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15446__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13134__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13175__I _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07761__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13984_ _06949_ _06950_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13834__A1 _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09502__A2 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14470__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12935_ _01434_ _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11696__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15596__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11624__S _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12866_ mod.u_cpu.cpu.state.ibus_cyc _06066_ _06046_ _06067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07901__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11448__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14605_ _00459_ net3 mod.u_cpu.rf_ram.memory\[385\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11817_ _05342_ mod.u_cpu.rf_ram.memory\[230\]\[0\] _05356_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15585_ _01356_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09266__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12797_ _06010_ mod.u_cpu.rf_ram.memory\[12\]\[0\] _06021_ _06022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14536_ _00390_ net3 mod.u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11748_ _05308_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09018__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14467_ _00321_ net3 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11679_ _05261_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13418_ _06351_ mod.u_cpu.rf_ram.memory\[339\]\[0\] _06506_ _06507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09569__A2 _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14398_ _00252_ net3 mod.u_cpu.rf_ram.memory\[488\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08241__A2 mod.u_cpu.rf_ram.memory\[524\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13349_ _06422_ _06445_ _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13794__B _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07910_ _01746_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15019_ _00873_ net3 mod.u_cpu.rf_ram.memory\[206\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08890_ mod.u_cpu.rf_ram.memory\[565\]\[1\] _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12876__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07841_ _01488_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14813__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08179__I _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _01661_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09511_ mod.u_cpu.rf_ram.memory\[9\]\[1\] _03735_ _03729_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _03663_ _03666_ _03669_ _03672_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14963__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_91_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _03489_ _03611_ _03612_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08324_ _02347_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15319__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ mod.u_cpu.rf_ram.memory\[533\]\[0\] _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12365__S _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08480__A2 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ _01508_ mod.u_cpu.rf_ram.memory\[452\]\[0\] _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08186_ _01705_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_4_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07137_ _01445_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14343__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15469__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12867__A2 _06066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09473__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14493__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14069__A1 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11508__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13116__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08310__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08791__I0 mod.u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10412__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11678__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09709_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10981_ _04784_ _04759_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12720_ _03698_ _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10350__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12651_ _05918_ mod.u_cpu.rf_ram.memory\[146\]\[0\] _05925_ _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11602_ _05208_ mod.u_cpu.rf_ram.memory\[266\]\[1\] _05206_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15370_ _01145_ net3 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12582_ _05515_ _05374_ _05879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14321_ _00175_ net3 mod.u_cpu.rf_ram.memory\[527\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09263__A4 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11533_ _05163_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14252_ _00106_ net3 mod.u_cpu.rf_ram.memory\[561\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11464_ _05114_ mod.u_cpu.rf_ram.memory\[288\]\[0\] _05115_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13203_ _06118_ _06309_ _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10415_ _04402_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11602__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08223__A2 mod.u_cpu.rf_ram.memory\[516\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14183_ _07026_ _07086_ _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11395_ _05069_ mod.u_cpu.rf_ram.memory\[300\]\[1\] _05067_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09420__A1 _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10346_ _04355_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13134_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _06253_ _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14836__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07982__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13065_ _06205_ mod.u_cpu.rf_ram.memory\[106\]\[0\] _06212_ _06213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10277_ _03769_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12016_ _03827_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08082__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14986__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08909__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13967_ _06937_ _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12918_ mod.u_cpu.rf_ram.memory\[389\]\[1\] _06005_ _06099_ _06101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13898_ _01435_ _06881_ _06847_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15637_ _01408_ net3 mod.u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12849_ _02523_ _03742_ _06054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15568_ _01339_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13991__B1 _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14519_ _00373_ net3 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10992__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15499_ _01270_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14366__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13301__C _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15611__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13594__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08214__A2 _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09411__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08845__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09962__A2 _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09991_ _03951_ _04087_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07973__A1 _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08942_ _03247_ mod.u_cpu.rf_ram.regzero _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12712__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08873_ _02478_ mod.u_cpu.rf_ram.memory\[556\]\[1\] _03179_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07725__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07824_ _02130_ _02131_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07820__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09478__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ _01960_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11264__S _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07686_ _01993_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07541__I _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15141__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09425_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] _03561_ _03656_ _03657_ _03409_ _03658_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14709__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13699__B _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09356_ _03598_ _03586_ _03594_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08307_ _02566_ mod.u_cpu.rf_ram.memory\[476\]\[1\] _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09287_ _03528_ _03539_ _03540_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__S _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _02477_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15291__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12537__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14859__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08169_ _02047_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__S0 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10200_ _04253_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09953__A2 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11180_ _04379_ _04779_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _04201_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10062_ _04153_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11899__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07716__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11512__A2 _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14870_ _00724_ net3 mod.u_cpu.rf_ram.memory\[251\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13821_ _06818_ _06819_ _06332_ _06820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14239__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13752_ _06666_ _06671_ _06756_ _06757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10964_ _04772_ mod.u_cpu.rf_ram.memory\[367\]\[1\] _04770_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07451__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12703_ mod.u_cpu.rf_ram.memory\[13\]\[0\] _05622_ _05959_ _05960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13683_ _06482_ _06475_ _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08692__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _04726_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14389__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15422_ _01197_ net3 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11028__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12634_ _05907_ mod.u_cpu.rf_ram.memory\[14\]\[1\] _05912_ _05914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15634__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12776__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10626__I1 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15353_ _01128_ net3 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12565_ _05867_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14304_ _00158_ net3 mod.u_cpu.rf_ram.memory\[535\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _05152_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15284_ _00043_ net4 mod.u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12496_ _05823_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13576__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14235_ _00089_ net3 mod.u_cpu.rf_ram.memory\[570\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10317__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11447_ _04831_ _05089_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11378_ _04995_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14166_ _06046_ _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13740__A3 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07955__A1 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13628__I _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10329_ _04326_ mod.u_cpu.rf_ram.memory\[46\]\[0\] _04342_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13117_ _06246_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14097_ _07031_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15014__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13879__I1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07626__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13048_ _06032_ _06201_ _06202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09841__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15164__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13363__I _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14999_ _00853_ net3 mod.u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07540_ _01457_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08457__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08132__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07361__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07471_ _01778_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14205__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09210_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] _03474_
+ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _03409_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12707__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09632__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10242__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08192__I _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09072_ _03374_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08023_ _01863_ _02330_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04092_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07536__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08925_ _02533_ mod.u_cpu.rf_ram.memory\[542\]\[1\] _03231_ _02537_ _03232_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15507__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11058__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12542__I1 mod.u_cpu.rf_ram.memory\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03151_ _03153_ _03162_ _01891_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08371__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08795__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _01635_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08787_ _01662_ _03093_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13273__I _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14531__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07738_ _01890_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08674__A2 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07669_ _01484_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09408_ _03642_ _03638_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10680_ _04542_ _04581_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14681__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10608__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09339_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12350_ _05711_ mod.u_cpu.rf_ram.memory\[181\]\[1\] _05717_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13707__B1 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11301_ _04999_ mod.u_cpu.rf_ram.memory\[315\]\[1\] _05004_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13558__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12281_ _05662_ mod.u_cpu.rf_ram.memory\[190\]\[0\] _05672_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15037__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14020_ _06975_ _06977_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13183__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _04957_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11169__S _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _04901_ mod.u_cpu.rf_ram.memory\[336\]\[0\] _04910_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12352__I _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10114_ _04189_ _04164_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11094_ _04802_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15187__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10045_ _04141_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14922_ _00776_ net3 mod.u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14853_ _00707_ net3 mod.u_cpu.rf_ram.memory\[261\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08752__I3 mod.u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13804_ _06803_ _06714_ _06804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14784_ _00638_ net3 mod.u_cpu.rf_ram.memory\[295\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11996_ _05480_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07181__I _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__I0 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12997__A1 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13735_ _06739_ _03424_ _06740_ _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12997__B2 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10947_ _04756_ mod.u_cpu.rf_ram.memory\[370\]\[1\] _04760_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__A2 _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13666_ _06415_ _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10878_ _01859_ _04714_ _04715_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12749__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15405_ _01180_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12617_ _05891_ mod.u_cpu.rf_ram.memory\[152\]\[1\] _05901_ _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09614__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13597_ _03659_ _03694_ _06619_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15336_ _01111_ net3 mod.u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12548_ _05855_ mod.u_cpu.rf_ram.memory\[163\]\[0\] _05856_ _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10047__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15267_ _00024_ net4 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09217__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12479_ _05694_ _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14210__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11024__I1 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14218_ _03699_ mod.u_cpu.rf_ram.memory\[249\]\[0\] _07106_ _07107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15198_ _01051_ net3 mod.u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14404__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07928__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14149_ _03822_ _05254_ _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07356__I _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08710_ _01991_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11488__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09690_ _03882_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14554__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08641_ _02111_ mod.u_cpu.rf_ram.memory\[172\]\[1\] _02947_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08187__I _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08572_ mod.u_cpu.rf_ram.memory\[279\]\[1\] _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07523_ mod.u_cpu.rf_ram.memory\[344\]\[0\] mod.u_cpu.rf_ram.memory\[345\]\[0\] mod.u_cpu.rf_ram.memory\[346\]\[0\]
+ mod.u_cpu.rf_ram.memory\[347\]\[0\] _01826_ _01830_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ _01700_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07385_ _01445_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13401__A2 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09124_ _03392_ _03420_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _03354_ _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08006_ _02298_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07919__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _03905_ _04062_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ _02449_ _03207_ _03214_ _02469_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09888_ _03823_ _04033_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08344__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08839_ _03142_ _03143_ _03144_ _03145_ _02391_ _01552_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_72_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08895__A2 mod.u_cpu.rf_ram.memory\[566\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _05379_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08097__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12979__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10801_ mod.u_cpu.rf_ram.memory\[393\]\[1\] _04661_ _04659_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12548__S _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11781_ _05332_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13640__A2 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13520_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _03669_ _06574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10732_ _04615_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13451_ _06528_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10663_ _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12402_ _05300_ _05726_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11403__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10594_ _04247_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13382_ _06457_ _06460_ _06477_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14427__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15121_ _00974_ net3 mod.u_cpu.rf_ram.memory\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12333_ _03879_ _05703_ _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15052_ _00906_ net3 mod.u_cpu.rf_ram.memory\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12264_ _05660_ mod.u_cpu.rf_ram.memory\[193\]\[1\] _05658_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14003_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _06964_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11706__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11215_ _04905_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12195_ _05609_ mod.u_cpu.rf_ram.memory\[202\]\[1\] _05612_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14577__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08583__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11146_ _04899_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11077_ _04852_ _04848_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08335__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _04128_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14905_ _00759_ net3 mod.u_cpu.rf_ram.memory\[232\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10142__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14836_ _00690_ net3 mod.u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14767_ _00621_ net3 mod.u_cpu.rf_ram.memory\[304\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09835__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11979_ _05469_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13631__A2 _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13718_ _06723_ _06123_ _06724_ _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15202__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11642__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14698_ _00552_ net3 mod.u_cpu.rf_ram.memory\[338\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13919__B1 _06896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13649_ _06404_ _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13395__A1 _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07170_ _01449_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15352__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15319_ _01098_ net3 mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11945__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08403__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07377__A2 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09811_ _03964_ mod.u_cpu.rf_ram.memory\[546\]\[1\] _03976_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12720__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _03923_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10508__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07814__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12122__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09673_ _03869_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _02074_ _02930_ _01602_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08555_ _01981_ _02858_ _02861_ _01929_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13551__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07506_ _01791_ _01800_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08486_ _02672_ _02792_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07437_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _01658_ _01668_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ _03405_ _03406_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07299_ _01539_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08801__A2 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08380__I _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ mod.u_cpu.cpu.decode.op22 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13689__A2 _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07368__A2 _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11000_ _04798_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12361__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13310__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12951_ _06126_ _03424_ _06127_ _06128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10150__I _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11902_ _05416_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15225__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12882_ _06073_ mod.u_cpu.rf_ram.memory\[99\]\[0\] _06077_ _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14621_ _00475_ net3 mod.u_cpu.rf_ram.memory\[377\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11833_ _03959_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11182__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14552_ _00406_ net3 mod.u_cpu.rf_ram.memory\[411\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _04227_ _05319_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13503_ _06560_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10715_ _01730_ _04603_ _04604_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15375__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14483_ _00337_ net3 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11695_ _04852_ _05255_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13377__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13377__B2 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13434_ _03507_ _06511_ _06514_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _06518_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10646_ _04281_ _04534_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11927__A2 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13365_ _03664_ _03663_ _06356_ _06461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10577_ _04250_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15104_ _00958_ net3 mod.u_cpu.rf_ram.memory\[174\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__I _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12316_ _05695_ _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13296_ _06313_ _06393_ _06389_ _06394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15035_ _00889_ net3 mod.u_cpu.rf_ram.memory\[200\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12727__I1 mod.u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12741__S _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12247_ _03967_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__10738__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12178_ _05575_ mod.u_cpu.rf_ram.memory\[204\]\[0\] _05601_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13636__I _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11129_ _04883_ mod.u_cpu.rf_ram.memory\[342\]\[0\] _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08859__A2 _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11163__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13572__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08666__S _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11863__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14101__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14819_ _00673_ net3 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09808__A1 _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11092__S _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10418__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08340_ _02559_ mod.u_cpu.rf_ram.memory\[508\]\[1\] _02646_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11466__I1 mod.u_cpu.rf_ram.memory\[288\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _02550_ mod.u_cpu.rf_ram.memory\[542\]\[0\] _02577_ _02578_ _02579_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07222_ _01505_ _01514_ _01526_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14742__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09036__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08795__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08133__C _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14892__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10235__I _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15248__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07986_ _01864_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09725_ _03910_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11066__I _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10657__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09656_ _03744_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14272__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _01481_ _02758_ _02913_ _01469_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15398__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09587_ _03801_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ mod.u_cpu.rf_ram.memory\[293\]\[1\] _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11082__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _01852_ _02768_ _02775_ _01887_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10500_ _04460_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11480_ _05127_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _04412_ _04380_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13150_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _06263_ _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10362_ _04209_ _04353_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12101_ _05549_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10293_ _03791_ _04303_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13081_ _05630_ _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09586__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12032_ _05501_ mod.u_cpu.rf_ram.memory\[19\]\[1\] _05503_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13456__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12360__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07454__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13134__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07761__A2 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13983_ mod.u_arbiter.i_wb_cpu_rdt\[8\] _06938_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14615__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12934_ mod.u_cpu.cpu.genblk3.csr.mie_mtie mod.u_cpu.cpu.genblk3.csr.mstatus_mie
+ mod.timer_irq _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11696__I1 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12893__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12865_ _06063_ _06065_ _06066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13598__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14604_ _00458_ net3 mod.u_cpu.rf_ram.memory\[385\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08285__I _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11816_ _05355_ _05335_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15584_ _01355_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14765__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12796_ _05870_ _03905_ _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07277__A1 _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14535_ _00389_ net3 mod.u_cpu.rf_ram.memory\[420\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11747_ _05304_ mod.u_cpu.rf_ram.memory\[23\]\[1\] _05306_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14466_ _00320_ net3 mod.u_cpu.rf_ram.memory\[454\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11678_ _05250_ mod.u_cpu.rf_ram.memory\[256\]\[1\] _05259_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13417_ _05732_ _04847_ _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10256__S _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _04547_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13070__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14397_ _00251_ net3 mod.u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08777__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13770__A1 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13348_ _06433_ _06440_ _06444_ _06401_ _06445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10584__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13279_ _06116_ _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08529__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09577__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15018_ _00872_ net3 mod.u_cpu.rf_ram.memory\[206\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07840_ _01482_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07364__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14295__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07771_ _02039_ _02062_ _02078_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_68_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15540__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09510_ _03734_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12884__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08701__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _03670_ _03403_ _03671_ _03252_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_65_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09372_ _03563_ mod.u_scanchain_local.module_data_in\[60\] _03517_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\]
+ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_80_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07268__A1 _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ _02039_ _02608_ _02629_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08254_ mod.u_cpu.rf_ram.memory\[528\]\[0\] mod.u_cpu.rf_ram.memory\[529\]\[0\] mod.u_cpu.rf_ram.memory\[530\]\[0\]
+ mod.u_cpu.rf_ram.memory\[531\]\[0\] _02560_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07967__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07205_ _01511_ _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08185_ _02470_ _02492_ _01447_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08768__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09955__S _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13761__A1 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07136_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15070__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14638__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07274__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14069__A2 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07969_ _01742_ _02268_ _02276_ _02207_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09708_ _03697_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11827__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14788__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10980_ _03903_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09639_ _03842_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _05293_ _05920_ _05925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12627__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11601_ _05177_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12581_ _05878_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10102__I1 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14320_ _00174_ net3 mod.u_cpu.rf_ram.memory\[527\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11532_ _05162_ mod.u_cpu.rf_ram.memory\[278\]\[1\] _05160_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14251_ _00105_ net3 mod.u_cpu.rf_ram.memory\[562\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12004__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11463_ _04838_ _04996_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__B _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13202_ _06308_ _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07449__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08759__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13752__A1 _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15413__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10414_ _04400_ mod.u_cpu.rf_ram.memory\[456\]\[0\] _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14182_ _03822_ _05124_ _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10566__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _05031_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13133_ _06256_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10345_ _04348_ mod.u_cpu.rf_ram.memory\[467\]\[0\] _04354_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13064_ _03918_ _06092_ _06212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _04306_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10318__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13186__I _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11366__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15563__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12015_ _05493_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07184__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08931__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13966_ _05801_ _06937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12917_ _06100_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12491__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13897_ _03342_ _06881_ _06856_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12848_ _06052_ _06053_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15636_ _01407_ net3 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15567_ _01338_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12779_ _05998_ mod.u_cpu.rf_ram.memory\[132\]\[1\] _06007_ _06009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13991__A1 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14518_ _00372_ net3 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15498_ _01269_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14449_ _00303_ net3 mod.u_cpu.rf_ram.memory\[463\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15093__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13743__A1 _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13594__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09411__A2 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08845__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _04102_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08941_ mod.u_cpu.rf_ram.rdata\[0\] _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11357__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08411__C _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10513__I _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _02479_ _03178_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08922__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14930__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__A2 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07823_ mod.u_cpu.rf_ram.memory\[165\]\[0\] _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07754_ _02045_ _02052_ _02056_ _02061_ _01818_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_53_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09478__A2 _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07489__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07685_ _01645_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07584__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09424_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _03648_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _03637_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__12609__I0 _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09355_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12234__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14310__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _02593_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08989__A1 _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15436__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09286_ _03535_ mod.u_scanchain_local.module_data_in\[46\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09650__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08237_ _02325_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07661__A1 _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07269__I _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13585__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08168_ _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08836__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14460__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11596__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15586__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07119_ mod.u_cpu.cpu.decode.co_mem_word _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07413__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08099_ mod.u_cpu.rf_ram.memory\[21\]\[0\] _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10130_ _04142_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _04148_ mod.u_cpu.rf_ram.memory\[508\]\[0\] _04152_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10423__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13820_ _06311_ _06458_ _06466_ _06372_ _06776_ _06819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07732__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13751_ _06323_ _06425_ _06326_ _06281_ _06330_ _06756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10963_ _04719_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11520__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12702_ _03728_ _04643_ _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13682_ _06692_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _04695_ mod.u_cpu.rf_ram.memory\[378\]\[0\] _04725_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15421_ _01196_ net3 mod.u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12633_ _05913_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11028__A2 _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12286__S _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__S _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09659__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15352_ _01127_ net3 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12776__A2 _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12564_ _05855_ mod.u_cpu.rf_ram.memory\[160\]\[0\] _05866_ _05867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14303_ _00157_ net3 mod.u_cpu.rf_ram.memory\[536\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _05147_ mod.u_cpu.rf_ram.memory\[281\]\[1\] _05150_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12085__I _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14803__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15283_ _00042_ net4 mod.u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12495_ _05822_ mod.u_cpu.rf_ram.memory\[170\]\[1\] _05820_ _05823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14234_ _00088_ net3 mod.u_cpu.rf_ram.memory\[570\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13725__B2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11446_ _05102_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14165_ _03670_ _07072_ _07074_ _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12813__I _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _05057_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14953__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13116_ _06230_ mod.u_cpu.rf_ram.memory\[0\]\[0\] _06245_ _06246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10328_ _04251_ _03886_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14096_ _07021_ mod.u_cpu.rf_ram.memory\[120\]\[0\] _07030_ _07031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09157__A1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14150__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13047_ _04067_ _05387_ _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10259_ _04293_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15309__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13644__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14998_ _00852_ net3 mod.u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12464__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13949_ _03438_ _06917_ _06919_ _06922_ _06923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08132__A2 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14333__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ _01757_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15459__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15619_ _01390_ net3 mod.u_cpu.rf_ram.memory\[247\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09140_ _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09632__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14483__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09071_ _03372_ _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08022_ mod.u_cpu.rf_ram.memory\[119\]\[0\] _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13567__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ _04091_ mod.u_cpu.rf_ram.memory\[522\]\[1\] _04088_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11339__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08924_ _02534_ _03230_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09943__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08855_ _03017_ _03154_ _03161_ _02852_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _02111_ mod.u_cpu.rf_ram.memory\[172\]\[0\] _02113_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08371__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08786_ mod.u_cpu.rf_ram.memory\[88\]\[1\] mod.u_cpu.rf_ram.memory\[89\]\[1\] mod.u_cpu.rf_ram.memory\[90\]\[1\]
+ mod.u_cpu.rf_ram.memory\[91\]\[1\] _01673_ _01855_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07737_ _02040_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07668_ _01739_ _01944_ _01975_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14826__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _01663_ _01906_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15421__D _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _03583_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07634__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09269_ _03524_ _03525_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__13707__A1 _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11300_ _05005_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14976__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13558__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12280_ _05428_ _05668_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13183__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11231_ mod.u_cpu.rf_ram.memory\[325\]\[0\] _04954_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ _04766_ _04906_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11249__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10153__I _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ _03842_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14132__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11093_ _04863_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09942__I _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10044_ _04140_ mod.u_cpu.rf_ram.memory\[511\]\[1\] _04138_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14921_ _00775_ net3 mod.u_cpu.rf_ram.memory\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14356__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14852_ _00706_ net3 mod.u_cpu.rf_ram.memory\[261\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15601__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07462__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13803_ _06424_ _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07960__I2 mod.u_cpu.rf_ram.memory\[250\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14783_ _00637_ net3 mod.u_cpu.rf_ram.memory\[296\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11995_ _05464_ mod.u_cpu.rf_ram.memory\[569\]\[1\] _05478_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13734_ _06723_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _06740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12997__A2 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10946_ _04761_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14199__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13665_ _06338_ _06659_ _06665_ _06676_ _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_189_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10877_ _04611_ _04714_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15404_ _01179_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12616_ _05902_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13596_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] _03694_ _06619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09614__A2 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15335_ _01110_ net3 mod.u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _05649_ _05831_ _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11421__A2 _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15266_ _00023_ net4 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12478_ _05811_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14217_ _04025_ _05263_ _07106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10264__S _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _05087_ mod.u_cpu.rf_ram.memory\[294\]\[1\] _05090_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15197_ _01050_ net3 mod.u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14148_ _07063_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08050__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07484__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09057__C _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15131__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14079_ _07019_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08896__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10998__I _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08640_ _02130_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15281__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07372__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12437__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08571_ _01962_ mod.u_cpu.rf_ram.memory\[276\]\[1\] _02877_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14849__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07522_ _01820_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07453_ _01759_ _01760_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11622__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14999__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07384_ _01678_ _01685_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11799__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09123_ _03362_ _03385_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09054_ _03356_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14229__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08005_ mod.u_cpu.rf_ram.memory\[125\]\[0\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09369__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08416__I0 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12212__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09963__S _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__A2 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11069__I _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10923__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09956_ _04080_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14379__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__S _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15624__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08907_ _02525_ _03210_ _03213_ _02467_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09887_ _03995_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11723__I0 _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ mod.u_cpu.rf_ram.memory\[56\]\[1\] mod.u_cpu.rf_ram.memory\[57\]\[1\] mod.u_cpu.rf_ram.memory\[58\]\[1\]
+ mod.u_cpu.rf_ram.memory\[59\]\[1\] _02242_ _02388_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12428__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _02283_ _03072_ _03075_ _02308_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _04531_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11780_ _05311_ mod.u_cpu.rf_ram.memory\[235\]\[0\] _05331_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__A2 _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10731_ _04598_ mod.u_cpu.rf_ram.memory\[404\]\[0\] _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07855__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15004__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13450_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _06525_ _06526_ _03541_ _06528_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10662_ _03993_ _04132_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12401_ _05695_ _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13381_ _06413_ _06461_ _06474_ _06476_ _06477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11403__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ _04521_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15120_ _00973_ net3 mod.u_cpu.rf_ram.memory\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09937__I _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12332_ _05706_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15154__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15051_ _00905_ net3 mod.u_cpu.rf_ram.memory\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12263_ _05634_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14002_ _06963_ _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07457__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11214_ _04944_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12194_ _05613_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14105__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ mod.u_cpu.rf_ram.memory\[33\]\[0\] _04658_ _04898_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11076_ _03750_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10517__I1 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11714__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ mod.u_cpu.rf_ram.memory\[513\]\[1\] _04111_ _04126_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14904_ _00758_ net3 mod.u_cpu.rf_ram.memory\[232\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07192__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10142__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__I1 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14835_ _00689_ net3 mod.u_cpu.rf_ram.memory\[270\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11643__S _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11978_ mod.u_cpu.rf_ram.memory\[549\]\[1\] _05468_ _05466_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14766_ _00620_ net3 mod.u_cpu.rf_ram.memory\[304\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09835__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13717_ _06723_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _06724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10929_ _03841_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14697_ _00551_ net3 mod.u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11642__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13919__A1 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13919__B2 _06897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13648_ _06289_ _06313_ _06361_ _06393_ _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13395__A2 _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13579_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] mod.u_arbiter.i_wb_cpu_dbus_adr\[23\]
+ _06609_ _06610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08271__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15318_ _01097_ net3 mod.u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13369__I _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12273__I _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15249_ _00074_ net4 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14521__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _03977_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__A2 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__B _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09741_ _03696_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14671__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09523__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _03862_ mod.u_cpu.rf_ram.memory\[561\]\[1\] _03867_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09523__B2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08623_ mod.u_cpu.rf_ram.memory\[156\]\[1\] mod.u_cpu.rf_ram.memory\[157\]\[1\] mod.u_cpu.rf_ram.memory\[158\]\[1\]
+ mod.u_cpu.rf_ram.memory\[159\]\[1\] _01925_ _02071_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15027__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _01938_ mod.u_cpu.rf_ram.memory\[318\]\[1\] _02860_ _01952_ _02861_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12130__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _01770_ _01801_ _01811_ _01812_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07837__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ mod.u_cpu.rf_ram.memory\[359\]\[1\] _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12830__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07436_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15177__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07367_ _01670_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09757__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _03398_ mod.u_cpu.cpu.state.ibus_cyc _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07298_ mod.u_cpu.rf_ram.memory\[504\]\[0\] mod.u_cpu.rf_ram.memory\[505\]\[0\] mod.u_cpu.rf_ram.memory\[506\]\[0\]
+ mod.u_cpu.rf_ram.memory\[507\]\[0\] _01605_ _01570_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_164_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13279__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12183__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09037_ _03337_ _03339_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08014__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09939_ _04033_ _04068_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11527__I _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12950_ _06116_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _06127_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13310__A2 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11901_ _05406_ mod.u_cpu.rf_ram.memory\[225\]\[1\] _05414_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12881_ _03968_ _06048_ _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14620_ _00474_ net3 mod.u_cpu.rf_ram.memory\[377\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11832_ _05310_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07740__I _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14551_ _00405_ net3 mod.u_cpu.rf_ram.memory\[412\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _05252_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11262__I _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13502_ _03648_ _06557_ _06558_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _06560_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10714_ _04542_ _04603_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14482_ _00336_ net3 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13898__B _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11694_ _05272_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13377__A2 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13433_ _06517_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10645_ _04522_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14544__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13364_ _06422_ _06459_ _06460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10576_ _04510_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10060__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15103_ _00957_ net3 mod.u_cpu.rf_ram.memory\[489\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12315_ _05694_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14225__D _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10606__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13295_ _06392_ _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15034_ _00888_ net3 mod.u_cpu.rf_ram.memory\[200\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12246_ _05648_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14694__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__A2 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12177_ _05325_ _05568_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11128_ _04741_ _04887_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11059_ _04838_ _04704_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11863__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14101__I1 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14818_ _00672_ net3 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07382__I3 mod.u_cpu.rf_ram.memory\[399\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09808__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07650__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14749_ _00603_ net3 mod.u_cpu.rf_ram.memory\[313\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12812__A1 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09284__A3 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _02139_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07221_ _01528_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07152_ _01460_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08795__A2 _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09744__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12731__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11551__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07985_ _01669_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09724_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14417__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ _03757_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08606_ _01470_ _02836_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09586_ _03800_ mod.u_cpu.rf_ram.memory\[570\]\[1\] _03798_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ mod.u_cpu.rf_ram.memory\[288\]\[1\] mod.u_cpu.rf_ram.memory\[289\]\[1\] mod.u_cpu.rf_ram.memory\[290\]\[1\]
+ mod.u_cpu.rf_ram.memory\[291\]\[1\] _01826_ _02164_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14567__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08483__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _01855_ _02771_ _02774_ _01631_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _01705_ mod.u_cpu.rf_ram.memory\[404\]\[0\] _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_168_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08399_ mod.u_cpu.rf_ram.memory\[439\]\[1\] _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13603__I0 mod.u_cpu.rf_ram.memory\[329\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10430_ _04106_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_195_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10361_ _04347_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12100_ _05404_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13080_ _06222_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10292_ _04318_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12031_ _05504_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12641__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07735__I _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] _06943_ _06949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11145__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _06062_ _03669_ _06111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12289__S _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15342__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13047__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12864_ _06064_ _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07470__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14603_ _00457_ net3 mod.u_cpu.rf_ram.memory\[386\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13598__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11815_ _03949_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15583_ _01354_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12795_ _06020_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14534_ _00388_ net3 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08474__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15492__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11746_ _02412_ _05306_ _05307_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_159_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14465_ _00319_ net3 mod.u_cpu.rf_ram.memory\[455\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11677_ _05260_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10408__I0 mod.u_cpu.rf_ram.memory\[457\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10628_ _04537_ mod.u_cpu.rf_ram.memory\[422\]\[1\] _04545_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13416_ _06505_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14396_ _00250_ net3 mod.u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10336__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13347_ _06442_ _06314_ _06443_ _06382_ _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__A2 mod.u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10559_ _04499_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _06306_ _06364_ _06370_ _06372_ _06375_ _06376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15017_ _00871_ net3 mod.u_cpu.rf_ram.memory\[207\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12229_ _05226_ _05594_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_170_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11167__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ _02065_ _02069_ _02073_ _02076_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09860__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12884__I1 mod.u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _03395_ _03331_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14086__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07380__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09371_ _03610_ _03608_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_75_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10647__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08322_ _02609_ _02619_ _02628_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07268__A2 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10272__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08253_ _02107_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09009__A3 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07204_ mod.u_cpu.rf_ram.memory\[453\]\[0\] _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08184_ _02471_ _02474_ _02490_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10024__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _01419_ _01443_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11072__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08768__A2 mod.u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15215__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11772__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08076__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15365__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13277__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07968_ _02174_ _02271_ _02275_ _01766_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08587__S _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09707_ _03893_ _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11827__A2 _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07899_ _01787_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13292__I _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10886__I0 _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09638_ _03841_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08319__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ _03700_ _03743_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11600_ _05207_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12580_ _05874_ mod.u_cpu.rf_ram.memory\[158\]\[1\] _05876_ _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08456__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10263__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11531_ _05107_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14250_ _00104_ net3 mod.u_cpu.rf_ram.memory\[562\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11462_ _05045_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12004__A2 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13201_ _06302_ _06303_ _06308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_165_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _04255_ _04373_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11063__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08054__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__S1 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14181_ _07085_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11393_ _05068_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09945__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13132_ mod.u_arbiter.i_wb_cpu_rdt\[18\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _06253_ _06256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10344_ _04352_ _04353_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11188__S _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13467__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13063_ _06211_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10275_ _04288_ mod.u_cpu.rf_ram.memory\[478\]\[1\] _04304_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10318__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ _05484_ mod.u_cpu.rf_ram.memory\[57\]\[1\] _05491_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10820__S _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14732__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13965_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _06917_ _06918_ _06935_ _06936_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12916_ mod.u_cpu.rf_ram.memory\[389\]\[0\] _05971_ _06099_ _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12491__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13896_ _06884_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15635_ _01406_ net3 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14882__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12847_ _02080_ _03742_ _06053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11651__S _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08447__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15566_ _01337_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12778_ _06008_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14517_ _00371_ net3 mod.u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13991__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12546__I _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11729_ _05287_ mod.u_cpu.rf_ram.memory\[242\]\[1\] _05294_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11450__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15497_ _01268_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15238__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14448_ _00302_ net3 mod.u_cpu.rf_ram.memory\[463\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12990__B _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13743__A2 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14379_ _00233_ net3 mod.u_cpu.rf_ram.memory\[498\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10801__I0 mod.u_cpu.rf_ram.memory\[393\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14262__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15388__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11098__S _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _01466_ _02914_ _03167_ _03246_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ mod.u_cpu.rf_ram.memory\[557\]\[1\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07308__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07822_ _01744_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13259__A1 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09590__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12306__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07753_ _02057_ _02060_ _01632_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14001__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09423_ _03564_ _03655_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _03597_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12234__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ mod.u_cpu.rf_ram.memory\[477\]\[1\] _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13982__A2 _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09285_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07110__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11360__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08236_ mod.u_cpu.rf_ram.memory\[520\]\[0\] mod.u_cpu.rf_ram.memory\[521\]\[0\] mod.u_cpu.rf_ram.memory\[522\]\[0\]
+ mod.u_cpu.rf_ram.memory\[523\]\[0\] _02507_ _02543_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14605__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13734__A2 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _01702_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11745__A1 _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07118_ mod.u_cpu.cpu.decode.op21 _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07413__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ _01644_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12191__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14755__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10060_ _03782_ _04143_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13750_ _03510_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _06754_ _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08677__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10962_ _01897_ _04770_ _04771_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13670__A1 _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12701_ _05958_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13681_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _06691_ _06658_ _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10893_ _04322_ _04709_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15420_ _01195_ net3 mod.u_cpu.rf_ram.memory\[349\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08429__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12632_ _05904_ mod.u_cpu.rf_ram.memory\[14\]\[0\] _05912_ _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13422__A1 _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10236__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12563_ _05417_ _05757_ _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15351_ _01126_ net3 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11270__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14302_ _00156_ net3 mod.u_cpu.rf_ram.memory\[536\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11514_ _05151_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12494_ _05806_ _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15282_ _00040_ net4 mod.u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14285__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14233_ _00087_ net3 mod.u_cpu.rf_ram.memory\[571\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15530__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11445_ _05087_ mod.u_cpu.rf_ram.memory\[291\]\[1\] _05100_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08288__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10815__S _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12784__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14164_ _03298_ _07073_ _07074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11376_ _05050_ mod.u_cpu.rf_ram.memory\[303\]\[1\] _05055_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08601__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10327_ _04341_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10614__I _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13115_ _06181_ _03986_ _06245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14095_ _03804_ _07014_ _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07195__I _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09157__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13046_ _06200_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10258_ _04288_ mod.u_cpu.rf_ram.memory\[480\]\[1\] _04291_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07168__A1 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07263__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _04244_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14997_ _00851_ net3 mod.u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08668__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13948_ _06920_ _06921_ _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13879_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_arbiter.i_wb_cpu_rdt\[8\] _06334_
+ _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15060__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15618_ _01389_ net3 mod.u_cpu.rf_ram.memory\[247\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14628__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15549_ _01320_ net3 mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11975__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09070_ _01434_ _01436_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08691__I1 mod.u_cpu.rf_ram.memory\[201\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14213__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08021_ _02134_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09585__I _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__B _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14778__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08422__C _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09972_ _04090_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12940__S _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08923_ mod.u_cpu.rf_ram.memory\[543\]\[1\] _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07159__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08854_ _02063_ _03157_ _03160_ _01695_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07805_ _01673_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _01696_ _03091_ _01720_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07736_ mod.u_cpu.rf_ram.memory\[128\]\[0\] mod.u_cpu.rf_ram.memory\[129\]\[0\] mod.u_cpu.rf_ram.memory\[130\]\[0\]
+ mod.u_cpu.rf_ram.memory\[131\]\[0\] _02041_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15403__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07667_ _01740_ _01955_ _01974_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_164_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09406_ _03623_ _03640_ _03641_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13404__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ mod.u_cpu.rf_ram.memory\[359\]\[0\] _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15553__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09337_ _03582_ _03579_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _03520_ _03521_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_127_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08219_ _02526_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11018__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ mod.u_arbiter.i_wb_cpu_rdt\[25\] mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] _03469_
+ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12766__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11230_ _04955_ _04922_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_49_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12391__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _04909_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07493__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12518__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10112_ _04188_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11092_ _04862_ mod.u_cpu.rf_ram.memory\[348\]\[1\] _04860_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11466__S _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10043_ _04090_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14920_ _00774_ net3 mod.u_cpu.rf_ram.memory\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09444__B _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08442__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07743__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14851_ _00705_ net3 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07570__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13802_ _06418_ _06466_ _06666_ _06443_ _06486_ _06802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_17_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15083__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13643__A1 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14782_ _00636_ net3 mod.u_cpu.rf_ram.memory\[296\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11994_ _05479_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13733_ _06723_ _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10945_ _04753_ mod.u_cpu.rf_ram.memory\[370\]\[0\] _04760_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13664_ _06672_ _06674_ _06675_ _06472_ _06134_ _06676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_10876_ _04307_ _04713_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10209__A1 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15403_ _01178_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11257__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12615_ _05887_ mod.u_cpu.rf_ram.memory\[152\]\[0\] _05901_ _05902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13595_ _06618_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15334_ _01109_ net3 mod.u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12546_ _05812_ _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14920__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15265_ _00022_ net4 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12477_ _05807_ mod.u_cpu.rf_ram.memory\[519\]\[1\] _05809_ _05811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12757__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14216_ _07105_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11428_ _05091_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15196_ _01049_ net3 mod.u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14147_ _07055_ mod.u_cpu.rf_ram.memory\[90\]\[1\] _07061_ _07063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11359_ _04959_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07484__S1 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14078_ _06578_ mod.u_cpu.rf_ram.memory\[299\]\[0\] _07018_ _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12134__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13029_ _06189_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14300__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15426__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07653__I _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09550__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07561__A1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08570_ _01963_ _02876_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09689__I0 _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12437__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10448__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07521_ mod.u_cpu.rf_ram.memory\[328\]\[0\] mod.u_cpu.rf_ram.memory\[329\]\[0\] mod.u_cpu.rf_ram.memory\[330\]\[0\]
+ mod.u_cpu.rf_ram.memory\[331\]\[0\] _01826_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__15576__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14450__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11903__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07452_ mod.u_cpu.rf_ram.memory\[423\]\[0\] _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07383_ _01688_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09122_ _03363_ _03416_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09053_ _03308_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07828__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08004_ mod.u_cpu.rf_ram.memory\[120\]\[0\] mod.u_cpu.rf_ram.memory\[121\]\[0\] mod.u_cpu.rf_ram.memory\[122\]\[0\]
+ mod.u_cpu.rf_ram.memory\[123\]\[0\] _02294_ _02295_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08416__I1 mod.u_cpu.rf_ram.memory\[409\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__I _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ mod.u_cpu.rf_ram.memory\[525\]\[1\] _03929_ _04078_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13322__B1 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _02533_ mod.u_cpu.rf_ram.memory\[518\]\[1\] _03212_ _02537_ _03213_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09886_ _04032_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08837_ mod.u_cpu.rf_ram.memory\[60\]\[1\] mod.u_cpu.rf_ram.memory\[61\]\[1\] mod.u_cpu.rf_ram.memory\[62\]\[1\]
+ mod.u_cpu.rf_ram.memory\[63\]\[1\] _02406_ _02218_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_18_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07552__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08768_ _02316_ mod.u_cpu.rf_ram.memory\[126\]\[1\] _03074_ _02306_ _03075_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _02026_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13514__B _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08699_ _02190_ _03005_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10730_ _04189_ _04599_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14943__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07855__A2 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11239__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10661_ _04567_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12400_ _05752_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13380_ _06139_ _06475_ _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10592_ _04514_ mod.u_cpu.rf_ram.memory\[427\]\[1\] _04519_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08804__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09852__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12331_ _05692_ mod.u_cpu.rf_ram.memory\[184\]\[1\] _05704_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15050_ _00904_ net3 mod.u_cpu.rf_ram.memory\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12262_ _05659_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09604__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14001_ _05801_ _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11213_ _04936_ mod.u_cpu.rf_ram.memory\[328\]\[1\] _04942_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput6 net6 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12193_ _05605_ mod.u_cpu.rf_ram.memory\[202\]\[0\] _05612_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14323__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15449__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11144_ _03809_ _03980_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14105__A2 _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12116__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13313__B1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11075_ _04851_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13864__A1 _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12911__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10026_ _04127_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14903_ _00757_ net3 mod.u_cpu.rf_ram.memory\[233\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14473__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15599__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14834_ _00688_ net3 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13616__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14765_ _00619_ net3 mod.u_cpu.rf_ram.memory\[305\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11977_ _05229_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13716_ _05784_ _06723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10928_ _04748_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14696_ _00550_ net3 mod.u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13647_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_arbiter.i_wb_cpu_rdt\[4\] _06334_
+ _06659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09048__A1 _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12755__S _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10859_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _04222_ _03724_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_72_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13578_ _03692_ _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10602__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15317_ _01096_ net3 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12529_ _05837_ mod.u_cpu.rf_ram.memory\[469\]\[1\] _05842_ _05845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08271__A2 mod.u_cpu.rf_ram.memory\[542\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15248_ _00063_ net4 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15179_ _01032_ net3 mod.u_cpu.rf_ram.memory\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13155__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14816__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__C _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ _03922_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

