// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire \mod.timer_irq ;
 wire \mod.u_arbiter.i_wb_cpu_ack ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \mod.u_arbiter.i_wb_cpu_dbus_we ;
 wire \mod.u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \mod.u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[0] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[10] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[11] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[12] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[13] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[14] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[15] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[16] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[17] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[18] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[19] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[1] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[20] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[21] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[22] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[23] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[24] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[25] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[26] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[27] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[28] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[29] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[2] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[30] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[31] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[3] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[4] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[5] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[6] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[7] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[8] ;
 wire \mod.u_arbiter.i_wb_cpu_rdt[9] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[0] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[10] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[11] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[12] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[13] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[14] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[15] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[16] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[17] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[18] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[19] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[1] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[20] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[21] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[22] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[23] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[24] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[25] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[26] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[27] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[28] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[29] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[2] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[30] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[31] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[3] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[4] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[5] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[6] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[7] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[8] ;
 wire \mod.u_arbiter.o_wb_cpu_adr[9] ;
 wire \mod.u_arbiter.o_wb_cpu_cyc ;
 wire \mod.u_arbiter.o_wb_cpu_we ;
 wire \mod.u_cpu.cpu.alu.add_cy_r ;
 wire \mod.u_cpu.cpu.alu.cmp_r ;
 wire \mod.u_cpu.cpu.alu.i_rs1 ;
 wire \mod.u_cpu.cpu.bne_or_bge ;
 wire \mod.u_cpu.cpu.branch_op ;
 wire \mod.u_cpu.cpu.bufreg.c_r ;
 wire \mod.u_cpu.cpu.bufreg.i_sh_signed ;
 wire \mod.u_cpu.cpu.bufreg.lsb[0] ;
 wire \mod.u_cpu.cpu.bufreg.lsb[1] ;
 wire \mod.u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \mod.u_cpu.cpu.csr_d_sel ;
 wire \mod.u_cpu.cpu.csr_imm ;
 wire \mod.u_cpu.cpu.ctrl.i_iscomp ;
 wire \mod.u_cpu.cpu.ctrl.i_jump ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \mod.u_cpu.cpu.decode.co_ebreak ;
 wire \mod.u_cpu.cpu.decode.co_mem_word ;
 wire \mod.u_cpu.cpu.decode.op21 ;
 wire \mod.u_cpu.cpu.decode.op22 ;
 wire \mod.u_cpu.cpu.decode.op26 ;
 wire \mod.u_cpu.cpu.decode.opcode[0] ;
 wire \mod.u_cpu.cpu.decode.opcode[1] ;
 wire \mod.u_cpu.cpu.decode.opcode[2] ;
 wire \mod.u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \mod.u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \mod.u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \mod.u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \mod.u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[0] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[1] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[2] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[3] ;
 wire \mod.u_cpu.cpu.immdec.imm11_7[4] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \mod.u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[0] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[1] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[2] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[3] ;
 wire \mod.u_cpu.cpu.immdec.imm24_20[4] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[0] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[1] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[2] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[3] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[4] ;
 wire \mod.u_cpu.cpu.immdec.imm30_25[5] ;
 wire \mod.u_cpu.cpu.immdec.imm31 ;
 wire \mod.u_cpu.cpu.immdec.imm7 ;
 wire \mod.u_cpu.cpu.mem_bytecnt[0] ;
 wire \mod.u_cpu.cpu.mem_bytecnt[1] ;
 wire \mod.u_cpu.cpu.mem_if.signbit ;
 wire \mod.u_cpu.cpu.o_wdata0 ;
 wire \mod.u_cpu.cpu.o_wdata1 ;
 wire \mod.u_cpu.cpu.o_wen0 ;
 wire \mod.u_cpu.cpu.o_wen1 ;
 wire \mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \mod.u_cpu.cpu.state.ibus_cyc ;
 wire \mod.u_cpu.cpu.state.init_done ;
 wire \mod.u_cpu.cpu.state.o_cnt[2] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[0] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[1] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[2] ;
 wire \mod.u_cpu.cpu.state.o_cnt_r[3] ;
 wire \mod.u_cpu.cpu.state.stage_two_req ;
 wire \mod.u_cpu.raddr[0] ;
 wire \mod.u_cpu.raddr[1] ;
 wire \mod.u_cpu.rf_ram.addr[0] ;
 wire \mod.u_cpu.rf_ram.addr[1] ;
 wire \mod.u_cpu.rf_ram.addr[2] ;
 wire \mod.u_cpu.rf_ram.addr[3] ;
 wire \mod.u_cpu.rf_ram.addr[4] ;
 wire \mod.u_cpu.rf_ram.addr[5] ;
 wire \mod.u_cpu.rf_ram.addr[6] ;
 wire \mod.u_cpu.rf_ram.addr[7] ;
 wire \mod.u_cpu.rf_ram.data[0] ;
 wire \mod.u_cpu.rf_ram.data[1] ;
 wire \mod.u_cpu.rf_ram.data[2] ;
 wire \mod.u_cpu.rf_ram.data[3] ;
 wire \mod.u_cpu.rf_ram.data[4] ;
 wire \mod.u_cpu.rf_ram.data[5] ;
 wire \mod.u_cpu.rf_ram.data[6] ;
 wire \mod.u_cpu.rf_ram.data[7] ;
 wire \mod.u_cpu.rf_ram.i_wdata[0] ;
 wire \mod.u_cpu.rf_ram.i_wdata[1] ;
 wire \mod.u_cpu.rf_ram.i_wdata[2] ;
 wire \mod.u_cpu.rf_ram.i_wdata[3] ;
 wire \mod.u_cpu.rf_ram.i_wdata[4] ;
 wire \mod.u_cpu.rf_ram.i_wdata[5] ;
 wire \mod.u_cpu.rf_ram.i_wdata[6] ;
 wire \mod.u_cpu.rf_ram.i_wdata[7] ;
 wire \mod.u_cpu.rf_ram.rdata[0] ;
 wire \mod.u_cpu.rf_ram.rdata[1] ;
 wire \mod.u_cpu.rf_ram.rdata[2] ;
 wire \mod.u_cpu.rf_ram.rdata[3] ;
 wire \mod.u_cpu.rf_ram.rdata[4] ;
 wire \mod.u_cpu.rf_ram.rdata[5] ;
 wire \mod.u_cpu.rf_ram.rdata[6] ;
 wire \mod.u_cpu.rf_ram.rdata[7] ;
 wire \mod.u_cpu.rf_ram.regzero ;
 wire \mod.u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \mod.u_cpu.rf_ram_if.rcnt[0] ;
 wire \mod.u_cpu.rf_ram_if.rcnt[1] ;
 wire \mod.u_cpu.rf_ram_if.rcnt[2] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[1] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[2] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[3] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[4] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[5] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[6] ;
 wire \mod.u_cpu.rf_ram_if.rdata0[7] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[0] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[1] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[2] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[3] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[4] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[5] ;
 wire \mod.u_cpu.rf_ram_if.rdata1[6] ;
 wire \mod.u_cpu.rf_ram_if.rgnt ;
 wire \mod.u_cpu.rf_ram_if.rreq_r ;
 wire \mod.u_cpu.rf_ram_if.rtrig0 ;
 wire \mod.u_cpu.rf_ram_if.rtrig1 ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \mod.u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \mod.u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \mod.u_cpu.rf_ram_if.wen0_r ;
 wire \mod.u_cpu.rf_ram_if.wen1_r ;
 wire \mod.u_cpu.rf_ram_if.wtrig0 ;
 wire \mod.u_scanchain_local.clk ;
 wire \mod.u_scanchain_local.clk_out ;
 wire \mod.u_scanchain_local.data_out ;
 wire \mod.u_scanchain_local.data_out_i ;
 wire \mod.u_scanchain_local.module_data_in[34] ;
 wire \mod.u_scanchain_local.module_data_in[35] ;
 wire \mod.u_scanchain_local.module_data_in[36] ;
 wire \mod.u_scanchain_local.module_data_in[37] ;
 wire \mod.u_scanchain_local.module_data_in[38] ;
 wire \mod.u_scanchain_local.module_data_in[39] ;
 wire \mod.u_scanchain_local.module_data_in[40] ;
 wire \mod.u_scanchain_local.module_data_in[41] ;
 wire \mod.u_scanchain_local.module_data_in[42] ;
 wire \mod.u_scanchain_local.module_data_in[43] ;
 wire \mod.u_scanchain_local.module_data_in[44] ;
 wire \mod.u_scanchain_local.module_data_in[45] ;
 wire \mod.u_scanchain_local.module_data_in[46] ;
 wire \mod.u_scanchain_local.module_data_in[47] ;
 wire \mod.u_scanchain_local.module_data_in[48] ;
 wire \mod.u_scanchain_local.module_data_in[49] ;
 wire \mod.u_scanchain_local.module_data_in[50] ;
 wire \mod.u_scanchain_local.module_data_in[51] ;
 wire \mod.u_scanchain_local.module_data_in[52] ;
 wire \mod.u_scanchain_local.module_data_in[53] ;
 wire \mod.u_scanchain_local.module_data_in[54] ;
 wire \mod.u_scanchain_local.module_data_in[55] ;
 wire \mod.u_scanchain_local.module_data_in[56] ;
 wire \mod.u_scanchain_local.module_data_in[57] ;
 wire \mod.u_scanchain_local.module_data_in[58] ;
 wire \mod.u_scanchain_local.module_data_in[59] ;
 wire \mod.u_scanchain_local.module_data_in[60] ;
 wire \mod.u_scanchain_local.module_data_in[61] ;
 wire \mod.u_scanchain_local.module_data_in[62] ;
 wire \mod.u_scanchain_local.module_data_in[63] ;
 wire \mod.u_scanchain_local.module_data_in[64] ;
 wire \mod.u_scanchain_local.module_data_in[65] ;
 wire \mod.u_scanchain_local.module_data_in[66] ;
 wire \mod.u_scanchain_local.module_data_in[67] ;
 wire \mod.u_scanchain_local.module_data_in[68] ;
 wire \mod.u_scanchain_local.module_data_in[69] ;
 wire \clknet_0_mod.u_scanchain_local.clk ;
 wire \clknet_3_0__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_1__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_2__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_3__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_4__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_5__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_6__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_3_7__leaf_mod.u_scanchain_local.clk ;
 wire \clknet_opt_1_0_mod.u_scanchain_local.clk ;
 wire \clknet_opt_1_1_mod.u_scanchain_local.clk ;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1331_ (.I(\mod.u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1332_ (.I(\mod.u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1333_ (.A1(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0822_),
    .A3(_0823_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1334_ (.I(_0824_),
    .ZN(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1335_ (.I(_0824_),
    .ZN(\mod.u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1336_ (.I(\mod.u_cpu.cpu.decode.opcode[2] ),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1337_ (.I(_0825_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1338_ (.I(\mod.u_cpu.cpu.branch_op ),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1339_ (.I(_0827_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1340_ (.A1(_0826_),
    .A2(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1341_ (.I(\mod.u_cpu.cpu.decode.co_mem_word ),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1342_ (.A1(_0830_),
    .A2(\mod.u_cpu.cpu.bne_or_bge ),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1343_ (.A1(\mod.u_cpu.cpu.csr_d_sel ),
    .A2(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1344_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_0829_),
    .A3(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1345_ (.I(\mod.u_cpu.cpu.decode.op26 ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1346_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1347_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1348_ (.I(_0830_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1349_ (.I(\mod.u_cpu.cpu.bne_or_bge ),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1350_ (.I(\mod.u_cpu.cpu.csr_d_sel ),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1351_ (.A1(_0837_),
    .A2(_0838_),
    .A3(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1352_ (.A1(_0829_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1353_ (.A1(_0836_),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1354_ (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1355_ (.A1(_0826_),
    .A2(_0828_),
    .A3(\mod.u_cpu.cpu.decode.op21 ),
    .A4(_0840_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1356_ (.A1(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1357_ (.A1(_0843_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1358_ (.A1(_0842_),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1359_ (.A1(_0833_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1360_ (.A1(_0824_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1361_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0824_),
    .B1(_0849_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1362_ (.A1(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .A2(_0848_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1363_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0824_),
    .B1(_0849_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1364_ (.A1(_0850_),
    .A2(_0851_),
    .A3(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1365_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0847_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1366_ (.A1(\mod.u_cpu.cpu.decode.op26 ),
    .A2(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A3(_0829_),
    .A4(_0840_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1367_ (.A1(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .A2(_0833_),
    .A3(_0854_),
    .A4(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1368_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .B(_0856_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1369_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0824_),
    .B1(_0849_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1370_ (.A1(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A3(_0844_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1371_ (.A1(_0835_),
    .A2(_0859_),
    .B(_0847_),
    .C(_0824_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1372_ (.A1(\mod.u_cpu.cpu.csr_imm ),
    .A2(_0824_),
    .B1(_0849_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .C(_0860_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1373_ (.A1(_0857_),
    .A2(_0858_),
    .A3(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1374_ (.A1(_0853_),
    .A2(_0862_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1375_ (.I(\mod.u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1376_ (.I(\mod.u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1377_ (.A1(_0863_),
    .A2(_0864_),
    .ZN(\mod.u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1378_ (.I(\mod.u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1379_ (.A1(\mod.u_cpu.rf_ram_if.wen1_r ),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1380_ (.A1(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0822_),
    .A3(_0823_),
    .A4(\mod.u_cpu.rf_ram_if.wen0_r ),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1381_ (.A1(_0866_),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1382_ (.I(_0868_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1383_ (.A1(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\mod.u_cpu.rf_ram_if.rcnt[1] ),
    .B(\mod.u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1384_ (.A1(_0868_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1385_ (.A1(\mod.u_cpu.raddr[0] ),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1386_ (.I(_0871_),
    .Z(\mod.u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1387_ (.A1(\mod.u_cpu.raddr[0] ),
    .A2(_0870_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1388_ (.A1(\mod.u_cpu.raddr[1] ),
    .A2(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1389_ (.I(_0873_),
    .Z(\mod.u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1390_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1391_ (.A1(_0874_),
    .A2(_0859_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1392_ (.A1(_0835_),
    .A2(_0846_),
    .B(_0865_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1393_ (.A1(_0865_),
    .A2(_0875_),
    .B(_0876_),
    .C(_0868_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1394_ (.A1(_0861_),
    .A2(_0868_),
    .B(_0877_),
    .ZN(\mod.u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1395_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1396_ (.A1(\mod.u_cpu.cpu.decode.op26 ),
    .A2(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A3(_0865_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1397_ (.A1(_0865_),
    .A2(_0878_),
    .B(_0859_),
    .C(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1398_ (.A1(_0868_),
    .A2(_0880_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1399_ (.A1(_0857_),
    .A2(_0868_),
    .B(_0881_),
    .ZN(\mod.u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1400_ (.A1(_0865_),
    .A2(_0846_),
    .A3(_0026_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1401_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[2] ),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1402_ (.A1(_0858_),
    .A2(_0868_),
    .B1(_0882_),
    .B2(_0883_),
    .ZN(\mod.u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1403_ (.I(_0882_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1404_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1405_ (.A1(_0852_),
    .A2(_0868_),
    .B(_0885_),
    .ZN(\mod.u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1406_ (.I(\mod.u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1407_ (.A1(_0850_),
    .A2(_0868_),
    .B1(_0882_),
    .B2(_0886_),
    .ZN(\mod.u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1408_ (.A1(_0851_),
    .A2(_0026_),
    .B(_0884_),
    .ZN(\mod.u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1409_ (.I(\mod.u_cpu.rf_ram.regzero ),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1410_ (.A1(_0866_),
    .A2(_0867_),
    .B(\mod.u_cpu.rf_ram.rdata[0] ),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1411_ (.I(\mod.u_cpu.rf_ram.data[0] ),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1412_ (.A1(_0889_),
    .A2(_0866_),
    .A3(_0867_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1413_ (.A1(_0888_),
    .A2(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1414_ (.I(_0891_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1415_ (.A1(_0887_),
    .A2(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .A3(_0017_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1416_ (.A1(\mod.u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_0824_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1417_ (.A1(_0892_),
    .A2(_0893_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1418_ (.I0(\mod.u_cpu.rf_ram.rdata[1] ),
    .I1(\mod.u_cpu.rf_ram.data[1] ),
    .S(_0026_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1419_ (.I(_0894_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1420_ (.A1(_0887_),
    .A2(_0018_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1421_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[2] ),
    .I1(_0895_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1422_ (.I(_0896_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1423_ (.I0(\mod.u_cpu.rf_ram.rdata[2] ),
    .I1(\mod.u_cpu.rf_ram.data[2] ),
    .S(_0026_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1424_ (.I(_0897_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1425_ (.A1(_0887_),
    .A2(_0019_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1426_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[3] ),
    .I1(_0898_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1427_ (.I(_0899_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1428_ (.I0(\mod.u_cpu.rf_ram.rdata[3] ),
    .I1(\mod.u_cpu.rf_ram.data[3] ),
    .S(_0026_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1429_ (.I(_0900_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1430_ (.A1(_0887_),
    .A2(_0020_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1431_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[4] ),
    .I1(_0901_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1432_ (.I(_0902_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1433_ (.I0(\mod.u_cpu.rf_ram.rdata[4] ),
    .I1(\mod.u_cpu.rf_ram.data[4] ),
    .S(_0026_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1434_ (.I(_0903_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1435_ (.A1(_0887_),
    .A2(_0021_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1436_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[5] ),
    .I1(_0904_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1437_ (.I(_0905_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1438_ (.I0(\mod.u_cpu.rf_ram.rdata[5] ),
    .I1(\mod.u_cpu.rf_ram.data[5] ),
    .S(_0026_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1439_ (.I(_0906_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1440_ (.A1(_0887_),
    .A2(_0022_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1441_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[6] ),
    .I1(_0907_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1442_ (.I(_0908_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1443_ (.I0(\mod.u_cpu.rf_ram.rdata[6] ),
    .I1(\mod.u_cpu.rf_ram.data[6] ),
    .S(_0026_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1444_ (.I(_0909_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1445_ (.A1(_0887_),
    .A2(_0023_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1446_ (.I0(\mod.u_cpu.rf_ram_if.rdata0[7] ),
    .I1(_0910_),
    .S(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1447_ (.I(_0911_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1448_ (.I(\mod.u_cpu.rf_ram_if.rtrig1 ),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1449_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[1] ),
    .I1(_0895_),
    .S(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1450_ (.I(_0913_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1451_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[2] ),
    .I1(_0898_),
    .S(_0912_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1452_ (.I(_0914_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1453_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[3] ),
    .I1(_0901_),
    .S(_0912_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1454_ (.I(_0915_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1455_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[4] ),
    .I1(_0904_),
    .S(_0912_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1456_ (.I(_0916_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1457_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[5] ),
    .I1(_0907_),
    .S(_0912_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1458_ (.I(_0917_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1459_ (.I0(\mod.u_cpu.rf_ram_if.rdata1[6] ),
    .I1(_0910_),
    .S(_0912_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1460_ (.I(_0918_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1461_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_0865_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1462_ (.I(_0919_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1463_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_0865_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1464_ (.I(_0920_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1465_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_0865_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1466_ (.I(_0921_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1467_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_0865_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1468_ (.I(_0922_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1469_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_0865_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1470_ (.I(_0923_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1471_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_0865_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1472_ (.I(_0924_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1473_ (.I0(\mod.u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\mod.u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_0865_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1474_ (.I(_0925_),
    .Z(\mod.u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1475_ (.I(\mod.u_cpu.cpu.decode.opcode[0] ),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1476_ (.A1(_0825_),
    .A2(_0828_),
    .A3(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1477_ (.I(\mod.u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1478_ (.A1(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .A2(_0928_),
    .A3(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1479_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1480_ (.A1(_0825_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1481_ (.A1(_0926_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1482_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1483_ (.A1(_0828_),
    .A2(_0933_),
    .B1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .B2(_0829_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1484_ (.A1(_0926_),
    .A2(_0931_),
    .B(_0932_),
    .C(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1485_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1486_ (.A1(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1487_ (.I(\mod.u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1488_ (.A1(_0825_),
    .A2(_0827_),
    .A3(\mod.u_cpu.cpu.csr_d_sel ),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1489_ (.A1(\mod.u_cpu.cpu.immdec.imm31 ),
    .A2(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1490_ (.A1(_0938_),
    .A2(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1491_ (.A1(_0926_),
    .A2(_0933_),
    .A3(_0931_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1492_ (.A1(_0926_),
    .A2(_0933_),
    .A3(\mod.u_cpu.cpu.immdec.imm11_7[0] ),
    .A4(_0931_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1493_ (.I(_0938_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1494_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_0942_),
    .B(_0943_),
    .C(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1495_ (.A1(_0941_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1496_ (.A1(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .A2(_0928_),
    .B(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1497_ (.A1(_0927_),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1498_ (.A1(_0837_),
    .A2(_0825_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1499_ (.I(\mod.u_cpu.cpu.state.stage_two_req ),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1500_ (.A1(\mod.u_cpu.cpu.csr_d_sel ),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(\mod.u_cpu.cpu.state.init_done ),
    .C(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1501_ (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1502_ (.A1(_0843_),
    .A2(\mod.u_cpu.cpu.state.init_done ),
    .A3(_0952_),
    .A4(_0828_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1503_ (.I(_0926_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1504_ (.A1(_0828_),
    .A2(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1505_ (.A1(_0837_),
    .A2(_0839_),
    .B(_0831_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1506_ (.A1(_0955_),
    .A2(_0956_),
    .B(_0825_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1507_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1508_ (.A1(_0957_),
    .A2(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1509_ (.A1(_0949_),
    .A2(_0951_),
    .B1(_0953_),
    .B2(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1510_ (.A1(_0864_),
    .A2(_0960_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1511_ (.A1(_0946_),
    .A2(_0948_),
    .B1(_0961_),
    .B2(_0927_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1512_ (.A1(_0937_),
    .A2(_0962_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1513_ (.A1(_0930_),
    .A2(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1514_ (.A1(\mod.u_cpu.cpu.alu.add_cy_r ),
    .A2(\mod.u_cpu.cpu.alu.i_rs1 ),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1515_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .A2(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_0831_),
    .C(_0827_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1516_ (.I(_0912_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1517_ (.A1(\mod.u_cpu.rf_ram.regzero ),
    .A2(_0967_),
    .A3(_0888_),
    .A4(_0890_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1518_ (.A1(_0967_),
    .A2(\mod.u_cpu.rf_ram_if.rdata1[0] ),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1519_ (.A1(_0933_),
    .A2(_0941_),
    .A3(_0945_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1520_ (.A1(_0933_),
    .A2(_0968_),
    .A3(_0969_),
    .B(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1521_ (.A1(_0966_),
    .A2(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1522_ (.A1(_0965_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1523_ (.A1(_0840_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1524_ (.I(\mod.u_cpu.cpu.alu.i_rs1 ),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1525_ (.A1(_0975_),
    .A2(_0971_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1526_ (.A1(_0975_),
    .A2(_0971_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1527_ (.A1(_0838_),
    .A2(_0976_),
    .B(_0977_),
    .C(\mod.u_cpu.cpu.csr_d_sel ),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1528_ (.A1(_0837_),
    .A2(_0976_),
    .B(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1529_ (.A1(_0864_),
    .A2(_0960_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1530_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_0929_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1531_ (.A1(_0830_),
    .A2(_0839_),
    .A3(\mod.u_cpu.cpu.alu.cmp_r ),
    .A4(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1532_ (.A1(_0980_),
    .A2(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1533_ (.A1(_0826_),
    .A2(_0955_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1534_ (.A1(_0974_),
    .A2(_0979_),
    .A3(_0983_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1535_ (.A1(_0968_),
    .A2(_0969_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1536_ (.A1(_0842_),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1537_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_0829_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1538_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1539_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1540_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_0832_),
    .A3(_0988_),
    .A4(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1541_ (.A1(_0938_),
    .A2(\mod.u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1542_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .A2(_0929_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1543_ (.A1(_0929_),
    .A2(_0992_),
    .B(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1544_ (.A1(_0991_),
    .A2(_0994_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1545_ (.I(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1546_ (.I(\mod.u_cpu.cpu.decode.op22 ),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1547_ (.A1(\mod.u_cpu.cpu.decode.op26 ),
    .A2(_0841_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1548_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_0997_),
    .A3(_0929_),
    .A4(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1549_ (.A1(_0996_),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1550_ (.I(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1551_ (.A1(_1001_),
    .A2(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1552_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .B(_0929_),
    .C(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1553_ (.I(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1554_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1555_ (.A1(_1004_),
    .A2(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1556_ (.A1(_0828_),
    .A2(_0954_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1557_ (.I(\mod.u_cpu.cpu.mem_if.signbit ),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1558_ (.A1(_0838_),
    .A2(_0928_),
    .B(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1559_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I2(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I3(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(_0863_),
    .S1(_0864_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1560_ (.A1(_0830_),
    .A2(_1009_),
    .B(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1561_ (.A1(_0830_),
    .A2(_1008_),
    .A3(_1009_),
    .B(_1011_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1562_ (.A1(\mod.u_cpu.cpu.csr_d_sel ),
    .A2(_1011_),
    .B(_0825_),
    .C(_0926_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1563_ (.A1(_1006_),
    .A2(_1007_),
    .B1(_0205_),
    .B2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1564_ (.A1(_0987_),
    .A2(_0995_),
    .A3(_1000_),
    .A4(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1565_ (.I(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1566_ (.A1(_0927_),
    .A2(_0964_),
    .B(_0985_),
    .C(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1567_ (.A1(_0930_),
    .A2(_0963_),
    .B(_0828_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1568_ (.A1(_0827_),
    .A2(_0961_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1569_ (.A1(_0859_),
    .A2(_1017_),
    .A3(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1570_ (.A1(_0859_),
    .A2(_1016_),
    .B(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1571_ (.I(_1020_),
    .ZN(\mod.u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1572_ (.A1(_0865_),
    .A2(\mod.u_cpu.rf_ram_if.wdata1_r[7] ),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1573_ (.A1(_0865_),
    .A2(_1020_),
    .B(_1021_),
    .ZN(\mod.u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1574_ (.I0(\mod.u_cpu.rf_ram.rdata[7] ),
    .I1(\mod.u_cpu.rf_ram.data[7] ),
    .S(_0026_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1575_ (.I(_1022_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1576_ (.A1(_0987_),
    .A2(_0995_),
    .A3(_1000_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1577_ (.A1(\mod.u_cpu.cpu.csr_d_sel ),
    .A2(\mod.u_cpu.cpu.csr_imm ),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1578_ (.A1(\mod.u_cpu.cpu.csr_d_sel ),
    .A2(_0975_),
    .B(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1579_ (.A1(_0837_),
    .A2(_1025_),
    .B(\mod.u_cpu.cpu.bne_or_bge ),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1580_ (.A1(_0831_),
    .A2(_1025_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1581_ (.A1(_0830_),
    .A2(\mod.u_cpu.cpu.bne_or_bge ),
    .B(_1027_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1582_ (.A1(_1023_),
    .A2(_1026_),
    .B(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1583_ (.A1(_0846_),
    .A2(_1029_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1584_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0846_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1585_ (.A1(_1030_),
    .A2(_1031_),
    .ZN(\mod.u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1586_ (.A1(\mod.u_cpu.cpu.alu.add_cy_r ),
    .A2(\mod.u_cpu.cpu.alu.i_rs1 ),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1587_ (.A1(_0965_),
    .A2(_0972_),
    .B(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1588_ (.A1(_0958_),
    .A2(_0966_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1589_ (.A1(_0990_),
    .A2(_1033_),
    .B(_1034_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1590_ (.I(io_in[9]),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1591_ (.I(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1592_ (.A1(_1036_),
    .A2(\mod.u_cpu.cpu.state.ibus_cyc ),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1593_ (.I(_1037_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1594_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1595_ (.I(_1039_),
    .Z(\mod.u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1596_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_1038_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1597_ (.I(_1040_),
    .Z(\mod.u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1598_ (.A1(_1036_),
    .A2(\mod.u_cpu.cpu.state.ibus_cyc ),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1599_ (.I(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1600_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1042_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1601_ (.I(\mod.u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1602_ (.I(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1603_ (.I(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1604_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_1046_),
    .B(_1041_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1605_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_1046_),
    .B(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1606_ (.A1(_1043_),
    .A2(_1048_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1607_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_1046_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1608_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A3(_1046_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1609_ (.A1(_1038_),
    .A2(_1050_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_1042_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1611_ (.A1(_1049_),
    .A2(_1051_),
    .B(_1052_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1612_ (.I(_1041_),
    .Z(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1613_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_1050_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1614_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_1042_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1615_ (.A1(_1053_),
    .A2(_1054_),
    .B(_1055_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1616_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A4(_1044_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1617_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1618_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_1042_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1619_ (.A1(_1053_),
    .A2(_1057_),
    .B(_1058_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1620_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_1056_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1621_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A3(_1056_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1622_ (.A1(_1038_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1623_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_1042_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1624_ (.A1(_1059_),
    .A2(_1061_),
    .B(_1062_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1625_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_1060_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1626_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_1042_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1627_ (.A1(_1053_),
    .A2(_1063_),
    .B(_1064_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1628_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1629_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_1056_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1630_ (.A1(_1065_),
    .A2(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(_1065_),
    .A2(_1066_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1632_ (.A1(_1038_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1633_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_1042_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1634_ (.A1(_1067_),
    .A2(_1069_),
    .B(_1070_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1635_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1636_ (.A1(_1071_),
    .A2(_1067_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1637_ (.I(_1041_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1638_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1639_ (.A1(_1053_),
    .A2(_1072_),
    .B(_1074_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1640_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1641_ (.A1(_1075_),
    .A2(_1071_),
    .A3(_1065_),
    .A4(_1066_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1642_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_1067_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1643_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_1073_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1644_ (.A1(_1053_),
    .A2(_1076_),
    .A3(_1077_),
    .B(_1078_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1645_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_1076_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1646_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_1076_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1647_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_1073_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1648_ (.A1(_1053_),
    .A2(_1079_),
    .A3(_1080_),
    .B(_1081_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1649_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_1079_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1650_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_1073_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1651_ (.A1(_1053_),
    .A2(_1082_),
    .B(_1083_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1652_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_1079_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1653_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A4(_1076_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1654_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_1073_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1655_ (.A1(_1042_),
    .A2(_1084_),
    .A3(_1085_),
    .B(_1086_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1656_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_1085_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1657_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_1085_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1658_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .A2(_1073_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1659_ (.A1(_1042_),
    .A2(_1087_),
    .A3(_1088_),
    .B(_1089_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1660_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_1088_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1661_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_1073_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1662_ (.A1(_1053_),
    .A2(_1090_),
    .B(_1091_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1663_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_1088_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1664_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A4(_1085_),
    .Z(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1665_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .A2(_1073_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1666_ (.A1(_1042_),
    .A2(_1092_),
    .A3(_1093_),
    .B(_1094_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1667_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_1093_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1668_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_1093_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1669_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_1073_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1670_ (.A1(_1042_),
    .A2(_1095_),
    .A3(_1096_),
    .B(_1097_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1671_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_1096_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1672_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .A2(_1073_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1673_ (.A1(_1053_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1674_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A4(_1093_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1675_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_1096_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1676_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_1041_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1677_ (.A1(_1042_),
    .A2(_1100_),
    .A3(_1101_),
    .B(_1102_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1678_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_1100_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1679_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_1100_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1680_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_1041_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1681_ (.A1(_1042_),
    .A2(_1103_),
    .A3(_1104_),
    .B(_1105_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1682_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_1104_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1683_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_1073_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1684_ (.A1(_1053_),
    .A2(_1106_),
    .B(_1107_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1685_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A4(_1100_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1686_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_1104_),
    .B(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1687_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_1041_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1688_ (.A1(_1042_),
    .A2(_1108_),
    .A3(_1109_),
    .B(_1110_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1689_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_1108_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1690_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_1108_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1691_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_1041_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1692_ (.A1(_1042_),
    .A2(_1111_),
    .A3(_1112_),
    .B(_1113_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1693_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_1111_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1694_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_1073_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1695_ (.A1(_1053_),
    .A2(_1114_),
    .B(_1115_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1696_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_1111_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1697_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_1116_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_1073_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1699_ (.A1(_1053_),
    .A2(_1117_),
    .B(_1118_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1700_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1701_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A4(_1108_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1702_ (.A1(_1119_),
    .A2(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1703_ (.A1(_1119_),
    .A2(_1120_),
    .Z(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1704_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_1041_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1705_ (.A1(_1042_),
    .A2(_1121_),
    .A3(_1122_),
    .B(_1123_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1706_ (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1707_ (.A1(_1124_),
    .A2(_1121_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1708_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_1073_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1709_ (.A1(_1053_),
    .A2(_1125_),
    .B(_1126_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1710_ (.A1(_1124_),
    .A2(_1119_),
    .A3(_1120_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1711_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1712_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_1073_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1713_ (.A1(_1053_),
    .A2(_1128_),
    .B(_1129_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1714_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_1127_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1715_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1716_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_1073_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1717_ (.A1(_1053_),
    .A2(_1131_),
    .B(_1132_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1718_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(_1127_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1719_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1720_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_1038_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1721_ (.A1(_1038_),
    .A2(_1134_),
    .B(_1135_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1722_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A3(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A4(_1127_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1723_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1724_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A2(_1038_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1725_ (.A1(_1038_),
    .A2(_1137_),
    .B(_1138_),
    .ZN(\mod.u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1726_ (.I(_0863_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1727_ (.A1(\mod.u_cpu.cpu.bne_or_bge ),
    .A2(_0864_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1728_ (.A1(_1139_),
    .A2(_1140_),
    .B(_0837_),
    .ZN(\mod.u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1729_ (.A1(_1139_),
    .A2(_0864_),
    .B(_0837_),
    .ZN(\mod.u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1730_ (.A1(_0863_),
    .A2(_1140_),
    .B(_0837_),
    .ZN(\mod.u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1731_ (.A1(_0874_),
    .A2(_0878_),
    .A3(_0883_),
    .A4(_0886_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1732_ (.A1(\mod.u_cpu.cpu.state.init_done ),
    .A2(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(_0957_),
    .A2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1734_ (.A1(_0825_),
    .A2(_0827_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1735_ (.A1(_0954_),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1736_ (.A1(_0825_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1737_ (.A1(_0926_),
    .A2(_1144_),
    .B(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1738_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_1141_),
    .B(_1143_),
    .C(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1739_ (.A1(_0859_),
    .A2(_1148_),
    .B(_0990_),
    .ZN(\mod.u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1740_ (.A1(_0847_),
    .A2(_0990_),
    .ZN(\mod.u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1741_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1742_ (.A1(_1004_),
    .A2(_1005_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1743_ (.A1(_0958_),
    .A2(_1143_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1744_ (.A1(_1149_),
    .A2(_1150_),
    .B(_1151_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1745_ (.I(_0936_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1746_ (.A1(_0937_),
    .A2(_0962_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1747_ (.A1(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_1152_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1748_ (.A1(_1151_),
    .A2(_1154_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1749_ (.A1(_0827_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(_0827_),
    .A2(_0954_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1751_ (.A1(\mod.u_cpu.cpu.alu.i_rs1 ),
    .A2(\mod.u_cpu.cpu.bufreg.c_r ),
    .A3(_1155_),
    .A4(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1752_ (.A1(\mod.u_cpu.cpu.alu.i_rs1 ),
    .A2(_1155_),
    .A3(_1156_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1753_ (.A1(\mod.u_cpu.cpu.bufreg.c_r ),
    .A2(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1754_ (.A1(_0954_),
    .A2(\mod.u_cpu.cpu.decode.opcode[1] ),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1755_ (.A1(_0827_),
    .A2(_0981_),
    .A3(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1756_ (.A1(_0826_),
    .A2(_0946_),
    .A3(_1159_),
    .A4(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1757_ (.I(_0960_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1758_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1759_ (.I(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1760_ (.A1(_1157_),
    .A2(_1162_),
    .B(_1165_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1761_ (.A1(_0933_),
    .A2(_1038_),
    .ZN(\mod.u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1762_ (.A1(_0830_),
    .A2(_0863_),
    .B1(_0864_),
    .B2(_0831_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1763_ (.A1(\mod.u_cpu.cpu.state.init_done ),
    .A2(_0990_),
    .A3(_1144_),
    .A4(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1764_ (.A1(_1053_),
    .A2(_1167_),
    .ZN(\mod.u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1765_ (.A1(_0957_),
    .A2(_1142_),
    .B(_0949_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1766_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A3(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1767_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_1169_),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1768_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1769_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1770_ (.A1(_0938_),
    .A2(_0837_),
    .A3(_0825_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1771_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_1173_),
    .B(_1168_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1772_ (.A1(_1168_),
    .A2(_1172_),
    .B(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1773_ (.A1(_0830_),
    .A2(_0839_),
    .A3(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1774_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_1041_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1775_ (.A1(_0827_),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1776_ (.A1(_0826_),
    .A2(_1176_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1777_ (.A1(_0843_),
    .A2(\mod.u_cpu.cpu.state.init_done ),
    .A3(_0990_),
    .A4(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1778_ (.I(_1044_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1779_ (.I(_1181_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1780_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_1038_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1781_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0215_),
    .B(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1782_ (.I(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1783_ (.A1(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\mod.u_cpu.cpu.state.stage_two_req ),
    .B(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1784_ (.A1(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0823_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1785_ (.I(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1786_ (.A1(_0221_),
    .A2(\mod.u_cpu.rf_ram_if.rcnt[1] ),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1787_ (.A1(_0220_),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1788_ (.A1(_0219_),
    .A2(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1789_ (.A1(_1180_),
    .A2(_0224_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1790_ (.A1(_1035_),
    .A2(_0219_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(_1180_),
    .A2(_0219_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1792_ (.A1(\mod.u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_0225_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1793_ (.A1(_0221_),
    .A2(_0822_),
    .A3(_0823_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1794_ (.A1(_0869_),
    .A2(_0225_),
    .A3(_0226_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1795_ (.A1(\mod.u_cpu.raddr[0] ),
    .A2(_0226_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1796_ (.A1(\mod.u_cpu.raddr[0] ),
    .A2(_0226_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1797_ (.A1(_1180_),
    .A2(_0219_),
    .A3(_0227_),
    .A4(_0228_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1798_ (.I(_0229_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1799_ (.A1(\mod.u_cpu.raddr[1] ),
    .A2(_0227_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1800_ (.A1(_0225_),
    .A2(_0230_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1801_ (.A1(_1036_),
    .A2(\mod.u_cpu.rf_ram_if.rreq_r ),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1802_ (.I(_0231_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1803_ (.I(_0024_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1804_ (.A1(\mod.u_cpu.rf_ram.regzero ),
    .A2(_0824_),
    .A3(_0232_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1805_ (.A1(\mod.u_cpu.rf_ram.regzero ),
    .A2(_0967_),
    .A3(_0232_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1806_ (.A1(_0938_),
    .A2(_0218_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1807_ (.A1(\mod.u_cpu.cpu.state.ibus_cyc ),
    .A2(_0233_),
    .B(_1035_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1808_ (.A1(_1151_),
    .A2(_0233_),
    .B(_0234_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1809_ (.I(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1810_ (.A1(_0938_),
    .A2(_1143_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1811_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\mod.timer_irq ),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1812_ (.A1(_0236_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1813_ (.A1(_0944_),
    .A2(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ),
    .B1(_0235_),
    .B2(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1814_ (.A1(_1035_),
    .A2(_0239_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1815_ (.A1(_1045_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1816_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1817_ (.A1(_1045_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[0] ),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1819_ (.A1(_0242_),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1820_ (.A1(_0241_),
    .A2(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1821_ (.A1(_0242_),
    .A2(_0243_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1822_ (.I(_0246_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1823_ (.A1(_1044_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1824_ (.A1(_1181_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_0248_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1825_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_1044_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1826_ (.I(_0250_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1827_ (.A1(_0249_),
    .A2(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1828_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_1045_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1829_ (.A1(_0247_),
    .A2(_0252_),
    .B(_0253_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1830_ (.A1(_0245_),
    .A2(_0254_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1831_ (.A1(_0218_),
    .A2(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1832_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0215_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1833_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(_1038_),
    .A3(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1834_ (.I(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1835_ (.A1(\mod.u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1836_ (.A1(_0256_),
    .A2(_0260_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1837_ (.A1(_0938_),
    .A2(_0846_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1838_ (.A1(_0833_),
    .A2(_0999_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1839_ (.A1(_0996_),
    .A2(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1840_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_0833_),
    .B(_0262_),
    .C(_0859_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1841_ (.A1(_0833_),
    .A2(_1029_),
    .B(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1842_ (.A1(_0261_),
    .A2(_0263_),
    .B(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1843_ (.I(_0266_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1844_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1845_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_0928_),
    .A3(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .A4(_0997_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1846_ (.A1(_0998_),
    .A2(_0267_),
    .A3(_0268_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1847_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(_0269_),
    .B(_1036_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1848_ (.A1(_1029_),
    .A2(_0269_),
    .B(_0270_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1849_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_0261_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1850_ (.A1(_0996_),
    .A2(_0261_),
    .B(_0271_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1851_ (.A1(_0952_),
    .A2(_1030_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1852_ (.A1(_0944_),
    .A2(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A3(_0832_),
    .A4(_0988_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1853_ (.A1(_0846_),
    .A2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1854_ (.I0(_0272_),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mcause31 ),
    .S(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1855_ (.I(_0275_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1856_ (.I(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1857_ (.A1(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_0276_),
    .B(_0845_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1858_ (.A1(_0938_),
    .A2(_0846_),
    .B1(_0929_),
    .B2(_0991_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1859_ (.I0(_0277_),
    .I1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .S(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1860_ (.I(_0279_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1861_ (.I(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1862_ (.A1(_0827_),
    .A2(_0933_),
    .B1(_0280_),
    .B2(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .C(_0845_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1863_ (.A1(_0278_),
    .A2(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1864_ (.A1(_0276_),
    .A2(_0278_),
    .B(_0282_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1865_ (.A1(_0952_),
    .A2(_0827_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1866_ (.A1(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .A2(_0859_),
    .B(_0278_),
    .C(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1867_ (.A1(_0280_),
    .A2(_0278_),
    .B(_0284_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1868_ (.I(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1869_ (.I(\mod.u_cpu.cpu.decode.co_ebreak ),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1870_ (.A1(_0286_),
    .A2(_0844_),
    .B(_0278_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1871_ (.A1(_0285_),
    .A2(_0278_),
    .B1(_0287_),
    .B2(_1030_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1872_ (.I(_0216_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1873_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1874_ (.I(_0289_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1875_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_0288_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1876_ (.I(_0290_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1877_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_0288_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1878_ (.I(_0291_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1879_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_0288_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1880_ (.I(_0292_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1881_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_0288_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1882_ (.I(_0293_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1883_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_0288_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1884_ (.I(_0294_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1885_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_0288_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1886_ (.I(_0295_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1887_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_0288_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1888_ (.I(_0296_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1889_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_0288_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1890_ (.I(_0297_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1891_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_0288_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1892_ (.I(_0298_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1893_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_0288_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1894_ (.I(_0299_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1895_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_0288_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1896_ (.I(_0300_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1897_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_0288_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1898_ (.I(_0301_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1899_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_0288_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1900_ (.I(_0302_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1901_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_0288_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1902_ (.I(_0303_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1903_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_0288_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1904_ (.I(_0304_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1905_ (.A1(\mod.u_arbiter.i_wb_cpu_ack ),
    .A2(\mod.u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1906_ (.A1(_1046_),
    .A2(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1907_ (.A1(_1035_),
    .A2(_0306_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1908_ (.A1(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_0259_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1909_ (.A1(_0258_),
    .A2(_0255_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1910_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_1046_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1911_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_1044_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1912_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_1044_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1913_ (.A1(_1044_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1914_ (.A1(_1181_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1915_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_1044_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1916_ (.I(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1917_ (.A1(_0313_),
    .A2(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1918_ (.A1(_0310_),
    .A2(_0311_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1919_ (.A1(_0316_),
    .A2(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1920_ (.A1(_1045_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1921_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1922_ (.A1(_0319_),
    .A2(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1923_ (.A1(_0310_),
    .A2(_0321_),
    .B(_0311_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1924_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_1045_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1925_ (.A1(_1044_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1926_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1927_ (.A1(_0323_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1928_ (.A1(_1045_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1929_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1930_ (.A1(_0327_),
    .A2(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1931_ (.A1(_0326_),
    .A2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1932_ (.A1(_0310_),
    .A2(_0311_),
    .B1(_0318_),
    .B2(_0322_),
    .C(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1933_ (.A1(_0319_),
    .A2(_0320_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1934_ (.A1(_0327_),
    .A2(_0328_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1935_ (.A1(_0251_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1936_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_1044_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1937_ (.A1(_0249_),
    .A2(_0325_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1938_ (.A1(_0329_),
    .A2(_0336_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1939_ (.A1(_0251_),
    .A2(_0332_),
    .B1(_0334_),
    .B2(_0335_),
    .C(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1940_ (.A1(_0323_),
    .A2(_0251_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(_0333_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1942_ (.A1(_0253_),
    .A2(_0247_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1943_ (.A1(_0332_),
    .A2(_0340_),
    .B(_0341_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1944_ (.A1(_0331_),
    .A2(_0338_),
    .B(_0342_),
    .C(_0258_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1945_ (.A1(_0308_),
    .A2(_0309_),
    .B(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1946_ (.A1(_0307_),
    .A2(_0344_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1947_ (.A1(_0990_),
    .A2(_1147_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1948_ (.A1(_0218_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1949_ (.A1(_1044_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1950_ (.A1(_1181_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1951_ (.A1(_0347_),
    .A2(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1952_ (.A1(_0347_),
    .A2(_0348_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1953_ (.A1(_0251_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1954_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_1045_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1955_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_1045_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1956_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_1045_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1957_ (.A1(_0316_),
    .A2(_0352_),
    .A3(_0353_),
    .A4(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1958_ (.I(_0335_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1959_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_1044_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1960_ (.A1(_0310_),
    .A2(_0311_),
    .A3(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1961_ (.A1(_0356_),
    .A2(_0350_),
    .A3(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1962_ (.A1(_0349_),
    .A2(_0355_),
    .B(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1963_ (.A1(_0321_),
    .A2(_0355_),
    .B(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1964_ (.A1(_0249_),
    .A2(_0351_),
    .B1(_0361_),
    .B2(_0252_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1965_ (.A1(_0339_),
    .A2(_0350_),
    .B(_0362_),
    .C(_0244_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1966_ (.A1(_0253_),
    .A2(_0244_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1967_ (.A1(_0249_),
    .A2(_0325_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1968_ (.A1(_0332_),
    .A2(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1969_ (.A1(_0330_),
    .A2(_0349_),
    .B1(_0351_),
    .B2(_0249_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1970_ (.A1(_0241_),
    .A2(_0244_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1971_ (.A1(_0337_),
    .A2(_0350_),
    .B1(_0366_),
    .B2(_0367_),
    .C(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1972_ (.A1(_0363_),
    .A2(_0364_),
    .A3(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1973_ (.A1(_0241_),
    .A2(_0247_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1974_ (.A1(_0252_),
    .A2(_0349_),
    .B1(_0354_),
    .B2(_0249_),
    .C(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1975_ (.A1(_0256_),
    .A2(_0370_),
    .A3(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1976_ (.A1(_0308_),
    .A2(_0349_),
    .B(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1977_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0259_),
    .B(_0346_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1978_ (.A1(_0874_),
    .A2(_0346_),
    .B1(_0374_),
    .B2(_0375_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1979_ (.I(_0258_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1980_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_0376_),
    .B1(_0308_),
    .B2(_0335_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1981_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_0346_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1982_ (.A1(_0325_),
    .A2(_0329_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1983_ (.A1(_0323_),
    .A2(_0251_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1984_ (.A1(_0379_),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1985_ (.A1(_0353_),
    .A2(_0365_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1986_ (.A1(_0356_),
    .A2(_0381_),
    .B(_0382_),
    .C(_0244_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1987_ (.A1(_0323_),
    .A2(_0355_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1988_ (.A1(_0245_),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1989_ (.A1(_0365_),
    .A2(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1990_ (.A1(_0254_),
    .A2(_0383_),
    .B1(_0386_),
    .B2(_0335_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1991_ (.A1(_0252_),
    .A2(_0335_),
    .B1(_0353_),
    .B2(_0249_),
    .C(_0371_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1992_ (.A1(_0376_),
    .A2(_0387_),
    .A3(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1993_ (.A1(_0346_),
    .A2(_0377_),
    .B(_0378_),
    .C(_0389_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1994_ (.I(_0218_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1995_ (.A1(_0249_),
    .A2(_0352_),
    .B1(_0357_),
    .B2(_0252_),
    .C1(_0365_),
    .C2(_0314_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1996_ (.A1(_0334_),
    .A2(_0365_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1997_ (.A1(_0352_),
    .A2(_0365_),
    .B1(_0392_),
    .B2(_0357_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1998_ (.A1(_0371_),
    .A2(_0391_),
    .B1(_0393_),
    .B2(_0368_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1999_ (.A1(_0245_),
    .A2(_0252_),
    .A3(_0355_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2000_ (.A1(_0254_),
    .A2(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2001_ (.A1(_0255_),
    .A2(_0394_),
    .B1(_0396_),
    .B2(_0357_),
    .C(_0376_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2002_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0345_),
    .B(_0218_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2003_ (.A1(_0883_),
    .A2(_0390_),
    .A3(_0345_),
    .B1(_0397_),
    .B2(_0398_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2004_ (.A1(_1045_),
    .A2(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2005_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2006_ (.A1(_0379_),
    .A2(_0341_),
    .B(_0396_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2007_ (.A1(\mod.u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_0345_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2008_ (.A1(_0886_),
    .A2(_0345_),
    .B(_0402_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2009_ (.A1(_0252_),
    .A2(_0333_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2010_ (.A1(_0249_),
    .A2(_0310_),
    .B(_0364_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2011_ (.A1(_0404_),
    .A2(_0368_),
    .B(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2012_ (.A1(_0245_),
    .A2(_0254_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2013_ (.I(_0407_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2014_ (.A1(_0258_),
    .A2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2015_ (.A1(_0376_),
    .A2(_0403_),
    .B1(_0406_),
    .B2(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2016_ (.A1(_0259_),
    .A2(_0400_),
    .A3(_0401_),
    .B(_0410_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2017_ (.A1(_0244_),
    .A2(_0249_),
    .A3(_0379_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2018_ (.A1(_0255_),
    .A2(_0380_),
    .A3(_0385_),
    .A4(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2019_ (.A1(_0390_),
    .A2(_0311_),
    .A3(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2020_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0259_),
    .B(_0346_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2021_ (.A1(_0886_),
    .A2(_0346_),
    .B1(_0413_),
    .B2(_0414_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2022_ (.A1(_0958_),
    .A2(_1143_),
    .B(_1035_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2023_ (.I(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2024_ (.A1(_1035_),
    .A2(_1151_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2025_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2026_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2027_ (.I(_0419_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2028_ (.A1(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2029_ (.I(_0420_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2030_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2031_ (.I(_0421_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2032_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2033_ (.I(_0422_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2034_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2035_ (.I(_0423_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2036_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2037_ (.I(_0424_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2038_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2039_ (.I(_0425_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2040_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2041_ (.I(_0426_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2042_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2043_ (.I(_0427_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2044_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2045_ (.I(_0428_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2046_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2047_ (.I(_0429_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2048_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2049_ (.I(_0430_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2050_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2051_ (.I(_0431_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2052_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2053_ (.I(_0432_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2054_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_0416_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2055_ (.I(_0433_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2056_ (.I(_0415_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2057_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_0434_),
    .B1(_0418_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2058_ (.I(_0435_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2059_ (.I(_0417_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2060_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2061_ (.I(_0437_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2062_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2063_ (.I(_0438_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2064_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2065_ (.I(_0439_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2066_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2067_ (.I(_0440_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2068_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2069_ (.I(_0441_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2070_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2071_ (.I(_0442_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2072_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2073_ (.I(_0443_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2074_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2075_ (.I(_0444_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2076_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2077_ (.I(_0445_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2078_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2079_ (.I(_0446_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2080_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2081_ (.I(_0447_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2082_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2083_ (.I(_0448_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2084_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2085_ (.I(_0449_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2086_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2087_ (.I(_0450_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2088_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_0434_),
    .B1(_0436_),
    .B2(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2089_ (.I(_0451_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2090_ (.A1(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_0416_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2091_ (.A1(\mod.u_cpu.cpu.ctrl.i_jump ),
    .A2(_1006_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2092_ (.A1(_0859_),
    .A2(_0833_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2093_ (.A1(\mod.u_cpu.cpu.ctrl.i_jump ),
    .A2(_0964_),
    .B(_0453_),
    .C(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2094_ (.A1(_0454_),
    .A2(_0930_),
    .A3(_0986_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2095_ (.A1(_0455_),
    .A2(_0456_),
    .B(_0436_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_0452_),
    .A2(_0457_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2097_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .B(_0929_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2098_ (.A1(_0960_),
    .A2(_1143_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2099_ (.A1(_1143_),
    .A2(_0458_),
    .B(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2100_ (.A1(_0864_),
    .A2(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2101_ (.A1(_1139_),
    .A2(_0460_),
    .B(_0461_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2102_ (.A1(_0826_),
    .A2(_0946_),
    .A3(_1161_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2103_ (.A1(_1159_),
    .A2(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2104_ (.A1(_1143_),
    .A2(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2105_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_1143_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2106_ (.A1(_0464_),
    .A2(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2107_ (.A1(_0460_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2108_ (.A1(_1139_),
    .A2(_0460_),
    .B(_0467_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2109_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_1164_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2110_ (.I(_0468_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2111_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_1164_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2112_ (.I(_0469_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2113_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_1164_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2114_ (.I(_0470_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2115_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_1164_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2116_ (.I(_0471_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2117_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_1164_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2118_ (.I(_0472_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2119_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_1164_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2120_ (.I(_0473_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2121_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_1164_),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2122_ (.I(_0474_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2123_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_1164_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2124_ (.I(_0475_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2125_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_1164_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2126_ (.I(_0476_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2127_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_1164_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2128_ (.I(_0477_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2129_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_1164_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2130_ (.I(_0478_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2131_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_1164_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2132_ (.I(_0479_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2133_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_1164_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2134_ (.I(_0480_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2135_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_1164_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2136_ (.I(_0481_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2137_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_1164_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2138_ (.I(_0482_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2139_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_1163_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2140_ (.I(_0483_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2141_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_1163_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2142_ (.I(_0484_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2143_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_1163_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2144_ (.I(_0485_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2145_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_1163_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2146_ (.I(_0486_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2147_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_1163_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2148_ (.I(_0487_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2149_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_1163_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2150_ (.I(_0488_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2151_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_1163_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2152_ (.I(_0489_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2153_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_1163_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2154_ (.I(_0490_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2155_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_1163_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2156_ (.I(_0491_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2157_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_1163_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2158_ (.I(_0492_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2159_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_1163_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2160_ (.I(_0493_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2161_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_1163_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2162_ (.I(_0494_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2163_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_1163_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2164_ (.I(_0495_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2165_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .S(_1163_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2166_ (.I(_0496_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2167_ (.A1(\mod.u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A3(_1143_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_0464_),
    .A2(_0497_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2169_ (.I0(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_0498_),
    .S(_1163_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2170_ (.I(_0499_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2171_ (.A1(_0837_),
    .A2(_0839_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2172_ (.I0(_0946_),
    .I1(_0986_),
    .S(\mod.u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2173_ (.A1(\mod.u_cpu.cpu.bne_or_bge ),
    .A2(\mod.u_cpu.cpu.csr_d_sel ),
    .B(_0830_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2174_ (.A1(_0501_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2175_ (.A1(\mod.u_cpu.cpu.alu.i_rs1 ),
    .A2(_0502_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2176_ (.A1(_1033_),
    .A2(_0503_),
    .A3(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2177_ (.I(\mod.u_cpu.cpu.alu.cmp_r ),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2178_ (.A1(_0506_),
    .A2(_0930_),
    .B(_0500_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2179_ (.A1(_0500_),
    .A2(_0505_),
    .B1(_0507_),
    .B2(_0973_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(\mod.u_cpu.cpu.alu.cmp_r ),
    .A2(_0990_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2181_ (.A1(_0990_),
    .A2(_0508_),
    .B(_0509_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2182_ (.A1(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A2(_0236_),
    .B(_0238_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2183_ (.I(_0510_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2184_ (.I(\mod.u_cpu.cpu.immdec.imm31 ),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_0332_),
    .A2(_0334_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2186_ (.A1(_0340_),
    .A2(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2187_ (.A1(_0251_),
    .A2(_0332_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2188_ (.A1(_0400_),
    .A2(_0311_),
    .A3(_0332_),
    .A4(_0330_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2189_ (.A1(_0514_),
    .A2(_0515_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2190_ (.A1(_0321_),
    .A2(_0337_),
    .B(_0368_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2191_ (.A1(_0513_),
    .A2(_0516_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2192_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_1046_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2193_ (.A1(_0408_),
    .A2(_0519_),
    .B(_0376_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2194_ (.A1(_0511_),
    .A2(_0259_),
    .B1(_0518_),
    .B2(_0520_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2195_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2196_ (.A1(_0826_),
    .A2(_0926_),
    .B(_0931_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2197_ (.A1(_0939_),
    .A2(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2198_ (.A1(_0958_),
    .A2(_0523_),
    .B(_0218_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2199_ (.I(_0524_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2200_ (.A1(_0333_),
    .A2(_0354_),
    .A3(_0380_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2201_ (.A1(_0249_),
    .A2(_0251_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2202_ (.A1(_0333_),
    .A2(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2203_ (.A1(_0335_),
    .A2(_0350_),
    .A3(_0358_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(_0528_),
    .A2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2205_ (.A1(_0379_),
    .A2(_0530_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2206_ (.A1(_0332_),
    .A2(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2207_ (.A1(_0244_),
    .A2(_0526_),
    .A3(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2208_ (.A1(_0321_),
    .A2(_0359_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2209_ (.A1(_0252_),
    .A2(_0355_),
    .A3(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2210_ (.A1(_0354_),
    .A2(_0527_),
    .B(_0241_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2211_ (.A1(_0354_),
    .A2(_0365_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2212_ (.A1(_0535_),
    .A2(_0536_),
    .B1(_0537_),
    .B2(_0364_),
    .C(_0256_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2213_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_1046_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2214_ (.A1(_0533_),
    .A2(_0538_),
    .B1(_0539_),
    .B2(_0308_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2215_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_0259_),
    .B(_0525_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2216_ (.A1(_0521_),
    .A2(_0525_),
    .B1(_0540_),
    .B2(_0541_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2217_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2218_ (.A1(_0528_),
    .A2(_0529_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2219_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_1045_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2220_ (.A1(_0544_),
    .A2(_0314_),
    .B(_0317_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2221_ (.A1(_0404_),
    .A2(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2222_ (.A1(_0329_),
    .A2(_0365_),
    .B1(_0543_),
    .B2(_0354_),
    .C(_0546_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2223_ (.A1(_0379_),
    .A2(_0368_),
    .B(_0255_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2224_ (.A1(_0245_),
    .A2(_0339_),
    .B1(_0548_),
    .B2(_0332_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2225_ (.A1(_0368_),
    .A2(_0547_),
    .B(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2226_ (.A1(_0390_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2227_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_0259_),
    .B(_0525_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2228_ (.A1(_0542_),
    .A2(_0525_),
    .B1(_0551_),
    .B2(_0552_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2229_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2230_ (.A1(_0314_),
    .A2(_0400_),
    .B(_0311_),
    .C(_0330_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2231_ (.A1(_0353_),
    .A2(_0543_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2232_ (.A1(_0512_),
    .A2(_0554_),
    .A3(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2233_ (.A1(_0247_),
    .A2(_0251_),
    .B1(_0341_),
    .B2(_0556_),
    .C(_0408_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2234_ (.A1(_0408_),
    .A2(_0333_),
    .B(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2235_ (.A1(_0390_),
    .A2(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2236_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_0376_),
    .B(_0525_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2237_ (.A1(_0553_),
    .A2(_0525_),
    .B1(_0559_),
    .B2(_0560_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2238_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2239_ (.I(_0352_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2240_ (.A1(_0318_),
    .A2(_0404_),
    .B1(_0562_),
    .B2(_0530_),
    .C(_0512_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2241_ (.A1(_0251_),
    .A2(_0408_),
    .B1(_0341_),
    .B2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2242_ (.A1(_0376_),
    .A2(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2243_ (.A1(\mod.u_cpu.cpu.csr_imm ),
    .A2(_0376_),
    .B(_0525_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2244_ (.A1(_0561_),
    .A2(_0525_),
    .B1(_0565_),
    .B2(_0566_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2245_ (.I(\mod.u_cpu.cpu.csr_imm ),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2246_ (.A1(_0339_),
    .A2(_0371_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2247_ (.A1(_0249_),
    .A2(_0332_),
    .A3(_0355_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2248_ (.A1(_0245_),
    .A2(_0325_),
    .A3(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2249_ (.A1(_0330_),
    .A2(_0365_),
    .B(_0349_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2250_ (.A1(_0544_),
    .A2(_0543_),
    .B(_0513_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2251_ (.A1(_0337_),
    .A2(_0350_),
    .B1(_0571_),
    .B2(_0572_),
    .C(_0368_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2252_ (.A1(_0351_),
    .A2(_0568_),
    .B1(_0570_),
    .B2(_0349_),
    .C(_0573_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2253_ (.A1(_0256_),
    .A2(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2254_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0376_),
    .B1(_0323_),
    .B2(_0308_),
    .C(_0524_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2255_ (.A1(_0567_),
    .A2(_0525_),
    .B1(_0575_),
    .B2(_0576_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2256_ (.I(\mod.u_arbiter.i_wb_cpu_rdt[0] ),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2257_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2258_ (.A1(_0215_),
    .A2(_0577_),
    .B(_0578_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2259_ (.A1(_0315_),
    .A2(_0529_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2260_ (.A1(_0528_),
    .A2(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2261_ (.A1(_0323_),
    .A2(_0379_),
    .A3(_0335_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2262_ (.A1(_0340_),
    .A2(_0512_),
    .A3(_0581_),
    .A4(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2263_ (.A1(_0335_),
    .A2(_0340_),
    .B(_0341_),
    .C(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2264_ (.A1(_0335_),
    .A2(_0569_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2265_ (.A1(_0253_),
    .A2(_0325_),
    .A3(_0585_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2266_ (.A1(_0247_),
    .A2(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2267_ (.A1(_0251_),
    .A2(_0335_),
    .B1(_0579_),
    .B2(_0252_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2268_ (.A1(_0584_),
    .A2(_0587_),
    .B1(_0588_),
    .B2(_0568_),
    .C(_0408_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2269_ (.A1(_0408_),
    .A2(_0579_),
    .B(_0589_),
    .C(_0258_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2270_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_0218_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2271_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_0525_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2272_ (.A1(_0525_),
    .A2(_0590_),
    .A3(_0591_),
    .B(_0592_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2273_ (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2274_ (.A1(_0379_),
    .A2(_0357_),
    .A3(_0527_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2275_ (.A1(_0532_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2276_ (.A1(_0357_),
    .A2(_0570_),
    .B1(_0595_),
    .B2(_0241_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2277_ (.A1(_0251_),
    .A2(_0357_),
    .A3(_0364_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2278_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2279_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_0408_),
    .C(_0598_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2280_ (.A1(_0364_),
    .A2(_0596_),
    .B(_0597_),
    .C(_0599_),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2281_ (.A1(_0390_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2282_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0376_),
    .B(_0525_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2283_ (.A1(_0593_),
    .A2(_0525_),
    .B1(_0601_),
    .B2(_0602_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2284_ (.A1(_0379_),
    .A2(_0527_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2285_ (.A1(_0400_),
    .A2(_0337_),
    .B1(_0532_),
    .B2(_0603_),
    .C(_0368_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2286_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2287_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .B(_0407_),
    .C(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2288_ (.A1(_0325_),
    .A2(_0371_),
    .B(_0606_),
    .C(_0218_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2289_ (.A1(_0310_),
    .A2(_0570_),
    .B(_0604_),
    .C(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2290_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_0218_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_0525_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2292_ (.A1(_0525_),
    .A2(_0608_),
    .A3(_0609_),
    .B(_0610_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2293_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .S(_1046_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2294_ (.A1(_0311_),
    .A2(_0337_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2295_ (.A1(_0532_),
    .A2(_0612_),
    .B(_0368_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2296_ (.A1(_0311_),
    .A2(_0570_),
    .B1(_0611_),
    .B2(_0408_),
    .C(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(_0827_),
    .A2(_0940_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2298_ (.A1(_0828_),
    .A2(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .B(_0218_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2299_ (.A1(_0218_),
    .A2(_0614_),
    .B1(_0615_),
    .B2(_0616_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2300_ (.I0(_0617_),
    .I1(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ),
    .S(_0525_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2301_ (.I(_0618_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2302_ (.A1(\mod.u_cpu.cpu.immdec.imm7 ),
    .A2(_0390_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2303_ (.A1(_0940_),
    .A2(_0990_),
    .B(_0376_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2304_ (.A1(_0990_),
    .A2(_0619_),
    .B1(_0620_),
    .B2(_0374_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2305_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2306_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .B(_0408_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2307_ (.A1(_0323_),
    .A2(_0325_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2308_ (.A1(_0332_),
    .A2(_0333_),
    .A3(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2309_ (.A1(_0340_),
    .A2(_0515_),
    .A3(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2310_ (.A1(_0321_),
    .A2(_0530_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2311_ (.A1(_0321_),
    .A2(_0529_),
    .B(_0527_),
    .C(_0333_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2312_ (.A1(_0354_),
    .A2(_0626_),
    .B1(_0627_),
    .B2(_0381_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2313_ (.A1(_0625_),
    .A2(_0628_),
    .B(_0342_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2314_ (.A1(_0244_),
    .A2(_0514_),
    .B(_0371_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2315_ (.A1(_0332_),
    .A2(_0371_),
    .B1(_0629_),
    .B2(_0630_),
    .C(_0255_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2316_ (.A1(_0621_),
    .A2(_0622_),
    .B(_0218_),
    .C(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2317_ (.A1(_0926_),
    .A2(_0933_),
    .A3(_1144_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2318_ (.A1(_0958_),
    .A2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2319_ (.A1(_0258_),
    .A2(_0634_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2320_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_0390_),
    .B(_0632_),
    .C(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2321_ (.A1(_0258_),
    .A2(_0634_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2322_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2323_ (.A1(_0636_),
    .A2(_0638_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2324_ (.I(\mod.u_cpu.cpu.immdec.imm30_25[1] ),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2325_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_1045_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _2326_ (.A1(_0325_),
    .A2(_0544_),
    .B1(_0336_),
    .B2(_0349_),
    .C1(_0640_),
    .C2(_0326_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2327_ (.A1(_0349_),
    .A2(_0365_),
    .B1(_0623_),
    .B2(_0354_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2328_ (.A1(_0253_),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2329_ (.A1(_0544_),
    .A2(_0529_),
    .B(_0627_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2330_ (.A1(_0334_),
    .A2(_0349_),
    .B1(_0365_),
    .B2(_0544_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2331_ (.A1(_0625_),
    .A2(_0644_),
    .A3(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2332_ (.A1(_0247_),
    .A2(_0643_),
    .B1(_0646_),
    .B2(_0517_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2333_ (.A1(_0364_),
    .A2(_0641_),
    .B(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2334_ (.A1(_0308_),
    .A2(_0640_),
    .B1(_0648_),
    .B2(_0409_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2335_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_0634_),
    .B(_0376_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2336_ (.A1(_0639_),
    .A2(_0637_),
    .B1(_0649_),
    .B2(_0650_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2337_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_0390_),
    .B(_0635_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2338_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_1045_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2339_ (.A1(_0353_),
    .A2(_0529_),
    .B(_0627_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2340_ (.A1(_0315_),
    .A2(_0392_),
    .B(_0625_),
    .C(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2341_ (.A1(_0335_),
    .A2(_0365_),
    .B1(_0623_),
    .B2(_0353_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2342_ (.A1(_0253_),
    .A2(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2343_ (.A1(_0517_),
    .A2(_0654_),
    .B1(_0656_),
    .B2(_0247_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2344_ (.A1(_0335_),
    .A2(_0339_),
    .B1(_0652_),
    .B2(_0252_),
    .C(_0371_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2345_ (.A1(_0408_),
    .A2(_0657_),
    .A3(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2346_ (.A1(_0408_),
    .A2(_0652_),
    .B(_0659_),
    .C(_0376_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2347_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_0637_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2348_ (.A1(_0651_),
    .A2(_0660_),
    .B(_0661_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2349_ (.A1(_0352_),
    .A2(_0529_),
    .B(_0627_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2350_ (.A1(_0334_),
    .A2(_0357_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2351_ (.A1(_0366_),
    .A2(_0625_),
    .A3(_0662_),
    .A4(_0663_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2352_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_1046_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2353_ (.A1(_0339_),
    .A2(_0357_),
    .B1(_0665_),
    .B2(_0252_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2354_ (.A1(_0371_),
    .A2(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2355_ (.A1(_0517_),
    .A2(_0664_),
    .B(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2356_ (.A1(_0218_),
    .A2(_0634_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2357_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_0637_),
    .B1(_0665_),
    .B2(_0308_),
    .C1(_0669_),
    .C2(\mod.u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2358_ (.A1(_0256_),
    .A2(_0668_),
    .B(_0670_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2359_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2360_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2361_ (.A1(_0310_),
    .A2(_0334_),
    .B(_0516_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2362_ (.A1(_0340_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2363_ (.A1(_0323_),
    .A2(_0310_),
    .B(_0364_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2364_ (.A1(_0323_),
    .A2(_0672_),
    .B(_0675_),
    .C(_0251_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2365_ (.A1(_0517_),
    .A2(_0674_),
    .B(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2366_ (.I(_0669_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2367_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_0635_),
    .B1(_0678_),
    .B2(\mod.u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2368_ (.A1(_0308_),
    .A2(_0672_),
    .B1(_0677_),
    .B2(_0409_),
    .C(_0679_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2369_ (.A1(_0825_),
    .A2(_0926_),
    .B(\mod.u_cpu.cpu.decode.opcode[1] ),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2370_ (.A1(_0940_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2371_ (.A1(_0521_),
    .A2(_0680_),
    .B(_0681_),
    .C(_1156_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2372_ (.A1(\mod.u_cpu.cpu.immdec.imm7 ),
    .A2(_1156_),
    .B(_0669_),
    .C(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2373_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_0637_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2374_ (.A1(_0344_),
    .A2(_0683_),
    .A3(_0684_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2375_ (.A1(_0829_),
    .A2(_1145_),
    .B(_0958_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2376_ (.A1(_0218_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2377_ (.A1(_0258_),
    .A2(_0685_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2378_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_0686_),
    .B1(_0687_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2379_ (.A1(_0540_),
    .A2(_0688_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2381_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2382_ (.A1(_0689_),
    .A2(_0690_),
    .B(_0255_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2383_ (.A1(_0249_),
    .A2(_0333_),
    .B(_0626_),
    .C(_0325_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2384_ (.A1(_0368_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2385_ (.A1(_0353_),
    .A2(_0626_),
    .B(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2386_ (.A1(_0245_),
    .A2(_0353_),
    .A3(_0527_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2387_ (.A1(_0371_),
    .A2(_0382_),
    .B(_0694_),
    .C(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2388_ (.A1(_0691_),
    .A2(_0696_),
    .B(_0390_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2389_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_0686_),
    .B1(_0687_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2390_ (.A1(_0697_),
    .A2(_0698_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2391_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_1045_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2392_ (.A1(_0323_),
    .A2(_0315_),
    .B1(_0562_),
    .B2(_0380_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2393_ (.A1(_0252_),
    .A2(_0699_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2394_ (.A1(_0245_),
    .A2(_0693_),
    .B(_0352_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2395_ (.A1(_0341_),
    .A2(_0626_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2396_ (.A1(_0371_),
    .A2(_0701_),
    .B(_0702_),
    .C(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2397_ (.A1(_0308_),
    .A2(_0699_),
    .B1(_0704_),
    .B2(_0409_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2398_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0686_),
    .B1(_0687_),
    .B2(\mod.u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_0705_),
    .A2(_0706_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2400_ (.A1(_0317_),
    .A2(_0404_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2401_ (.A1(_0241_),
    .A2(_0336_),
    .B(_0313_),
    .C(_0244_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2402_ (.A1(_0544_),
    .A2(_0626_),
    .A3(_0707_),
    .B1(_0708_),
    .B2(_0693_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2403_ (.A1(_1046_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2404_ (.A1(_0215_),
    .A2(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2405_ (.A1(_0325_),
    .A2(_0711_),
    .B(_0675_),
    .C(_0339_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2406_ (.A1(_0256_),
    .A2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2407_ (.A1(_0376_),
    .A2(_0685_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2408_ (.I(\mod.u_cpu.cpu.immdec.imm24_20[4] ),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(_0715_),
    .A2(_0686_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(_0308_),
    .A2(_0711_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2411_ (.A1(\mod.u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_0714_),
    .B(_0716_),
    .C(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2412_ (.A1(_0709_),
    .A2(_0713_),
    .B(_0718_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2413_ (.I0(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_1045_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2414_ (.A1(_0308_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2415_ (.A1(_0381_),
    .A2(_0543_),
    .A3(_0707_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2416_ (.A1(_0311_),
    .A2(_0334_),
    .B(_0626_),
    .C(_0247_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2417_ (.A1(_0315_),
    .A2(_0721_),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2418_ (.A1(_0249_),
    .A2(_0311_),
    .B1(_0719_),
    .B2(_0252_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2419_ (.A1(_0247_),
    .A2(_0314_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2420_ (.A1(_0364_),
    .A2(_0724_),
    .B1(_0725_),
    .B2(_0253_),
    .C(_0256_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2421_ (.A1(\mod.u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_0376_),
    .B1(_0723_),
    .B2(_0726_),
    .C(_0687_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2422_ (.A1(_0715_),
    .A2(_0687_),
    .B1(_0720_),
    .B2(_0727_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2423_ (.A1(_0834_),
    .A2(_0390_),
    .B(_0649_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2424_ (.A1(_0997_),
    .A2(_0390_),
    .B(_0705_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2425_ (.A1(\mod.u_cpu.cpu.decode.op21 ),
    .A2(_0259_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2426_ (.A1(_0697_),
    .A2(_0728_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2427_ (.A1(\mod.u_cpu.cpu.decode.co_ebreak ),
    .A2(_0259_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2428_ (.A1(_0540_),
    .A2(_0729_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2429_ (.A1(_0838_),
    .A2(_0390_),
    .B(_0551_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2430_ (.A1(_0837_),
    .A2(_0390_),
    .B(_0559_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2431_ (.A1(_0839_),
    .A2(_0390_),
    .B(_0565_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2432_ (.A1(_0245_),
    .A2(_0252_),
    .A3(_0355_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2433_ (.A1(_0730_),
    .A2(_0534_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2434_ (.A1(_0408_),
    .A2(_0354_),
    .B1(_0531_),
    .B2(_0341_),
    .C(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2435_ (.A1(_0926_),
    .A2(_0259_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2436_ (.A1(_0259_),
    .A2(_0732_),
    .B(_0733_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2437_ (.A1(_0334_),
    .A2(_0341_),
    .B1(_0353_),
    .B2(_0408_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2438_ (.A1(\mod.u_cpu.cpu.decode.opcode[1] ),
    .A2(_0259_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2439_ (.A1(_0259_),
    .A2(_0734_),
    .B(_0735_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2440_ (.A1(_0241_),
    .A2(_0384_),
    .A3(_0534_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2441_ (.A1(_0244_),
    .A2(_0251_),
    .A3(_0736_),
    .B1(_0381_),
    .B2(_0368_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2442_ (.A1(_0390_),
    .A2(_0255_),
    .A3(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2443_ (.A1(_0825_),
    .A2(_0259_),
    .B1(_0308_),
    .B2(_0352_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2444_ (.A1(_0738_),
    .A2(_0739_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2445_ (.A1(_0247_),
    .A2(_0249_),
    .B1(_0408_),
    .B2(_0313_),
    .C(_0258_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2446_ (.A1(_0368_),
    .A2(_0721_),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2447_ (.A1(_0933_),
    .A2(_0390_),
    .B(_0741_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2448_ (.A1(_0408_),
    .A2(_0314_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2449_ (.A1(_0341_),
    .A2(_0381_),
    .B(_0395_),
    .C(_0376_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2450_ (.A1(_0828_),
    .A2(_0259_),
    .B1(_0742_),
    .B2(_0743_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2451_ (.I(_1177_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2452_ (.A1(_0863_),
    .A2(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .B(_0928_),
    .C(_0864_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2453_ (.A1(_0863_),
    .A2(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2454_ (.A1(_0958_),
    .A2(_0745_),
    .A3(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2455_ (.A1(_0949_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2456_ (.A1(_1177_),
    .A2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2457_ (.I(_0749_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2458_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2459_ (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2460_ (.A1(_0949_),
    .A2(_0747_),
    .B(_1177_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2461_ (.A1(_0752_),
    .A2(_1168_),
    .B(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2462_ (.A1(_0751_),
    .A2(_1168_),
    .B(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2463_ (.A1(_0577_),
    .A2(_0744_),
    .B1(_0750_),
    .B2(_0751_),
    .C(_0755_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2464_ (.I(_0753_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2465_ (.I(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2466_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2467_ (.A1(_1168_),
    .A2(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2468_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_1168_),
    .B(_0757_),
    .C(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2469_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_0744_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2470_ (.A1(_0760_),
    .A2(_0761_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2471_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .B(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2472_ (.A1(_1168_),
    .A2(_1169_),
    .A3(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2473_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_1168_),
    .B(_0757_),
    .C(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2474_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_0744_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2475_ (.A1(_0764_),
    .A2(_0765_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2476_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_1169_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2477_ (.A1(_1168_),
    .A2(_1170_),
    .A3(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2478_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1168_),
    .B(_0757_),
    .C(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2479_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .A2(_0744_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(_0768_),
    .A2(_0769_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2481_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_1170_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2482_ (.A1(_1168_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2483_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_1168_),
    .B(_0757_),
    .C(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2484_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_0744_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2485_ (.A1(_0772_),
    .A2(_0773_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2486_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_0744_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2487_ (.A1(_1175_),
    .A2(_0757_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2488_ (.A1(_0774_),
    .A2(_0775_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2489_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .C2(_0750_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2490_ (.I(_0776_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(_0749_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2492_ (.I(_1177_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2493_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_0757_),
    .B1(_0777_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .C1(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .C2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2494_ (.I(_0779_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2495_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .C2(_0750_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2496_ (.I(_0780_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2497_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .C2(_0750_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2498_ (.I(_0781_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2499_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .C2(_0750_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2500_ (.I(_0782_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2501_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .C2(_0750_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2502_ (.I(_0783_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2503_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .C2(_0750_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2504_ (.I(_0784_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2505_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .C2(_0750_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2506_ (.I(_0785_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2507_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_0744_),
    .B1(_0757_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .C1(_0777_),
    .C2(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2508_ (.I(_0786_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2509_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_0744_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .C1(_0777_),
    .C2(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2510_ (.I(_0787_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2511_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .C2(_0750_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2512_ (.I(_0788_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2513_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .C2(_0750_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2514_ (.I(_0789_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2515_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .C2(_0777_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2516_ (.I(_0790_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2517_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .C2(_0777_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2518_ (.I(_0791_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2519_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .C2(_0777_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2520_ (.I(_0792_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2521_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .C2(_0777_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2522_ (.I(_0793_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2523_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .C2(_0777_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2524_ (.I(_0794_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2525_ (.A1(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_0757_),
    .B1(_0777_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .C1(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .C2(_0778_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2526_ (.I(_0795_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2527_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .C2(_0777_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2528_ (.I(_0796_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2529_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .C2(_0777_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2530_ (.I(_0797_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2531_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .C2(_0777_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2532_ (.I(_0798_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2533_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .C2(_0777_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2534_ (.I(_0799_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2535_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .C2(_0777_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2536_ (.I(_0800_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2537_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .C2(_0777_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2538_ (.I(_0801_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2539_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_0778_),
    .B1(_0756_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .C1(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .C2(_0777_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2540_ (.I(_0802_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2541_ (.A1(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_0744_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2542_ (.A1(_0501_),
    .A2(_0757_),
    .B1(_0750_),
    .B2(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2543_ (.A1(_0803_),
    .A2(_0804_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2544_ (.A1(_0938_),
    .A2(\mod.u_cpu.cpu.state.init_done ),
    .B(_1036_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2545_ (.A1(_0938_),
    .A2(_1143_),
    .B(_0805_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2546_ (.A1(_1036_),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2547_ (.I(_0806_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2548_ (.A1(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .A2(_0928_),
    .A3(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .A4(_0210_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2549_ (.I(_0807_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2550_ (.A1(_0944_),
    .A2(\mod.u_cpu.cpu.ctrl.i_jump ),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2551_ (.A1(_0838_),
    .A2(_0508_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2552_ (.A1(_0944_),
    .A2(_1143_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2553_ (.A1(_0926_),
    .A2(_0809_),
    .B(_0810_),
    .C(_0827_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2554_ (.A1(_0808_),
    .A2(_0811_),
    .B(_1035_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2555_ (.A1(_0825_),
    .A2(_0827_),
    .A3(_1166_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2556_ (.A1(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_0944_),
    .B1(_0810_),
    .B2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2557_ (.A1(_1035_),
    .A2(_0813_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2558_ (.I(\mod.u_cpu.rf_ram_if.rgnt ),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2559_ (.A1(_0814_),
    .A2(_1180_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2560_ (.A1(_0944_),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .B1(_0990_),
    .B2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2561_ (.A1(_1035_),
    .A2(_0816_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2562_ (.A1(_1036_),
    .A2(\mod.u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(_0817_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2564_ (.A1(_1035_),
    .A2(_1001_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2565_ (.A1(\mod.u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\mod.u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2566_ (.A1(_1035_),
    .A2(_0267_),
    .A3(_0818_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2567_ (.A1(_0928_),
    .A2(_0267_),
    .B(_1036_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2568_ (.A1(_0928_),
    .A2(_0267_),
    .B(_0819_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2569_ (.A1(_0928_),
    .A2(_0267_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2570_ (.A1(\mod.u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2571_ (.A1(_1035_),
    .A2(_0821_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2572_ (.A1(_0944_),
    .A2(_1035_),
    .A3(_1143_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2573_ (.D(_0027_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2574_ (.D(_0000_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2575_ (.D(_0001_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2576_ (.D(_0002_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2577_ (.D(_0003_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2578_ (.D(_0004_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2579_ (.D(_0005_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2580_ (.D(_0006_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2581_ (.D(_0007_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2582_ (.D(_0008_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2583_ (.D(_0009_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2584_ (.D(_0010_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2585_ (.D(_0011_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2586_ (.D(_0012_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2587_ (.D(_0028_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2588_ (.D(\mod.u_cpu.cpu.o_wen1 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2589_ (.D(\mod.u_cpu.cpu.o_wen0 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2590_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2591_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2592_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2593_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2594_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2595_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2596_ (.D(\mod.u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2597_ (.D(\mod.u_cpu.cpu.o_wdata1 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2598_ (.D(_0029_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2599_ (.D(_0030_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2600_ (.D(_0031_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2601_ (.D(_0032_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2602_ (.D(\mod.u_cpu.rf_ram_if.rtrig0 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2603_ (.D(_0033_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2604_ (.D(_0034_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2605_ (.D(_0035_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2606_ (.D(\mod.u_cpu.rf_ram_if.wtrig0 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2607_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2608_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2609_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2610_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2611_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2612_ (.D(\mod.u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2613_ (.D(\mod.u_cpu.cpu.o_wdata0 ),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2614_ (.D(_0036_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2615_ (.D(_0025_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2616_ (.D(_0017_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2617_ (.D(_0018_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2618_ (.D(_0019_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2619_ (.D(_0020_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2620_ (.D(_0021_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2621_ (.D(_0022_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2622_ (.D(_0023_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2623_ (.D(_0024_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2624_ (.D(_0037_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2625_ (.D(_0038_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2626_ (.D(_0039_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2627_ (.D(_0040_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2628_ (.D(_0041_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2629_ (.D(_0042_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2630_ (.D(_0043_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2631_ (.D(_0044_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2632_ (.D(_0045_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2633_ (.D(_0046_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2634_ (.D(_0047_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2635_ (.D(_0048_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2636_ (.D(_0049_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2637_ (.D(_0050_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2638_ (.D(_0051_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2639_ (.D(_0052_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2640_ (.D(_0053_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2641_ (.D(_0054_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2642_ (.D(_0055_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2643_ (.D(_0056_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2644_ (.D(_0057_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2645_ (.D(_0058_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2646_ (.D(_0059_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2647_ (.D(_0060_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2648_ (.D(_0061_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2649_ (.D(_0062_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2650_ (.D(_0063_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2651_ (.D(_0064_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2652_ (.D(_0065_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2653_ (.D(_0066_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2654_ (.D(_0067_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2655_ (.D(_0068_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2656_ (.D(_0069_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2657_ (.D(_0013_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2658_ (.D(_0070_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2659_ (.D(_0071_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2660_ (.D(_0072_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2661_ (.D(_0073_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2662_ (.D(_0074_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2663_ (.D(_0075_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2664_ (.D(_0076_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2665_ (.D(_0077_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2666_ (.D(_0078_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2667_ (.D(_0079_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2668_ (.D(_0080_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2669_ (.D(_0081_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2670_ (.D(_0082_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2671_ (.D(_0083_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2672_ (.D(_0084_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2673_ (.D(_0085_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2674_ (.D(_0086_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2675_ (.D(_0087_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2676_ (.D(_0088_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2677_ (.D(_0089_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2678_ (.D(_0090_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2679_ (.D(_0091_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2680_ (.D(_0092_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2681_ (.D(_0093_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2682_ (.D(_0094_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2683_ (.D(_0095_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2684_ (.D(_0096_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2685_ (.D(_0097_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2686_ (.D(_0098_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2687_ (.D(_0099_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2688_ (.D(_0100_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2689_ (.D(_0101_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2690_ (.D(_0015_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2691_ (.D(_0016_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2692_ (.D(_0102_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2693_ (.D(_0103_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2694_ (.D(_0014_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2695_ (.D(_0104_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2696_ (.D(_0105_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2697_ (.D(_0106_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2698_ (.D(_0107_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2699_ (.D(_0108_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2700_ (.D(_0109_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2701_ (.D(_0110_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2702_ (.D(_0111_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2703_ (.D(_0112_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2704_ (.D(_0113_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2705_ (.D(_0114_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2706_ (.D(_0115_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2707_ (.D(_0116_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2708_ (.D(_0117_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2709_ (.D(_0118_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2710_ (.D(_0119_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2711_ (.D(_0120_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2712_ (.D(_0121_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2713_ (.D(_0122_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2714_ (.D(_0123_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2715_ (.D(_0124_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2716_ (.D(_0125_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2717_ (.D(_0126_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2718_ (.D(_0127_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2719_ (.D(_0128_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2720_ (.D(_0129_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2721_ (.D(_0130_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2722_ (.D(_0131_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2723_ (.D(_0132_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2724_ (.D(_0133_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2725_ (.D(_0134_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2726_ (.D(_0135_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2727_ (.D(_0136_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2728_ (.D(_0137_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2729_ (.D(_0138_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2730_ (.D(_0139_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2731_ (.D(_0140_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2732_ (.D(_0141_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2733_ (.D(_0142_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2734_ (.D(_0143_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2735_ (.D(_0144_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2736_ (.D(_0145_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2737_ (.D(_0146_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2738_ (.D(_0147_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2739_ (.D(_0148_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2740_ (.D(_0149_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2741_ (.D(_0150_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2742_ (.D(_0151_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2743_ (.D(_0152_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2744_ (.D(_0153_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2745_ (.D(_0154_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2746_ (.D(_0155_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2747_ (.D(_0156_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2748_ (.D(_0157_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2749_ (.D(_0158_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2750_ (.D(_0159_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2751_ (.D(_0160_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2752_ (.D(_0161_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2753_ (.D(_0162_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2754_ (.D(_0163_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2755_ (.D(_0164_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2756_ (.D(_0165_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2757_ (.D(_0166_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2758_ (.D(_0167_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2759_ (.D(_0168_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2760_ (.D(_0169_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2761_ (.D(_0170_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2762_ (.D(_0171_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2763_ (.D(_0172_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2764_ (.D(_0173_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2765_ (.D(_0174_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2766_ (.D(_0175_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2767_ (.D(_0176_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2768_ (.D(_0177_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2769_ (.D(_0178_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2770_ (.D(_0179_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2771_ (.D(_0180_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2772_ (.D(_0181_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2773_ (.D(_0182_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2774_ (.D(_0183_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2775_ (.D(_0184_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2776_ (.D(_0185_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2777_ (.D(_0186_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2778_ (.D(_0187_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2779_ (.D(_0188_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2780_ (.D(_0189_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2781_ (.D(_0190_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2782_ (.D(_0191_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2783_ (.D(_0192_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2784_ (.D(_0193_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2785_ (.D(_0194_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2786_ (.D(_0195_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2787_ (.D(_0196_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2788_ (.D(_0197_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2789_ (.D(_0198_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2790_ (.D(_0199_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2791_ (.D(_0200_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2792_ (.D(_0201_),
    .CLK(io_in[12]),
    .Q(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2793_ (.D(_0202_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2794_ (.D(_0203_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2795_ (.D(_0204_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2796_ (.D(_0205_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2797_ (.D(_0206_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2798_ (.D(_0207_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2799_ (.D(_0208_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2800_ (.D(_0209_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2801_ (.D(_0210_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2802_ (.D(_0211_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2803_ (.D(_0212_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2804_ (.D(_0213_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _2805_ (.D(_0214_),
    .CLK(io_in[12]),
    .Q(\mod.u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2806_ (.Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2807_ (.Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2808_ (.Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2809_ (.Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2810_ (.Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2811_ (.Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2812_ (.Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2813_ (.Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2814_ (.Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2815_ (.Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2816_ (.Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2817_ (.Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2818_ (.Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2819_ (.Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2820_ (.Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2821_ (.Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2822_ (.Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2823_ (.Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2824_ (.Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2825_ (.Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2826_ (.Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2827_ (.Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2828_ (.Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2829_ (.Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2830_ (.Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2831_ (.Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2832_ (.Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2833_ (.Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2834_ (.Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2835_ (.Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2836_ (.Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2837_ (.Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2838_ (.Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2839_ (.Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2840_ (.Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2841_ (.Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2842_ (.Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2843_ (.Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2844_ (.Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2845_ (.Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2846_ (.Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2847_ (.Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2848_ (.Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2849_ (.Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2850_ (.Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2851_ (.Z(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2852_ (.Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2853_ (.Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2854_ (.Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2855_ (.Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2856_ (.Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2857_ (.Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2858_ (.Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2859_ (.Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2860_ (.Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2861_ (.Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2862_ (.Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2863_ (.Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2864_ (.Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2865_ (.Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2866_ (.Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2867_ (.Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2868_ (.Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2869_ (.Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2870_ (.Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2871_ (.Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2872_ (.Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2873_ (.Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2874_ (.Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2875_ (.Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2876_ (.Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2877_ (.Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2878_ (.Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _2879_ (.Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2880_ (.ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2881_ (.ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2882_ (.ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2883_ (.ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2884_ (.ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2885_ (.ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2886_ (.ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2887_ (.ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2888_ (.ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2889_ (.ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2890_ (.ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2891_ (.ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2892_ (.ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2893_ (.ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2894_ (.ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2895_ (.ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2896_ (.ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2897_ (.ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2898_ (.ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2899_ (.ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2900_ (.ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2901_ (.ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2902_ (.ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2903_ (.ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2904_ (.ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2905_ (.ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2906_ (.ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2907_ (.ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2908_ (.ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2909_ (.ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2910_ (.ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2911_ (.ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2912_ (.ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2913_ (.ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2914_ (.ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2915_ (.ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2916_ (.ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2917_ (.ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2918_ (.ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2919_ (.ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2920_ (.ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2921_ (.ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2922_ (.ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2923_ (.ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2924_ (.ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2925_ (.ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2926_ (.ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2927_ (.ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2928_ (.ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2929_ (.ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2930_ (.ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2931_ (.ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2932_ (.ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2933_ (.ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2934_ (.ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2935_ (.ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2936_ (.ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2937_ (.ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2938_ (.ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2939_ (.ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2940_ (.ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2941_ (.ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2942_ (.ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2943_ (.ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2944_ (.ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2945_ (.ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2946_ (.ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2947_ (.ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2948_ (.ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2949_ (.ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2950_ (.ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2951_ (.ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2952_ (.ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2953_ (.ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2954_ (.ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2955_ (.ZN(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2956_ (.ZN(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2957_ (.ZN(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2958_ (.ZN(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2959_ (.ZN(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2960_ (.ZN(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2961_ (.ZN(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2962_ (.ZN(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2963_ (.ZN(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2964_ (.ZN(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2965_ (.ZN(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2966_ (.ZN(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2967_ (.ZN(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2968_ (.ZN(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2969_ (.ZN(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2970_ (.ZN(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2971_ (.ZN(io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2972_ (.ZN(io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2973_ (.ZN(io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2974_ (.ZN(io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2975_ (.ZN(io_oeb[20]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2976_ (.ZN(io_oeb[21]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2977_ (.ZN(io_oeb[22]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2978_ (.ZN(io_oeb[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2979_ (.ZN(io_oeb[24]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2980_ (.ZN(io_oeb[25]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2981_ (.ZN(io_oeb[26]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2982_ (.ZN(io_oeb[27]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2983_ (.ZN(io_oeb[28]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2984_ (.ZN(io_oeb[29]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2985_ (.ZN(io_oeb[30]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2986_ (.ZN(io_oeb[31]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2987_ (.ZN(io_oeb[32]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2988_ (.ZN(io_oeb[33]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2989_ (.ZN(io_oeb[34]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2990_ (.ZN(io_oeb[35]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2991_ (.ZN(io_oeb[36]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2992_ (.ZN(io_oeb[37]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2993_ (.ZN(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2994_ (.ZN(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2995_ (.ZN(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2996_ (.ZN(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2997_ (.ZN(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2998_ (.ZN(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _2999_ (.ZN(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3000_ (.ZN(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3001_ (.ZN(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3002_ (.ZN(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3003_ (.ZN(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3004_ (.ZN(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3005_ (.ZN(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3006_ (.ZN(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3007_ (.ZN(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3008_ (.ZN(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3009_ (.ZN(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3010_ (.ZN(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3011_ (.ZN(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3012_ (.ZN(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3013_ (.ZN(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3014_ (.ZN(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3015_ (.ZN(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3016_ (.ZN(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3017_ (.ZN(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3018_ (.ZN(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3019_ (.ZN(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3020_ (.ZN(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3021_ (.ZN(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3022_ (.ZN(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3023_ (.ZN(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3024_ (.ZN(io_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3025_ (.ZN(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3026_ (.ZN(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3027_ (.ZN(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3028_ (.ZN(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3029_ (.ZN(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3030_ (.ZN(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3031_ (.ZN(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3032_ (.ZN(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3033_ (.ZN(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3034_ (.ZN(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3035_ (.ZN(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3036_ (.ZN(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3037_ (.ZN(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3038_ (.ZN(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3039_ (.ZN(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3040_ (.ZN(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3041_ (.ZN(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3042_ (.ZN(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3043_ (.ZN(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3044_ (.ZN(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3045_ (.ZN(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3046_ (.ZN(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3047_ (.ZN(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3048_ (.ZN(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3049_ (.ZN(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3050_ (.ZN(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3051_ (.ZN(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3052_ (.ZN(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3053_ (.ZN(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3054_ (.ZN(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3055_ (.ZN(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3056_ (.ZN(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3057_ (.ZN(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3058_ (.ZN(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3059_ (.ZN(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3060_ (.ZN(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3061_ (.ZN(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3062_ (.ZN(la_data_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3063_ (.ZN(la_data_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3064_ (.ZN(la_data_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3065_ (.ZN(la_data_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3066_ (.ZN(la_data_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3067_ (.ZN(la_data_out[38]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3068_ (.ZN(la_data_out[39]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3069_ (.ZN(la_data_out[40]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3070_ (.ZN(la_data_out[41]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3071_ (.ZN(la_data_out[42]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3072_ (.ZN(la_data_out[43]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3073_ (.ZN(la_data_out[44]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3074_ (.ZN(la_data_out[45]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3075_ (.ZN(la_data_out[46]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3076_ (.ZN(la_data_out[47]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3077_ (.ZN(la_data_out[48]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3078_ (.ZN(la_data_out[49]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3079_ (.ZN(la_data_out[50]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3080_ (.ZN(la_data_out[51]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3081_ (.ZN(la_data_out[52]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3082_ (.ZN(la_data_out[53]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3083_ (.ZN(la_data_out[54]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3084_ (.ZN(la_data_out[55]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3085_ (.ZN(la_data_out[56]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3086_ (.ZN(la_data_out[57]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3087_ (.ZN(la_data_out[58]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3088_ (.ZN(la_data_out[59]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3089_ (.ZN(la_data_out[60]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3090_ (.ZN(la_data_out[61]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3091_ (.ZN(la_data_out[62]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3092_ (.ZN(la_data_out[63]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3093_ (.ZN(user_irq[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3094_ (.ZN(user_irq[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3095_ (.ZN(user_irq[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3096_ (.ZN(wbs_ack_o));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3097_ (.ZN(wbs_dat_o[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3098_ (.ZN(wbs_dat_o[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3099_ (.ZN(wbs_dat_o[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3100_ (.ZN(wbs_dat_o[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3101_ (.ZN(wbs_dat_o[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3102_ (.ZN(wbs_dat_o[5]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3103_ (.ZN(wbs_dat_o[6]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3104_ (.ZN(wbs_dat_o[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3105_ (.ZN(wbs_dat_o[8]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3106_ (.ZN(wbs_dat_o[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3107_ (.ZN(wbs_dat_o[10]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3108_ (.ZN(wbs_dat_o[11]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3109_ (.ZN(wbs_dat_o[12]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3110_ (.ZN(wbs_dat_o[13]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3111_ (.ZN(wbs_dat_o[14]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3112_ (.ZN(wbs_dat_o[15]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3113_ (.ZN(wbs_dat_o[16]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3114_ (.ZN(wbs_dat_o[17]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3115_ (.ZN(wbs_dat_o[18]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3116_ (.ZN(wbs_dat_o[19]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3117_ (.ZN(wbs_dat_o[20]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3118_ (.ZN(wbs_dat_o[21]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3119_ (.ZN(wbs_dat_o[22]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3120_ (.ZN(wbs_dat_o[23]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3121_ (.ZN(wbs_dat_o[24]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3122_ (.ZN(wbs_dat_o[25]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3123_ (.ZN(wbs_dat_o[26]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3124_ (.ZN(wbs_dat_o[27]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3125_ (.ZN(wbs_dat_o[28]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3126_ (.ZN(wbs_dat_o[29]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3127_ (.ZN(wbs_dat_o[30]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _3128_ (.ZN(wbs_dat_o[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3129_ (.I(\mod.u_scanchain_local.clk_out ),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3130_ (.I(\mod.u_scanchain_local.data_out ),
    .Z(io_out[14]));
 gf180mcu_fd_ip_sram__sram256x8m8wm1 \mod.u_cpu.rf_ram.RAM0  (.CEN(_1256_),
    .CLK(io_in[12]),
    .GWEN(_0026_),
    .A({\mod.u_cpu.rf_ram.addr[7] ,
    \mod.u_cpu.rf_ram.addr[6] ,
    \mod.u_cpu.rf_ram.addr[5] ,
    \mod.u_cpu.rf_ram.addr[4] ,
    \mod.u_cpu.rf_ram.addr[3] ,
    \mod.u_cpu.rf_ram.addr[2] ,
    \mod.u_cpu.rf_ram.addr[1] ,
    \mod.u_cpu.rf_ram.addr[0] }),
    .D({\mod.u_cpu.rf_ram.i_wdata[7] ,
    \mod.u_cpu.rf_ram.i_wdata[6] ,
    \mod.u_cpu.rf_ram.i_wdata[5] ,
    \mod.u_cpu.rf_ram.i_wdata[4] ,
    \mod.u_cpu.rf_ram.i_wdata[3] ,
    \mod.u_cpu.rf_ram.i_wdata[2] ,
    \mod.u_cpu.rf_ram.i_wdata[1] ,
    \mod.u_cpu.rf_ram.i_wdata[0] }),
    .Q({\mod.u_cpu.rf_ram.data[7] ,
    \mod.u_cpu.rf_ram.data[6] ,
    \mod.u_cpu.rf_ram.data[5] ,
    \mod.u_cpu.rf_ram.data[4] ,
    \mod.u_cpu.rf_ram.data[3] ,
    \mod.u_cpu.rf_ram.data[2] ,
    \mod.u_cpu.rf_ram.data[1] ,
    \mod.u_cpu.rf_ram.data[0] }),
    .WEN({_0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_,
    _0026_}));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \mod.u_scanchain_local.input_buf_clk  (.I(io_in[8]),
    .Z(\mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \mod.u_scanchain_local.out_flop  (.D(\mod.u_scanchain_local.module_data_in[69] ),
    .CLKN(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \mod.u_scanchain_local.output_buffers[2]  (.I(\mod.u_scanchain_local.data_out_i ),
    .Z(\mod.u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \mod.u_scanchain_local.output_buffers[3]  (.I(\clknet_opt_1_1_mod.u_scanchain_local.clk ),
    .Z(\mod.u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[0]  (.D(io_in[10]),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_cyc ),
    .CLK(\clknet_3_2__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[10]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[11]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[12]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[13]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[14]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[15]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[16]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[17]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[18]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[19]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[1]  (.D(\mod.timer_irq ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_we ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[20]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[21]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[22]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[23]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[24]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[25]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[26]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[27]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[28]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[29]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[2]  (.D(\mod.u_arbiter.i_wb_cpu_ack ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[30]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[31]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[32]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[33]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[34]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[35]  (.D(\mod.u_scanchain_local.module_data_in[34] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[36]  (.D(\mod.u_scanchain_local.module_data_in[35] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[37]  (.D(\mod.u_scanchain_local.module_data_in[36] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[38]  (.D(\mod.u_scanchain_local.module_data_in[37] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[39]  (.D(\mod.u_scanchain_local.module_data_in[38] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[3]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[40]  (.D(\mod.u_scanchain_local.module_data_in[39] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[41]  (.D(\mod.u_scanchain_local.module_data_in[40] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[42]  (.D(\mod.u_scanchain_local.module_data_in[41] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(\clknet_3_0__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[43]  (.D(\mod.u_scanchain_local.module_data_in[42] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[44]  (.D(\mod.u_scanchain_local.module_data_in[43] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[45]  (.D(\mod.u_scanchain_local.module_data_in[44] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[46]  (.D(\mod.u_scanchain_local.module_data_in[45] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[47]  (.D(\mod.u_scanchain_local.module_data_in[46] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[48]  (.D(\mod.u_scanchain_local.module_data_in[47] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(\clknet_3_5__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[49]  (.D(\mod.u_scanchain_local.module_data_in[48] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[4]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[50]  (.D(\mod.u_scanchain_local.module_data_in[49] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[51]  (.D(\mod.u_scanchain_local.module_data_in[50] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[52]  (.D(\mod.u_scanchain_local.module_data_in[51] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[53]  (.D(\mod.u_scanchain_local.module_data_in[52] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[54]  (.D(\mod.u_scanchain_local.module_data_in[53] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[55]  (.D(\mod.u_scanchain_local.module_data_in[54] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[56]  (.D(\mod.u_scanchain_local.module_data_in[55] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(\clknet_3_7__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[57]  (.D(\mod.u_scanchain_local.module_data_in[56] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[58]  (.D(\mod.u_scanchain_local.module_data_in[57] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[59]  (.D(\mod.u_scanchain_local.module_data_in[58] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[5]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[60]  (.D(\mod.u_scanchain_local.module_data_in[59] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[61]  (.D(\mod.u_scanchain_local.module_data_in[60] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(\clknet_3_2__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[62]  (.D(\mod.u_scanchain_local.module_data_in[61] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[63]  (.D(\mod.u_scanchain_local.module_data_in[62] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[64]  (.D(\mod.u_scanchain_local.module_data_in[63] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(\clknet_3_6__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[65]  (.D(\mod.u_scanchain_local.module_data_in[64] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[66]  (.D(\mod.u_scanchain_local.module_data_in[65] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(\clknet_3_2__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[67]  (.D(\mod.u_scanchain_local.module_data_in[66] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(\clknet_3_2__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[68]  (.D(\mod.u_scanchain_local.module_data_in[67] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[69]  (.D(\mod.u_scanchain_local.module_data_in[68] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(\clknet_3_3__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[6]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[7]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[8]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(\clknet_3_4__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \mod.u_scanchain_local.scan_flop[9]  (.D(\mod.u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(io_in[11]),
    .SI(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(\clknet_3_1__leaf_mod.u_scanchain_local.clk ),
    .Q(\mod.u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_494 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_495 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_496 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_497 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_498 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_499 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_500 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_501 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_502 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_503 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_504 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_505 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_506 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_507 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_508 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_509 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_510 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_511 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_512 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_513 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_514 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_515 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_516 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_517 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_518 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_519 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_520 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_521 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_522 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_0_mod.u_scanchain_local.clk  (.I(\mod.u_scanchain_local.clk ),
    .Z(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_0__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_1__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_2__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_3__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_4__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_5__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_6__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_3_7__f_mod.u_scanchain_local.clk  (.I(\clknet_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_opt_1_0_mod.u_scanchain_local.clk  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ),
    .Z(\clknet_opt_1_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 \clkbuf_opt_1_1_mod.u_scanchain_local.clk  (.I(\clknet_opt_1_0_mod.u_scanchain_local.clk ),
    .Z(\clknet_opt_1_1_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__D (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A2 (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__D (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__A2 (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__D (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__A2 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__D (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__A2 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A2 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A3 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__A2 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__S (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[0]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[1]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[2]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[3]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_GWEN  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[4]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[5]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[7]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_WEN[6]  (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A2 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A2 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__C (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__I (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__A1 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__B (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__B2 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__B (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__C (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__C (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__C (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__C (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__B2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__B2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__B2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__B2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__I (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__C (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2201__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A1 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A2 (.I(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__B2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A2 (.I(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__B2 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A1 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__B (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__C (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__B (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__C (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2406__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__C (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__C (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__C (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__C (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__I (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A2 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1889__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__S (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__B1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__B2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__B2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__B2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A2 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A1 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__B (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__B (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A2 (.I(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__B (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__C2 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__B1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1922__A2 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__B1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1940__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__C (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1937__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1927__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A1 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A2 (.I(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__C (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A4 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1932__C (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__B2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2206__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A3 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2187__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__C (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1935__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__B1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__B2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__B2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__B1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__C (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__C (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__B2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__B (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__B1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__B1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__B (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A2 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A3 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__B (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__B (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__B2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2252__B2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__B (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__B2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__I (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__B2 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__B1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A3 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__B2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__B2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__A4 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A3 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__A3 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1999__A3 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__B2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__B2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__B1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A3 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__B (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A3 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2212__B2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__B (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1972__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1995__C1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__B (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__C (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__C (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__B (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__B2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__C (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__C (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2246__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__C (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__C (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__B2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__B1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__C (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__C (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__B (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__B (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__B (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__C (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A3 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__A1 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__B2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__B (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__B1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2188__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__B1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__B (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__I (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__B2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__B (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__B2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__B (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__C (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__C (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__B2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__B2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2054__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2034__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__B1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2064__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__B1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A2 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2343__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__B2 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__B (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__B1 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__C (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2199__I (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__S (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2215__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__A3 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__B (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A3 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__A2 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__B2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__B1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__B (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__B1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__B (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__B1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__B2 (.I(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2242__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__B (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__B1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__B1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A2 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__C (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__C (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__B1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__I0 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__B (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2383__B (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2312__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2320__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__C1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__B1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__B1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__B (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__C1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__B (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2377__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__C (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__B1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__B1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__B (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__B1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__B (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__C2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__B1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__B (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__B1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__C2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__C1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__C1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__C2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__C2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__C (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1335__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1334__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A3 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__B (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__B (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1337__I (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__A1 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__C (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__C (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1339__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__B (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A4 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1340__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__B2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A3 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1344__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__B (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1348__I (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__B2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__B (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__B (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A2 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__B (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__B (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__B (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1528__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2431__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2171__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1773__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1351__A3 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__B1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__B1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__B1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__B1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__A3 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__C (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1569__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__B (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1391__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__A2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__I (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__S0 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__C (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2100__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__B1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__S1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1461__S (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A3 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__B (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1379__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1399__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1398__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1394__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__C (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1382__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A3 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__B2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A4 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__B2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1445__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1435__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1455__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1453__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__S (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__C (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1503__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__A3 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__B (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__B (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__B1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__B (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A3 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1519__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1491__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__I (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__C (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__I0 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__B (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1509__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A3 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__B (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__A3 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2172__I1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2094__A3 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A3 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__B (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__A4 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A4 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A4 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A4 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A2 (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__I (.I(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__B (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__B (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__B (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__B (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__B (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__B (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A1 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1637__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__B (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1705__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__S (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A4 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2004__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__S (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__S (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__S (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__S (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__S (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__S (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A3 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__A1 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A4 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A4 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__A3 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A3 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A3 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2104__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__B (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__A3 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A3 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__C (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__B (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2149__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__S (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2131__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__S (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__I (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__B (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__B (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__I (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__B (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__I (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1775__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A4 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A2 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__I (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_CEN  (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[0]_D  (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[67]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[68]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[69]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[66]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[63]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[64]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[65]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[57]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[58]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[59]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[60]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[61]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[62]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[56]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[55]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[54]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[38]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[3]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[4]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[5]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[39]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[2]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[1]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[0]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[41]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[40]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[43]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[42]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[53]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[52]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[10]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[14]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[21]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[12]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[20]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[17]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[19]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[11]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[18]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[6]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[7]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[8]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[9]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[16]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[15]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[22]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[23]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[24]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[25]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[26]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[27]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[28]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[13]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[29]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[30]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[31]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[32]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[33]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[37]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[34]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[35]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[36]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[46]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[47]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[48]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[49]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[50]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[51]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[44]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[45]_SE  (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2615__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_CLK  (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2738__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2748__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2677__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2771__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2790__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__CLK (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.input_buf_clk_I  (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[1]_D  (.I(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A3 (.I(\mod.timer_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[2]_D  (.I(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A1 (.I(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__A1 (.I(\mod.u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2125__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2153__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1698__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2109__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2105__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2169__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[6]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__I (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A3 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I0 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[21]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__C2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[22]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[23]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[24]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[7]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2466__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__I (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[26]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[27]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[30]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I3 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[31]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[33]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[8]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__B (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[36]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[37]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[9]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[10]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[11]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[12]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[13]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__B2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[14]_SI  (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__C1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__I2 (.I(\mod.u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1554__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__A1 (.I(\mod.u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[3]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__I (.I(\mod.u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[13]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[14]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[15]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[16]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[17]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[18]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[22]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[4]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[24]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[25]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[26]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__C1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[28]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[30]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[5]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[33]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[6]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1955__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[7]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1954__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[8]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[9]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[11]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__I1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[12]_D  (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A1 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A2 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I0 (.I(\mod.u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A1 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__A2 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__I (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A2 (.I(\mod.u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1727__A1 (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__A2 (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__B (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__I (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1342__A2 (.I(\mod.u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2167__A1 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A1 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__A2 (.I(\mod.u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A2 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__A1 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A1 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__C (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A1 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A3 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__I (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1343__A1 (.I(\mod.u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2245__I (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2243__A1 (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__A1 (.I(\mod.u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A2 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(\mod.u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__B2 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A3 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__A2 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(\mod.u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__I (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A1 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1540__A1 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1483__B1 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1396__A2 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__A2 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1347__A1 (.I(\mod.u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A1 (.I(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1355__A3 (.I(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__A1 (.I(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1344__A1 (.I(\mod.u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__I1 (.I(\mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__I (.I(\mod.u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A2 (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A2 (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__I (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__A2 (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1356__A1 (.I(\mod.u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1395__I (.I(\mod.u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2007__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1404__A1 (.I(\mod.u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1369__A1 (.I(\mod.u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2378__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1365__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__I (.I(\mod.u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1361__B2 (.I(\mod.u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(\mod.u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(\mod.u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(\mod.u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A3 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A3 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1558__B (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__B (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A3 (.I(\mod.u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__A1 (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__B2 (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__A1 (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__I (.I(\mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A2 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A2 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1502__A2 (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__B (.I(\mod.u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A2 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__A1 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__A3 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A3 (.I(\mod.u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[0]  (.I(\mod.u_cpu.rf_ram.addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[1]  (.I(\mod.u_cpu.rf_ram.addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[2]  (.I(\mod.u_cpu.rf_ram.addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[3]  (.I(\mod.u_cpu.rf_ram.addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[4]  (.I(\mod.u_cpu.rf_ram.addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[5]  (.I(\mod.u_cpu.rf_ram.addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[6]  (.I(\mod.u_cpu.rf_ram.addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_A[7]  (.I(\mod.u_cpu.rf_ram.addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__I (.I(\mod.u_cpu.rf_ram.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1418__I1 (.I(\mod.u_cpu.rf_ram.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1423__I1 (.I(\mod.u_cpu.rf_ram.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__I1 (.I(\mod.u_cpu.rf_ram.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__I1 (.I(\mod.u_cpu.rf_ram.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__I1 (.I(\mod.u_cpu.rf_ram.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1443__I1 (.I(\mod.u_cpu.rf_ram.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__I1 (.I(\mod.u_cpu.rf_ram.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[0]  (.I(\mod.u_cpu.rf_ram.i_wdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[1]  (.I(\mod.u_cpu.rf_ram.i_wdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[2]  (.I(\mod.u_cpu.rf_ram.i_wdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[3]  (.I(\mod.u_cpu.rf_ram.i_wdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[4]  (.I(\mod.u_cpu.rf_ram.i_wdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[5]  (.I(\mod.u_cpu.rf_ram.i_wdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[6]  (.I(\mod.u_cpu.rf_ram.i_wdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_cpu.rf_ram.RAM0_D[7]  (.I(\mod.u_cpu.rf_ram.i_wdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2602__D (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1436__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1426__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1421__S (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A2 (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__A2 (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__A1 (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1362__A1 (.I(\mod.u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__D (.I(\mod.u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__I0 (.I(\mod.u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__D (.I(\mod.u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__I0 (.I(\mod.u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__D (.I(\mod.u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__I1 (.I(\mod.u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__D (.I(\mod.u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__I1 (.I(\mod.u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__D (.I(\mod.u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__I1 (.I(\mod.u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__D (.I(\mod.u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1572__A2 (.I(\mod.u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_0_mod.u_scanchain_local.clk_I  (.I(\mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.output_buffers[2]_I  (.I(\mod.u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[37]_D  (.I(\mod.u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[38]_D  (.I(\mod.u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.out_flop_D  (.I(\mod.u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_7__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_6__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_5__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_4__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_3__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_2__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_1__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_3_0__f_mod.u_scanchain_local.clk_I  (.I(\clknet_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[15]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[18]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[19]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[2]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[3]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[40]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[41]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[42]_CLK  (.I(\clknet_3_0__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[13]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[17]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[20]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[21]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[23]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[24]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[35]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[37]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[7]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[9]_CLK  (.I(\clknet_3_1__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_opt_1_0_mod.u_scanchain_local.clk_I  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[0]_CLK  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[61]_CLK  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[66]_CLK  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[67]_CLK  (.I(\clknet_3_2__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[1]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[38]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[39]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[65]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[68]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[69]_CLK  (.I(\clknet_3_3__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[10]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[11]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[28]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[30]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[44]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[45]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[47]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[4]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[5]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[6]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[8]_CLK  (.I(\clknet_3_4__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[12]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[14]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[16]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[22]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[25]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[26]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[27]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[29]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[31]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[32]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[33]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[34]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[36]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[46]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[48]_CLK  (.I(\clknet_3_5__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.out_flop_CLKN  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[55]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[57]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[58]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[59]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[60]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[62]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[63]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[64]_CLK  (.I(\clknet_3_6__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[43]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[49]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[50]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[51]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[52]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[53]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[54]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.scan_flop[56]_CLK  (.I(\clknet_3_7__leaf_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_clkbuf_opt_1_1_mod.u_scanchain_local.clk_I  (.I(\clknet_opt_1_0_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mod.u_scanchain_local.output_buffers[3]_I  (.I(\clknet_opt_1_1_mod.u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
endmodule

